-------------------------------------------------------------------------------
-- Synchronous ROM with generic memory and data sizes
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity rom is
    generic(ADDRESS_BITS: positive;
            DATA_LENGTH:  positive;
            SELECT_ROM:  integer := 0); -- Select which ROM to use
    port(-- Control signals
         Clk: in std_logic;
         Re:  in std_logic;
         
         -- Input signals
         Addr: in std_logic_vector (ADDRESS_BITS - 1 downto 0);
         
         -- Output
         Dout: out std_logic_vector (DATA_LENGTH - 1 downto 0);
         initial_addr_2: out std_logic_vector (ADDRESS_BITS - 1 downto 0);
         initial_addr_3: out std_logic_vector (ADDRESS_BITS - 1 downto 0));
end rom;

architecture Behavioral of rom is

    type MemoryBank is array(0 to 2**ADDRESS_BITS - 1)
                    of std_logic_vector(DATA_LENGTH - 1 downto 0);
    signal bank: MemoryBank;


begin

	gen_rom_0: if SELECT_ROM = 0 generate
		bank <= (
			0 => x"00000005",
			1 => x"00000009",
			2 => x"0000000d",
			3 => x"00000011",
			4 => x"00000015",
			5 => x"00000019",
			6 => x"0000001d",
			7 => x"00000021",
			8 => x"00000025",
			9 => x"00000029",
			10 => x"0000002d",
			11 => x"00000031",
			12 => x"00000035",
			13 => x"00000039",
			14 => x"0000003d",
			15 => x"00000041",
			16 => x"00000045",
			17 => x"00000049",
			18 => x"0000004d",
			19 => x"00000051",
			20 => x"00000055",
			21 => x"00000059",
			22 => x"0000005d",
			23 => x"00000061",
			24 => x"00000065",
			25 => x"00000069",
			26 => x"0000006d",
			27 => x"00000071",
			28 => x"00000075",
			29 => x"00000079",
			30 => x"0000007d",
			31 => x"00000081",
			32 => x"00000085",
			33 => x"00000089",
			34 => x"0000008d",
			35 => x"00000091",
			36 => x"00000095",
			37 => x"0f05da04",
			38 => x"000000a1",
			39 => x"ffe600a1",
			40 => x"0f058504",
			41 => x"000000ad",
			42 => x"fff200ad",
			43 => x"0007e504",
			44 => x"ffe700b9",
			45 => x"000000b9",
			46 => x"0007e504",
			47 => x"ffed00c5",
			48 => x"000000c5",
			49 => x"0f058504",
			50 => x"000000d1",
			51 => x"ffee00d1",
			52 => x"0f05d208",
			53 => x"0e032004",
			54 => x"000000e5",
			55 => x"000e00e5",
			56 => x"ffe100e5",
			57 => x"0007ba08",
			58 => x"0f055a04",
			59 => x"00000101",
			60 => x"ff990101",
			61 => x"0e032604",
			62 => x"00000101",
			63 => x"00160101",
			64 => x"0006ce04",
			65 => x"ff0c011d",
			66 => x"06014d08",
			67 => x"09002504",
			68 => x"007f011d",
			69 => x"0000011d",
			70 => x"0000011d",
			71 => x"0900270c",
			72 => x"06014d08",
			73 => x"0505f604",
			74 => x"00000139",
			75 => x"00880139",
			76 => x"00000139",
			77 => x"ff320139",
			78 => x"0100160c",
			79 => x"0e02bd04",
			80 => x"00000155",
			81 => x"0f05da04",
			82 => x"000b0155",
			83 => x"00000155",
			84 => x"00000155",
			85 => x"0f05da0c",
			86 => x"0c056304",
			87 => x"00000171",
			88 => x"0c05be04",
			89 => x"00230171",
			90 => x"00000171",
			91 => x"00000171",
			92 => x"0f05da0c",
			93 => x"0c05be08",
			94 => x"0c052804",
			95 => x"0000018d",
			96 => x"001e018d",
			97 => x"0000018d",
			98 => x"0000018d",
			99 => x"0900270c",
			100 => x"0f05da08",
			101 => x"0006ce04",
			102 => x"000001a9",
			103 => x"000601a9",
			104 => x"000001a9",
			105 => x"000001a9",
			106 => x"0007ba08",
			107 => x"09002004",
			108 => x"000001cd",
			109 => x"fec501cd",
			110 => x"0c059b08",
			111 => x"0208f704",
			112 => x"00cf01cd",
			113 => x"000001cd",
			114 => x"000001cd",
			115 => x"0415f304",
			116 => x"fe9301f1",
			117 => x"0208900c",
			118 => x"03037b04",
			119 => x"000001f1",
			120 => x"09002704",
			121 => x"013101f1",
			122 => x"000001f1",
			123 => x"000001f1",
			124 => x"01001810",
			125 => x"0c05be0c",
			126 => x"0505ea04",
			127 => x"00000215",
			128 => x"0f05da04",
			129 => x"00750215",
			130 => x"00000215",
			131 => x"00000215",
			132 => x"ff200215",
			133 => x"0f05da10",
			134 => x"0705d20c",
			135 => x"0c052504",
			136 => x"00000239",
			137 => x"09002604",
			138 => x"00620239",
			139 => x"00000239",
			140 => x"00000239",
			141 => x"ff620239",
			142 => x"01001810",
			143 => x"0c05a40c",
			144 => x"07054504",
			145 => x"0000025d",
			146 => x"0f05da04",
			147 => x"002d025d",
			148 => x"0000025d",
			149 => x"0000025d",
			150 => x"ffbc025d",
			151 => x"0f05d210",
			152 => x"0e032604",
			153 => x"00000281",
			154 => x"09002508",
			155 => x"0c05be04",
			156 => x"00250281",
			157 => x"00000281",
			158 => x"00000281",
			159 => x"ffd90281",
			160 => x"09002710",
			161 => x"0c056304",
			162 => x"000002a5",
			163 => x"0c05be08",
			164 => x"0f05d204",
			165 => x"002a02a5",
			166 => x"000002a5",
			167 => x"000002a5",
			168 => x"000002a5",
			169 => x"0007a908",
			170 => x"09002004",
			171 => x"000002d1",
			172 => x"ff8502d1",
			173 => x"0e032004",
			174 => x"000002d1",
			175 => x"0c05be08",
			176 => x"09002704",
			177 => x"004102d1",
			178 => x"000002d1",
			179 => x"000002d1",
			180 => x"0006ce04",
			181 => x"fe6d02fd",
			182 => x"0100160c",
			183 => x"0f05d208",
			184 => x"0208f004",
			185 => x"016d02fd",
			186 => x"000002fd",
			187 => x"000002fd",
			188 => x"0f058504",
			189 => x"004302fd",
			190 => x"ff3202fd",
			191 => x"0007ca0c",
			192 => x"01001408",
			193 => x"0e033404",
			194 => x"fea50331",
			195 => x"01ba0331",
			196 => x"fe660331",
			197 => x"0208bb04",
			198 => x"01a20331",
			199 => x"041a1404",
			200 => x"fe860331",
			201 => x"02090004",
			202 => x"01e50331",
			203 => x"ff870331",
			204 => x"0007e50c",
			205 => x"09002108",
			206 => x"0303a004",
			207 => x"fe6c036d",
			208 => x"04a3036d",
			209 => x"fe5d036d",
			210 => x"0208dd0c",
			211 => x"0f05b608",
			212 => x"0f059f04",
			213 => x"02e3036d",
			214 => x"01d8036d",
			215 => x"053a036d",
			216 => x"0705be04",
			217 => x"01ca036d",
			218 => x"fe49036d",
			219 => x"0007a908",
			220 => x"09001f04",
			221 => x"000003a1",
			222 => x"fe6803a1",
			223 => x"0f058504",
			224 => x"019703a1",
			225 => x"06014d08",
			226 => x"02091304",
			227 => x"01aa03a1",
			228 => x"000003a1",
			229 => x"0a040504",
			230 => x"fe9903a1",
			231 => x"010c03a1",
			232 => x"0007a908",
			233 => x"09002004",
			234 => x"000003dd",
			235 => x"fe7403dd",
			236 => x"0c059b0c",
			237 => x"0208f708",
			238 => x"0007ba04",
			239 => x"000003dd",
			240 => x"01d603dd",
			241 => x"000003dd",
			242 => x"02089f04",
			243 => x"00c403dd",
			244 => x"06014d04",
			245 => x"000003dd",
			246 => x"ff6803dd",
			247 => x"08053208",
			248 => x"09001f04",
			249 => x"00000411",
			250 => x"fe670411",
			251 => x"0208b404",
			252 => x"01990411",
			253 => x"06014904",
			254 => x"01f50411",
			255 => x"0a040908",
			256 => x"0b05b604",
			257 => x"00000411",
			258 => x"fe820411",
			259 => x"00f30411",
			260 => x"0007ba08",
			261 => x"0f058504",
			262 => x"00000445",
			263 => x"ff590445",
			264 => x"0705d210",
			265 => x"0f05d20c",
			266 => x"09002004",
			267 => x"00000445",
			268 => x"09002604",
			269 => x"004e0445",
			270 => x"00000445",
			271 => x"00000445",
			272 => x"00000445",
			273 => x"0007a908",
			274 => x"09002004",
			275 => x"00000479",
			276 => x"ff7c0479",
			277 => x"0e032004",
			278 => x"00000479",
			279 => x"0c05be0c",
			280 => x"0f05d208",
			281 => x"09002704",
			282 => x"004b0479",
			283 => x"00000479",
			284 => x"00000479",
			285 => x"00000479",
			286 => x"09002714",
			287 => x"0705d210",
			288 => x"0505ea04",
			289 => x"000004a5",
			290 => x"0f05da08",
			291 => x"0b05e904",
			292 => x"005304a5",
			293 => x"000004a5",
			294 => x"000004a5",
			295 => x"000004a5",
			296 => x"ff4604a5",
			297 => x"0f05da14",
			298 => x"0e032004",
			299 => x"000004d1",
			300 => x"0c05be0c",
			301 => x"01001a08",
			302 => x"01001304",
			303 => x"000004d1",
			304 => x"002504d1",
			305 => x"000004d1",
			306 => x"000004d1",
			307 => x"ffc304d1",
			308 => x"0007ca0c",
			309 => x"09002108",
			310 => x"03035304",
			311 => x"fe8d0515",
			312 => x"01dd0515",
			313 => x"fe630515",
			314 => x"0208c70c",
			315 => x"04190f04",
			316 => x"02fa0515",
			317 => x"0007f604",
			318 => x"011b0515",
			319 => x"01e20515",
			320 => x"06014d04",
			321 => x"03630515",
			322 => x"0d066b04",
			323 => x"01070515",
			324 => x"fe550515",
			325 => x"0007e50c",
			326 => x"09002108",
			327 => x"0303a004",
			328 => x"fe700559",
			329 => x"03720559",
			330 => x"fe5e0559",
			331 => x"0208dd10",
			332 => x"0e033e0c",
			333 => x"03040504",
			334 => x"02920559",
			335 => x"0f05ad04",
			336 => x"01a00559",
			337 => x"feba0559",
			338 => x"03900559",
			339 => x"06015304",
			340 => x"01b30559",
			341 => x"fe4d0559",
			342 => x"0007a908",
			343 => x"09002004",
			344 => x"0000059d",
			345 => x"fe73059d",
			346 => x"0c059b0c",
			347 => x"0208f708",
			348 => x"0007ba04",
			349 => x"0000059d",
			350 => x"01e4059d",
			351 => x"0000059d",
			352 => x"02089f04",
			353 => x"00d5059d",
			354 => x"06014d04",
			355 => x"0000059d",
			356 => x"0d066d04",
			357 => x"0000059d",
			358 => x"ff4f059d",
			359 => x"0007ca0c",
			360 => x"09002108",
			361 => x"03035304",
			362 => x"fe9f05e9",
			363 => x"017905e9",
			364 => x"fe6405e9",
			365 => x"0208c710",
			366 => x"04190f04",
			367 => x"02b805e9",
			368 => x"0f058504",
			369 => x"01c905e9",
			370 => x"0007f604",
			371 => x"000005e9",
			372 => x"015b05e9",
			373 => x"06014d04",
			374 => x"02ea05e9",
			375 => x"0d066b04",
			376 => x"00bb05e9",
			377 => x"fe5f05e9",
			378 => x"09002718",
			379 => x"0505ea04",
			380 => x"ff550625",
			381 => x"0208b904",
			382 => x"01910625",
			383 => x"0d06af08",
			384 => x"01001204",
			385 => x"00000625",
			386 => x"ff620625",
			387 => x"0d06b904",
			388 => x"00a40625",
			389 => x"00000625",
			390 => x"0a040c04",
			391 => x"fe6b0625",
			392 => x"00000625",
			393 => x"09002718",
			394 => x"0705d214",
			395 => x"0505ea04",
			396 => x"00000661",
			397 => x"0f05d20c",
			398 => x"01001808",
			399 => x"0208f004",
			400 => x"01090661",
			401 => x"00000661",
			402 => x"00000661",
			403 => x"00000661",
			404 => x"00000661",
			405 => x"0a040c04",
			406 => x"fe8f0661",
			407 => x"00000661",
			408 => x"0900271c",
			409 => x"0505f604",
			410 => x"fef606a5",
			411 => x"0f058504",
			412 => x"01a106a5",
			413 => x"06014d08",
			414 => x"0007f604",
			415 => x"000006a5",
			416 => x"01a906a5",
			417 => x"0705a904",
			418 => x"012f06a5",
			419 => x"0a040204",
			420 => x"fe9f06a5",
			421 => x"000006a5",
			422 => x"0a040c04",
			423 => x"fe6906a5",
			424 => x"000006a5",
			425 => x"0007d80c",
			426 => x"09002108",
			427 => x"0006ce04",
			428 => x"fe7806f9",
			429 => x"01ce06f9",
			430 => x"fe6006f9",
			431 => x"09002518",
			432 => x"0d06af14",
			433 => x"03040508",
			434 => x"0f059f04",
			435 => x"022f06f9",
			436 => x"014a06f9",
			437 => x"06015304",
			438 => x"02dd06f9",
			439 => x"0208d604",
			440 => x"006206f9",
			441 => x"fe5106f9",
			442 => x"049506f9",
			443 => x"0208c904",
			444 => x"014a06f9",
			445 => x"fe6006f9",
			446 => x"09002724",
			447 => x"0007ba10",
			448 => x"0e033408",
			449 => x"09002004",
			450 => x"0000074d",
			451 => x"ffc3074d",
			452 => x"06014204",
			453 => x"0083074d",
			454 => x"0000074d",
			455 => x"06013404",
			456 => x"03ae074d",
			457 => x"0c05b80c",
			458 => x"0007ca04",
			459 => x"0000074d",
			460 => x"0f05da04",
			461 => x"015e074d",
			462 => x"0000074d",
			463 => x"0000074d",
			464 => x"0a040c04",
			465 => x"fe71074d",
			466 => x"0000074d",
			467 => x"0007d814",
			468 => x"01001410",
			469 => x"0e033408",
			470 => x"00075404",
			471 => x"fe7a07a9",
			472 => x"ffe507a9",
			473 => x"0a03cc04",
			474 => x"02b707a9",
			475 => x"ffb007a9",
			476 => x"fe6207a9",
			477 => x"0208f718",
			478 => x"0e034314",
			479 => x"03040508",
			480 => x"0f059f04",
			481 => x"01f607a9",
			482 => x"00d807a9",
			483 => x"00081208",
			484 => x"01001804",
			485 => x"fe8407a9",
			486 => x"000007a9",
			487 => x"00e207a9",
			488 => x"037707a9",
			489 => x"fe8c07a9",
			490 => x"0900272c",
			491 => x"01001720",
			492 => x"0007ca10",
			493 => x"0e033408",
			494 => x"09002004",
			495 => x"0000080d",
			496 => x"ffab080d",
			497 => x"06014504",
			498 => x"00a8080d",
			499 => x"0000080d",
			500 => x"0c05bc0c",
			501 => x"01001608",
			502 => x"02090004",
			503 => x"0178080d",
			504 => x"0000080d",
			505 => x"0000080d",
			506 => x"0000080d",
			507 => x"05069104",
			508 => x"0000080d",
			509 => x"08054204",
			510 => x"04f9080d",
			511 => x"0000080d",
			512 => x"08056f04",
			513 => x"fe6f080d",
			514 => x"0000080d",
			515 => x"0006ce04",
			516 => x"fe8b084b",
			517 => x"0705d218",
			518 => x"09002614",
			519 => x"0f05d210",
			520 => x"0100180c",
			521 => x"0208f008",
			522 => x"0c052e04",
			523 => x"0000084b",
			524 => x"011c084b",
			525 => x"0000084b",
			526 => x"0000084b",
			527 => x"0000084b",
			528 => x"0000084b",
			529 => x"0000084b",
			530 => x"0000084d",
			531 => x"00000851",
			532 => x"00000855",
			533 => x"00000859",
			534 => x"0000085d",
			535 => x"00000861",
			536 => x"00000865",
			537 => x"00000869",
			538 => x"0000086d",
			539 => x"00000871",
			540 => x"00000875",
			541 => x"00000879",
			542 => x"0000087d",
			543 => x"00000881",
			544 => x"00000885",
			545 => x"00000889",
			546 => x"0000088d",
			547 => x"00000891",
			548 => x"00000895",
			549 => x"00000899",
			550 => x"0000089d",
			551 => x"000008a1",
			552 => x"000008a5",
			553 => x"000008a9",
			554 => x"000008ad",
			555 => x"000008b1",
			556 => x"000008b5",
			557 => x"000008b9",
			558 => x"000008bd",
			559 => x"000008c1",
			560 => x"000008c5",
			561 => x"000008c9",
			562 => x"000008cd",
			563 => x"000008d1",
			564 => x"000008d5",
			565 => x"000008d9",
			566 => x"000008dd",
			567 => x"0f05da04",
			568 => x"000008e9",
			569 => x"ffea08e9",
			570 => x"0f058504",
			571 => x"000008f5",
			572 => x"fff408f5",
			573 => x"0007e504",
			574 => x"ffea0901",
			575 => x"00000901",
			576 => x"0007e504",
			577 => x"ffef090d",
			578 => x"0000090d",
			579 => x"0f058504",
			580 => x"00000919",
			581 => x"ffe90919",
			582 => x"0007ba08",
			583 => x"0f058504",
			584 => x"0000092d",
			585 => x"ffe2092d",
			586 => x"0000092d",
			587 => x"0007ba08",
			588 => x"0f055a04",
			589 => x"00000949",
			590 => x"ffa00949",
			591 => x"0e032604",
			592 => x"00000949",
			593 => x"00130949",
			594 => x"0100180c",
			595 => x"0208f008",
			596 => x"0505ea04",
			597 => x"00000965",
			598 => x"007a0965",
			599 => x"00000965",
			600 => x"ff160965",
			601 => x"0007f60c",
			602 => x"0f056704",
			603 => x"00000981",
			604 => x"0a040c04",
			605 => x"ff8a0981",
			606 => x"00000981",
			607 => x"00000981",
			608 => x"0100160c",
			609 => x"0e02bd04",
			610 => x"0000099d",
			611 => x"0f05da04",
			612 => x"000b099d",
			613 => x"0000099d",
			614 => x"0000099d",
			615 => x"0f05da0c",
			616 => x"0c05be08",
			617 => x"0c052804",
			618 => x"000009b9",
			619 => x"002509b9",
			620 => x"000009b9",
			621 => x"000009b9",
			622 => x"0900270c",
			623 => x"0f05da08",
			624 => x"0804a304",
			625 => x"000009d5",
			626 => x"000609d5",
			627 => x"000009d5",
			628 => x"000009d5",
			629 => x"0f05da0c",
			630 => x"07054504",
			631 => x"000009f1",
			632 => x"01001804",
			633 => x"001209f1",
			634 => x"000009f1",
			635 => x"000009f1",
			636 => x"0007ba08",
			637 => x"09002004",
			638 => x"00000a15",
			639 => x"fecc0a15",
			640 => x"0c059b08",
			641 => x"0208f704",
			642 => x"00c10a15",
			643 => x"00000a15",
			644 => x"00000a15",
			645 => x"0f05da10",
			646 => x"06014d0c",
			647 => x"07054504",
			648 => x"00000a39",
			649 => x"09002504",
			650 => x"00920a39",
			651 => x"00000a39",
			652 => x"00000a39",
			653 => x"fef90a39",
			654 => x"0006ce04",
			655 => x"ff3b0a5d",
			656 => x"06014d0c",
			657 => x"09002508",
			658 => x"07057304",
			659 => x"00000a5d",
			660 => x"00810a5d",
			661 => x"00000a5d",
			662 => x"00000a5d",
			663 => x"01001810",
			664 => x"0c05a40c",
			665 => x"07054504",
			666 => x"00000a81",
			667 => x"0f05da04",
			668 => x"00370a81",
			669 => x"00000a81",
			670 => x"00000a81",
			671 => x"ffb00a81",
			672 => x"0f05da10",
			673 => x"0c059b0c",
			674 => x"0705d208",
			675 => x"0c052504",
			676 => x"00000aa5",
			677 => x"00240aa5",
			678 => x"00000aa5",
			679 => x"00000aa5",
			680 => x"ffbe0aa5",
			681 => x"0f05d210",
			682 => x"0e032004",
			683 => x"00000ac9",
			684 => x"0c05be08",
			685 => x"07055d04",
			686 => x"00000ac9",
			687 => x"00180ac9",
			688 => x"00000ac9",
			689 => x"ffdb0ac9",
			690 => x"09002710",
			691 => x"0c056304",
			692 => x"00000aed",
			693 => x"0c05be08",
			694 => x"0f05d204",
			695 => x"00230aed",
			696 => x"00000aed",
			697 => x"00000aed",
			698 => x"00000aed",
			699 => x"0007ba08",
			700 => x"0f055a04",
			701 => x"00000b19",
			702 => x"ff920b19",
			703 => x"0e032604",
			704 => x"00000b19",
			705 => x"0c05be08",
			706 => x"0c057d04",
			707 => x"00000b19",
			708 => x"001f0b19",
			709 => x"00000b19",
			710 => x"09002714",
			711 => x"02087e08",
			712 => x"0505ea04",
			713 => x"00000b45",
			714 => x"00ee0b45",
			715 => x"0705a904",
			716 => x"00060b45",
			717 => x"0d06ad04",
			718 => x"ffe80b45",
			719 => x"00000b45",
			720 => x"feac0b45",
			721 => x"01001610",
			722 => x"0505ea04",
			723 => x"ffb10b79",
			724 => x"0f05b608",
			725 => x"0c05bc04",
			726 => x"017c0b79",
			727 => x"00000b79",
			728 => x"00000b79",
			729 => x"0a03f704",
			730 => x"fe6c0b79",
			731 => x"0f059f04",
			732 => x"00570b79",
			733 => x"00000b79",
			734 => x"0007a908",
			735 => x"09001f04",
			736 => x"00000bad",
			737 => x"fe670bad",
			738 => x"0f058504",
			739 => x"019c0bad",
			740 => x"06014d08",
			741 => x"02091304",
			742 => x"01bc0bad",
			743 => x"00000bad",
			744 => x"0a040504",
			745 => x"fe860bad",
			746 => x"01430bad",
			747 => x"0007ba08",
			748 => x"09002104",
			749 => x"00000be1",
			750 => x"fe780be1",
			751 => x"02089804",
			752 => x"01ba0be1",
			753 => x"0705ba08",
			754 => x"0705b804",
			755 => x"003d0be1",
			756 => x"00000be1",
			757 => x"06014d04",
			758 => x"00000be1",
			759 => x"ff770be1",
			760 => x"01001818",
			761 => x"06014d0c",
			762 => x"0505f604",
			763 => x"00000c1d",
			764 => x"09002504",
			765 => x"01900c1d",
			766 => x"00000c1d",
			767 => x"0a040208",
			768 => x"02087c04",
			769 => x"00000c1d",
			770 => x"ff650c1d",
			771 => x"00a80c1d",
			772 => x"0a040c04",
			773 => x"fe7f0c1d",
			774 => x"00000c1d",
			775 => x"09002714",
			776 => x"0705d210",
			777 => x"0505ea04",
			778 => x"00000c51",
			779 => x"0f05d208",
			780 => x"01001804",
			781 => x"01290c51",
			782 => x"00000c51",
			783 => x"00000c51",
			784 => x"00000c51",
			785 => x"0a040c04",
			786 => x"fe880c51",
			787 => x"00000c51",
			788 => x"08053208",
			789 => x"09002004",
			790 => x"00000c85",
			791 => x"ff6a0c85",
			792 => x"0705d210",
			793 => x"09002004",
			794 => x"00000c85",
			795 => x"0f05d208",
			796 => x"09002604",
			797 => x"00390c85",
			798 => x"00000c85",
			799 => x"00000c85",
			800 => x"00000c85",
			801 => x"0c056308",
			802 => x"08055c04",
			803 => x"ffbf0cb9",
			804 => x"00000cb9",
			805 => x"0705d210",
			806 => x"0900260c",
			807 => x"0c059b08",
			808 => x"0f05ca04",
			809 => x"002b0cb9",
			810 => x"00000cb9",
			811 => x"00000cb9",
			812 => x"00000cb9",
			813 => x"00000cb9",
			814 => x"0006ce04",
			815 => x"ff4f0ce5",
			816 => x"0705d210",
			817 => x"0900260c",
			818 => x"01001808",
			819 => x"0c052e04",
			820 => x"00000ce5",
			821 => x"00720ce5",
			822 => x"00000ce5",
			823 => x"00000ce5",
			824 => x"00000ce5",
			825 => x"0f05da14",
			826 => x"09002610",
			827 => x"0c05bd0c",
			828 => x"0505f604",
			829 => x"00000d11",
			830 => x"01001804",
			831 => x"001b0d11",
			832 => x"00000d11",
			833 => x"00000d11",
			834 => x"00000d11",
			835 => x"00000d11",
			836 => x"0006ce04",
			837 => x"fe6f0d45",
			838 => x"01001610",
			839 => x"0c05be0c",
			840 => x"0f05d208",
			841 => x"0208f004",
			842 => x"01580d45",
			843 => x"00000d45",
			844 => x"00000d45",
			845 => x"00000d45",
			846 => x"0f058504",
			847 => x"00110d45",
			848 => x"ff650d45",
			849 => x"0007e50c",
			850 => x"09002108",
			851 => x"0303a004",
			852 => x"fe750d89",
			853 => x"02c40d89",
			854 => x"fe5f0d89",
			855 => x"0208dd10",
			856 => x"0e033e0c",
			857 => x"03040504",
			858 => x"02580d89",
			859 => x"0f05ad04",
			860 => x"01670d89",
			861 => x"fec90d89",
			862 => x"03410d89",
			863 => x"0705be04",
			864 => x"01770d89",
			865 => x"fe520d89",
			866 => x"0007a908",
			867 => x"01001304",
			868 => x"00000dcd",
			869 => x"fe760dcd",
			870 => x"0c059b0c",
			871 => x"0208f708",
			872 => x"0007ba04",
			873 => x"00000dcd",
			874 => x"01c50dcd",
			875 => x"00000dcd",
			876 => x"02089f04",
			877 => x"00b30dcd",
			878 => x"06014d04",
			879 => x"00000dcd",
			880 => x"0d066d04",
			881 => x"00000dcd",
			882 => x"ff790dcd",
			883 => x"09002718",
			884 => x"0505f604",
			885 => x"ff250e09",
			886 => x"0f058504",
			887 => x"01990e09",
			888 => x"06014d08",
			889 => x"0007f604",
			890 => x"00000e09",
			891 => x"017d0e09",
			892 => x"0705a904",
			893 => x"01030e09",
			894 => x"fed50e09",
			895 => x"0a040c04",
			896 => x"fe6a0e09",
			897 => x"00000e09",
			898 => x"0007ca18",
			899 => x"09002114",
			900 => x"06012108",
			901 => x"0f050304",
			902 => x"00000e55",
			903 => x"025d0e55",
			904 => x"01001208",
			905 => x"09001f04",
			906 => x"00350e55",
			907 => x"00000e55",
			908 => x"fe930e55",
			909 => x"fe650e55",
			910 => x"0208bb04",
			911 => x"01ae0e55",
			912 => x"06014a04",
			913 => x"02420e55",
			914 => x"041a5004",
			915 => x"fe720e55",
			916 => x"00000e55",
			917 => x"0006ce04",
			918 => x"feb20e99",
			919 => x"06014d0c",
			920 => x"09002508",
			921 => x"07057304",
			922 => x"00000e99",
			923 => x"01000e99",
			924 => x"00000e99",
			925 => x"0705a908",
			926 => x"0303f504",
			927 => x"00480e99",
			928 => x"00000e99",
			929 => x"06016008",
			930 => x"0303e504",
			931 => x"00000e99",
			932 => x"ffe20e99",
			933 => x"00000e99",
			934 => x"0900271c",
			935 => x"0505f604",
			936 => x"ff0c0edd",
			937 => x"0f058504",
			938 => x"019d0edd",
			939 => x"06014d08",
			940 => x"0007f604",
			941 => x"00000edd",
			942 => x"01920edd",
			943 => x"0705a904",
			944 => x"011b0edd",
			945 => x"0a040204",
			946 => x"fead0edd",
			947 => x"00000edd",
			948 => x"0a040c04",
			949 => x"fe690edd",
			950 => x"00000edd",
			951 => x"0007d814",
			952 => x"01001410",
			953 => x"0e033408",
			954 => x"00075404",
			955 => x"fe760f31",
			956 => x"ffdb0f31",
			957 => x"0a03cc04",
			958 => x"03140f31",
			959 => x"ff970f31",
			960 => x"fe610f31",
			961 => x"0208f714",
			962 => x"0e034310",
			963 => x"0208bb04",
			964 => x"020e0f31",
			965 => x"06015204",
			966 => x"02b70f31",
			967 => x"0b05c704",
			968 => x"01020f31",
			969 => x"fe3f0f31",
			970 => x"03b90f31",
			971 => x"fe840f31",
			972 => x"0007e514",
			973 => x"09002108",
			974 => x"00075404",
			975 => x"fe640f8d",
			976 => x"0b0a0f8d",
			977 => x"0a03fc04",
			978 => x"fe5a0f8d",
			979 => x"08052e04",
			980 => x"fe950f8d",
			981 => x"02530f8d",
			982 => x"0208f718",
			983 => x"0f05ca14",
			984 => x"0c05b80c",
			985 => x"0f05ad08",
			986 => x"0f059f04",
			987 => x"04270f8d",
			988 => x"02bc0f8d",
			989 => x"09e20f8d",
			990 => x"0208b904",
			991 => x"03fa0f8d",
			992 => x"fe6d0f8d",
			993 => x"09a10f8d",
			994 => x"fe6f0f8d",
			995 => x"0007ca0c",
			996 => x"09002108",
			997 => x"03035304",
			998 => x"fe950fe1",
			999 => x"01a70fe1",
			1000 => x"fe630fe1",
			1001 => x"0208f01c",
			1002 => x"0c05b814",
			1003 => x"09002710",
			1004 => x"0f05ad08",
			1005 => x"0208bb04",
			1006 => x"01d50fe1",
			1007 => x"001e0fe1",
			1008 => x"08055c04",
			1009 => x"067c0fe1",
			1010 => x"02720fe1",
			1011 => x"feca0fe1",
			1012 => x"0208b904",
			1013 => x"01840fe1",
			1014 => x"fe640fe1",
			1015 => x"fe860fe1",
			1016 => x"0008122c",
			1017 => x"0007e51c",
			1018 => x"09001f08",
			1019 => x"0a036304",
			1020 => x"c9c51045",
			1021 => x"dd161045",
			1022 => x"09002108",
			1023 => x"0a036304",
			1024 => x"c9b81045",
			1025 => x"d53c1045",
			1026 => x"0a03fc04",
			1027 => x"c9a61045",
			1028 => x"0a040504",
			1029 => x"cc6a1045",
			1030 => x"c9e11045",
			1031 => x"0208ad04",
			1032 => x"f4841045",
			1033 => x"0c059b04",
			1034 => x"d7291045",
			1035 => x"0208c904",
			1036 => x"cd621045",
			1037 => x"c9b81045",
			1038 => x"0f05b604",
			1039 => x"f63b1045",
			1040 => x"d53c1045",
			1041 => x"0007ca0c",
			1042 => x"09002108",
			1043 => x"03033b04",
			1044 => x"feac109b",
			1045 => x"017a109b",
			1046 => x"fe64109b",
			1047 => x"0f05d21c",
			1048 => x"09002718",
			1049 => x"0007cf04",
			1050 => x"04d0109b",
			1051 => x"0007f608",
			1052 => x"0208ad04",
			1053 => x"01da109b",
			1054 => x"fe99109b",
			1055 => x"0d06ad08",
			1056 => x"0d067704",
			1057 => x"01c8109b",
			1058 => x"010c109b",
			1059 => x"02d0109b",
			1060 => x"ff67109b",
			1061 => x"fe9a109b",
			1062 => x"0000109d",
			1063 => x"000010a1",
			1064 => x"000010a5",
			1065 => x"000010a9",
			1066 => x"000010ad",
			1067 => x"000010b1",
			1068 => x"000010b5",
			1069 => x"000010b9",
			1070 => x"000010bd",
			1071 => x"000010c1",
			1072 => x"000010c5",
			1073 => x"000010c9",
			1074 => x"000010cd",
			1075 => x"000010d1",
			1076 => x"000010d5",
			1077 => x"000010d9",
			1078 => x"000010dd",
			1079 => x"000010e1",
			1080 => x"000010e5",
			1081 => x"000010e9",
			1082 => x"000010ed",
			1083 => x"000010f1",
			1084 => x"000010f5",
			1085 => x"000010f9",
			1086 => x"000010fd",
			1087 => x"00001101",
			1088 => x"00001105",
			1089 => x"00001109",
			1090 => x"0000110d",
			1091 => x"00001111",
			1092 => x"00001115",
			1093 => x"00001119",
			1094 => x"0000111d",
			1095 => x"00001121",
			1096 => x"00001125",
			1097 => x"00001129",
			1098 => x"0000112d",
			1099 => x"0f05da04",
			1100 => x"00001139",
			1101 => x"ffec1139",
			1102 => x"0f058504",
			1103 => x"00001145",
			1104 => x"ffff1145",
			1105 => x"0007e504",
			1106 => x"ffed1151",
			1107 => x"00001151",
			1108 => x"0f058504",
			1109 => x"0000115d",
			1110 => x"ffec115d",
			1111 => x"00075404",
			1112 => x"fef21171",
			1113 => x"02087e04",
			1114 => x"006f1171",
			1115 => x"00001171",
			1116 => x"0f058504",
			1117 => x"00001185",
			1118 => x"09001f04",
			1119 => x"00001185",
			1120 => x"ffd81185",
			1121 => x"0006ce04",
			1122 => x"fe9c11a1",
			1123 => x"02089008",
			1124 => x"09002704",
			1125 => x"011111a1",
			1126 => x"000011a1",
			1127 => x"000011a1",
			1128 => x"0100180c",
			1129 => x"0505ea04",
			1130 => x"000011bd",
			1131 => x"06014d04",
			1132 => x"008811bd",
			1133 => x"000011bd",
			1134 => x"ff2911bd",
			1135 => x"0007f60c",
			1136 => x"0f056704",
			1137 => x"000011d9",
			1138 => x"0a040c04",
			1139 => x"ff9211d9",
			1140 => x"000011d9",
			1141 => x"000011d9",
			1142 => x"0100160c",
			1143 => x"0415f304",
			1144 => x"000011f5",
			1145 => x"0f05da04",
			1146 => x"000911f5",
			1147 => x"000011f5",
			1148 => x"000011f5",
			1149 => x"0f05da0c",
			1150 => x"0c05be08",
			1151 => x"0c052804",
			1152 => x"00001211",
			1153 => x"00221211",
			1154 => x"00001211",
			1155 => x"00001211",
			1156 => x"0900270c",
			1157 => x"0f05da08",
			1158 => x"0006ce04",
			1159 => x"0000122d",
			1160 => x"0006122d",
			1161 => x"0000122d",
			1162 => x"0000122d",
			1163 => x"0900270c",
			1164 => x"02089008",
			1165 => x"0505f604",
			1166 => x"00001251",
			1167 => x"01211251",
			1168 => x"00001251",
			1169 => x"0a040c04",
			1170 => x"fe971251",
			1171 => x"00001251",
			1172 => x"0007ba08",
			1173 => x"0f055a04",
			1174 => x"00001275",
			1175 => x"fed41275",
			1176 => x"0c059b08",
			1177 => x"0208f704",
			1178 => x"00b01275",
			1179 => x"00001275",
			1180 => x"00001275",
			1181 => x"0f05da10",
			1182 => x"06014d0c",
			1183 => x"0c052504",
			1184 => x"00001299",
			1185 => x"09002504",
			1186 => x"00891299",
			1187 => x"00001299",
			1188 => x"00001299",
			1189 => x"ff021299",
			1190 => x"0f05da10",
			1191 => x"0705d20c",
			1192 => x"0c052504",
			1193 => x"000012bd",
			1194 => x"09002604",
			1195 => x"006a12bd",
			1196 => x"000012bd",
			1197 => x"000012bd",
			1198 => x"ff5912bd",
			1199 => x"01001810",
			1200 => x"0c05a40c",
			1201 => x"0505ea04",
			1202 => x"000012e1",
			1203 => x"0f05da04",
			1204 => x"003212e1",
			1205 => x"000012e1",
			1206 => x"000012e1",
			1207 => x"ffb612e1",
			1208 => x"0f05da10",
			1209 => x"0e032004",
			1210 => x"00001305",
			1211 => x"09002708",
			1212 => x"0c05be04",
			1213 => x"00221305",
			1214 => x"00001305",
			1215 => x"00001305",
			1216 => x"ffc81305",
			1217 => x"0f05d210",
			1218 => x"0e032004",
			1219 => x"00001329",
			1220 => x"0c05be08",
			1221 => x"07055d04",
			1222 => x"00001329",
			1223 => x"00151329",
			1224 => x"00001329",
			1225 => x"ffde1329",
			1226 => x"0007ba08",
			1227 => x"09002104",
			1228 => x"00001355",
			1229 => x"fe7d1355",
			1230 => x"02089804",
			1231 => x"01951355",
			1232 => x"05065f04",
			1233 => x"00221355",
			1234 => x"03042604",
			1235 => x"ffbd1355",
			1236 => x"00001355",
			1237 => x"0c056308",
			1238 => x"08055c04",
			1239 => x"ffc41381",
			1240 => x"00001381",
			1241 => x"0705d20c",
			1242 => x"09002608",
			1243 => x"0c059b04",
			1244 => x"00261381",
			1245 => x"00001381",
			1246 => x"00001381",
			1247 => x"00001381",
			1248 => x"0417c304",
			1249 => x"fee913ad",
			1250 => x"06014d08",
			1251 => x"09002504",
			1252 => x"007c13ad",
			1253 => x"000013ad",
			1254 => x"02087e04",
			1255 => x"000013ad",
			1256 => x"0f057204",
			1257 => x"000013ad",
			1258 => x"ffe013ad",
			1259 => x"09002514",
			1260 => x"06014d08",
			1261 => x"00076604",
			1262 => x"000013e1",
			1263 => x"008413e1",
			1264 => x"0f057204",
			1265 => x"000013e1",
			1266 => x"00083c04",
			1267 => x"ffe013e1",
			1268 => x"000013e1",
			1269 => x"0f058504",
			1270 => x"000013e1",
			1271 => x"fede13e1",
			1272 => x"0007a908",
			1273 => x"09001f04",
			1274 => x"00001415",
			1275 => x"fe681415",
			1276 => x"0f058504",
			1277 => x"01991415",
			1278 => x"06014d08",
			1279 => x"02091304",
			1280 => x"01b41415",
			1281 => x"00001415",
			1282 => x"0705a904",
			1283 => x"01581415",
			1284 => x"fea11415",
			1285 => x"08053208",
			1286 => x"01001204",
			1287 => x"00001449",
			1288 => x"fe7a1449",
			1289 => x"02089804",
			1290 => x"01a61449",
			1291 => x"0705ba08",
			1292 => x"0c059d04",
			1293 => x"002c1449",
			1294 => x"00001449",
			1295 => x"06014d04",
			1296 => x"00001449",
			1297 => x"ff7c1449",
			1298 => x"01001818",
			1299 => x"06014d0c",
			1300 => x"0505f604",
			1301 => x"00001485",
			1302 => x"09002504",
			1303 => x"016f1485",
			1304 => x"00001485",
			1305 => x"0a040208",
			1306 => x"02087c04",
			1307 => x"00001485",
			1308 => x"ff7e1485",
			1309 => x"00841485",
			1310 => x"0a040c04",
			1311 => x"fe851485",
			1312 => x"00001485",
			1313 => x"0f05da18",
			1314 => x"06014d0c",
			1315 => x"07055d04",
			1316 => x"000014b9",
			1317 => x"09002504",
			1318 => x"00e814b9",
			1319 => x"000014b9",
			1320 => x"0705a908",
			1321 => x"05065f04",
			1322 => x"002114b9",
			1323 => x"000014b9",
			1324 => x"000014b9",
			1325 => x"fec014b9",
			1326 => x"0007ba08",
			1327 => x"0f058504",
			1328 => x"000014ed",
			1329 => x"ff6a14ed",
			1330 => x"01001504",
			1331 => x"000014ed",
			1332 => x"0f05d20c",
			1333 => x"09002608",
			1334 => x"01001804",
			1335 => x"003814ed",
			1336 => x"000014ed",
			1337 => x"000014ed",
			1338 => x"000014ed",
			1339 => x"0006ce04",
			1340 => x"feb91519",
			1341 => x"0c059b10",
			1342 => x"0208f70c",
			1343 => x"09002608",
			1344 => x"0705d204",
			1345 => x"00da1519",
			1346 => x"00001519",
			1347 => x"00001519",
			1348 => x"00001519",
			1349 => x"00001519",
			1350 => x"08051304",
			1351 => x"ff821545",
			1352 => x"0e032004",
			1353 => x"00001545",
			1354 => x"08052704",
			1355 => x"00001545",
			1356 => x"0c05be08",
			1357 => x"0f05d204",
			1358 => x"00521545",
			1359 => x"00001545",
			1360 => x"00001545",
			1361 => x"0f05da14",
			1362 => x"09002610",
			1363 => x"0c05bd0c",
			1364 => x"0505f604",
			1365 => x"00001571",
			1366 => x"01001804",
			1367 => x"00181571",
			1368 => x"00001571",
			1369 => x"00001571",
			1370 => x"00001571",
			1371 => x"00001571",
			1372 => x"09002718",
			1373 => x"02087e08",
			1374 => x"0505ea04",
			1375 => x"000015a5",
			1376 => x"00fd15a5",
			1377 => x"0f05ad04",
			1378 => x"000015a5",
			1379 => x"0f05da08",
			1380 => x"0705ea04",
			1381 => x"002e15a5",
			1382 => x"000015a5",
			1383 => x"000015a5",
			1384 => x"fea715a5",
			1385 => x"0007ba0c",
			1386 => x"09002108",
			1387 => x"0804a304",
			1388 => x"ff4015f1",
			1389 => x"000015f1",
			1390 => x"fe6715f1",
			1391 => x"0d06770c",
			1392 => x"09002708",
			1393 => x"0b05d804",
			1394 => x"01ae15f1",
			1395 => x"001f15f1",
			1396 => x"000015f1",
			1397 => x"06014d08",
			1398 => x"02091304",
			1399 => x"01b615f1",
			1400 => x"000015f1",
			1401 => x"02089f04",
			1402 => x"015f15f1",
			1403 => x"fe7a15f1",
			1404 => x"0900271c",
			1405 => x"0e03200c",
			1406 => x"00082608",
			1407 => x"09001f04",
			1408 => x"00001635",
			1409 => x"ffa31635",
			1410 => x"00921635",
			1411 => x"0208f00c",
			1412 => x"0c05be08",
			1413 => x"01001804",
			1414 => x"01661635",
			1415 => x"00001635",
			1416 => x"00001635",
			1417 => x"00001635",
			1418 => x"0a040c04",
			1419 => x"fe821635",
			1420 => x"00001635",
			1421 => x"09002718",
			1422 => x"07055d04",
			1423 => x"ff3a1671",
			1424 => x"0208b904",
			1425 => x"019a1671",
			1426 => x"0d06af08",
			1427 => x"01001204",
			1428 => x"00001671",
			1429 => x"ff4c1671",
			1430 => x"0d06b904",
			1431 => x"00b11671",
			1432 => x"00001671",
			1433 => x"0a040c04",
			1434 => x"fe6b1671",
			1435 => x"00001671",
			1436 => x"0007ca18",
			1437 => x"09002114",
			1438 => x"06012108",
			1439 => x"0f050304",
			1440 => x"000016bd",
			1441 => x"020316bd",
			1442 => x"01001208",
			1443 => x"09001f04",
			1444 => x"002716bd",
			1445 => x"000016bd",
			1446 => x"fea616bd",
			1447 => x"fe6616bd",
			1448 => x"0208bb04",
			1449 => x"01a816bd",
			1450 => x"06014a04",
			1451 => x"022416bd",
			1452 => x"041a5004",
			1453 => x"fe7a16bd",
			1454 => x"000016bd",
			1455 => x"0006ce04",
			1456 => x"fe6e16f9",
			1457 => x"01001614",
			1458 => x"0c05be10",
			1459 => x"0f05d20c",
			1460 => x"0007ba08",
			1461 => x"00078b04",
			1462 => x"009e16f9",
			1463 => x"000016f9",
			1464 => x"017c16f9",
			1465 => x"000016f9",
			1466 => x"000016f9",
			1467 => x"0f058504",
			1468 => x"002916f9",
			1469 => x"ff4b16f9",
			1470 => x"0415f304",
			1471 => x"fe72173d",
			1472 => x"02087e0c",
			1473 => x"03037b04",
			1474 => x"0000173d",
			1475 => x"09002804",
			1476 => x"01f0173d",
			1477 => x"0000173d",
			1478 => x"08054e04",
			1479 => x"ff97173d",
			1480 => x"0100160c",
			1481 => x"0c05a408",
			1482 => x"0208f704",
			1483 => x"012c173d",
			1484 => x"0000173d",
			1485 => x"0000173d",
			1486 => x"0000173d",
			1487 => x"0007ba0c",
			1488 => x"09002108",
			1489 => x"0f052f04",
			1490 => x"ff241791",
			1491 => x"00001791",
			1492 => x"fe661791",
			1493 => x"0d067708",
			1494 => x"09002704",
			1495 => x"01af1791",
			1496 => x"00001791",
			1497 => x"02089f04",
			1498 => x"018a1791",
			1499 => x"041a320c",
			1500 => x"0e037004",
			1501 => x"fe721791",
			1502 => x"0d06c504",
			1503 => x"003d1791",
			1504 => x"00001791",
			1505 => x"02091104",
			1506 => x"01ca1791",
			1507 => x"00001791",
			1508 => x"0007ca0c",
			1509 => x"09002108",
			1510 => x"03033b04",
			1511 => x"feb917f5",
			1512 => x"015217f5",
			1513 => x"fe6517f5",
			1514 => x"0208d61c",
			1515 => x"0c05b810",
			1516 => x"0f05ad0c",
			1517 => x"0f058504",
			1518 => x"01ba17f5",
			1519 => x"0d067704",
			1520 => x"016617f5",
			1521 => x"000017f5",
			1522 => x"030117f5",
			1523 => x"02089f04",
			1524 => x"016e17f5",
			1525 => x"0b05e804",
			1526 => x"009717f5",
			1527 => x"ff0617f5",
			1528 => x"0705cf08",
			1529 => x"09002504",
			1530 => x"027017f5",
			1531 => x"feec17f5",
			1532 => x"fe7817f5",
			1533 => x"09002724",
			1534 => x"02087e08",
			1535 => x"0505ea04",
			1536 => x"00001841",
			1537 => x"010b1841",
			1538 => x"0f05ad0c",
			1539 => x"06014e04",
			1540 => x"00001841",
			1541 => x"0a040204",
			1542 => x"ffd51841",
			1543 => x"00001841",
			1544 => x"0a03e304",
			1545 => x"00001841",
			1546 => x"0f05da08",
			1547 => x"0705ea04",
			1548 => x"00401841",
			1549 => x"00001841",
			1550 => x"00001841",
			1551 => x"fea11841",
			1552 => x"0007d818",
			1553 => x"0100140c",
			1554 => x"00075404",
			1555 => x"fe6418ad",
			1556 => x"0a03d104",
			1557 => x"057518ad",
			1558 => x"fec518ad",
			1559 => x"0a03fc04",
			1560 => x"fe5b18ad",
			1561 => x"08052e04",
			1562 => x"fe9f18ad",
			1563 => x"01f718ad",
			1564 => x"0208f71c",
			1565 => x"0c05ba14",
			1566 => x"0e034a10",
			1567 => x"03041d0c",
			1568 => x"0f05b608",
			1569 => x"0f059f04",
			1570 => x"035e18ad",
			1571 => x"015a18ad",
			1572 => x"06c118ad",
			1573 => x"00a818ad",
			1574 => x"05cc18ad",
			1575 => x"0208c904",
			1576 => x"02d718ad",
			1577 => x"fe7418ad",
			1578 => x"fe6e18ad",
			1579 => x"0007ca0c",
			1580 => x"09002108",
			1581 => x"03033b04",
			1582 => x"fec81923",
			1583 => x"012e1923",
			1584 => x"fe651923",
			1585 => x"0f05d22c",
			1586 => x"0c05b81c",
			1587 => x"01001610",
			1588 => x"0e03430c",
			1589 => x"0303f504",
			1590 => x"01b91923",
			1591 => x"03040e04",
			1592 => x"00e11923",
			1593 => x"00001923",
			1594 => x"029a1923",
			1595 => x"0303f504",
			1596 => x"01911923",
			1597 => x"04196d04",
			1598 => x"00001923",
			1599 => x"fea61923",
			1600 => x"06015204",
			1601 => x"018e1923",
			1602 => x"06015f08",
			1603 => x"0b05d804",
			1604 => x"00001923",
			1605 => x"fe9d1923",
			1606 => x"00001923",
			1607 => x"feb11923",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(530, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(1062, initial_addr_3'length));
	end generate gen_rom_0;

	gen_rom_1: if SELECT_ROM = 1 generate
		bank <= (
			0 => x"00000005",
			1 => x"00000009",
			2 => x"0000000d",
			3 => x"00000011",
			4 => x"00000015",
			5 => x"00000019",
			6 => x"0000001d",
			7 => x"00000021",
			8 => x"00000025",
			9 => x"00000029",
			10 => x"0000002d",
			11 => x"00000031",
			12 => x"00000035",
			13 => x"00000039",
			14 => x"0000003d",
			15 => x"00000041",
			16 => x"00000045",
			17 => x"00000049",
			18 => x"0000004d",
			19 => x"00000051",
			20 => x"00000055",
			21 => x"00000059",
			22 => x"0000005d",
			23 => x"00000061",
			24 => x"00000065",
			25 => x"00000069",
			26 => x"0000006d",
			27 => x"00000071",
			28 => x"00000075",
			29 => x"00000079",
			30 => x"0000007d",
			31 => x"00000081",
			32 => x"00000085",
			33 => x"00000089",
			34 => x"0000008d",
			35 => x"00000091",
			36 => x"00000095",
			37 => x"00000099",
			38 => x"0705a404",
			39 => x"ff3700a5",
			40 => x"000000a5",
			41 => x"040e6304",
			42 => x"ffa400b1",
			43 => x"000000b1",
			44 => x"01004504",
			45 => x"000000bd",
			46 => x"ffa900bd",
			47 => x"09004f04",
			48 => x"000000c9",
			49 => x"ffd100c9",
			50 => x"09003904",
			51 => x"000000d5",
			52 => x"ffdd00d5",
			53 => x"0705a404",
			54 => x"ffe500e1",
			55 => x"000000e1",
			56 => x"05064108",
			57 => x"04192604",
			58 => x"ff2d00f5",
			59 => x"000000f5",
			60 => x"000000f5",
			61 => x"01003608",
			62 => x"02087e04",
			63 => x"00000109",
			64 => x"00060109",
			65 => x"ff590109",
			66 => x"0705d208",
			67 => x"02091904",
			68 => x"ffef011d",
			69 => x"0000011d",
			70 => x"0000011d",
			71 => x"0b056508",
			72 => x"0e032004",
			73 => x"00000139",
			74 => x"ff810139",
			75 => x"06016004",
			76 => x"00070139",
			77 => x"00000139",
			78 => x"09004f08",
			79 => x"0007f604",
			80 => x"00120155",
			81 => x"00000155",
			82 => x"04116204",
			83 => x"ffd20155",
			84 => x"00000155",
			85 => x"0b056504",
			86 => x"ff8e0171",
			87 => x"06016308",
			88 => x"06014904",
			89 => x"00000171",
			90 => x"002b0171",
			91 => x"00000171",
			92 => x"0705a404",
			93 => x"ff9e018d",
			94 => x"02087e04",
			95 => x"0000018d",
			96 => x"020a2004",
			97 => x"002b018d",
			98 => x"0000018d",
			99 => x"0d06770c",
			100 => x"0c059b08",
			101 => x"0b05d604",
			102 => x"ffe001a9",
			103 => x"000001a9",
			104 => x"000001a9",
			105 => x"000001a9",
			106 => x"07056108",
			107 => x"04192604",
			108 => x"ff2001cd",
			109 => x"000001cd",
			110 => x"06016308",
			111 => x"06014904",
			112 => x"000001cd",
			113 => x"003501cd",
			114 => x"000001cd",
			115 => x"040e6304",
			116 => x"fee601f1",
			117 => x"0f05da04",
			118 => x"000001f1",
			119 => x"0c050704",
			120 => x"000001f1",
			121 => x"01007304",
			122 => x"009601f1",
			123 => x"000001f1",
			124 => x"0208a404",
			125 => x"ffd90215",
			126 => x"0100470c",
			127 => x"09001f04",
			128 => x"00000215",
			129 => x"0e030004",
			130 => x"00000215",
			131 => x"001b0215",
			132 => x"00000215",
			133 => x"0705a904",
			134 => x"ffcc0239",
			135 => x"0100790c",
			136 => x"09001f04",
			137 => x"00000239",
			138 => x"0d065104",
			139 => x"00000239",
			140 => x"00170239",
			141 => x"00000239",
			142 => x"07056108",
			143 => x"0418f304",
			144 => x"fec90265",
			145 => x"00000265",
			146 => x"0100710c",
			147 => x"0f059f04",
			148 => x"00000265",
			149 => x"08056f04",
			150 => x"00ab0265",
			151 => x"00000265",
			152 => x"00000265",
			153 => x"01004514",
			154 => x"0f05c308",
			155 => x"06014d04",
			156 => x"ffeb0291",
			157 => x"00000291",
			158 => x"0c050b04",
			159 => x"00000291",
			160 => x"01001304",
			161 => x"00000291",
			162 => x"006b0291",
			163 => x"fef40291",
			164 => x"04116204",
			165 => x"feb802bd",
			166 => x"06014904",
			167 => x"000002bd",
			168 => x"0008260c",
			169 => x"0f070f08",
			170 => x"0f057204",
			171 => x"000002bd",
			172 => x"00dd02bd",
			173 => x"000002bd",
			174 => x"000002bd",
			175 => x"01004518",
			176 => x"0f05c308",
			177 => x"06014d04",
			178 => x"fff502f1",
			179 => x"000002f1",
			180 => x"02085404",
			181 => x"000002f1",
			182 => x"0303e504",
			183 => x"000002f1",
			184 => x"00049c04",
			185 => x"000002f1",
			186 => x"005c02f1",
			187 => x"fefd02f1",
			188 => x"09005d1c",
			189 => x"0d06470c",
			190 => x"03041d08",
			191 => x"0b05b804",
			192 => x"ff63032d",
			193 => x"0000032d",
			194 => x"0000032d",
			195 => x"02087e04",
			196 => x"0000032d",
			197 => x"041a3208",
			198 => x"09001f04",
			199 => x"0000032d",
			200 => x"010a032d",
			201 => x"0000032d",
			202 => x"fe8f032d",
			203 => x"0100451c",
			204 => x"0c059b10",
			205 => x"03052b0c",
			206 => x"0705d208",
			207 => x"0b05e904",
			208 => x"ff950369",
			209 => x"00000369",
			210 => x"00000369",
			211 => x"00000369",
			212 => x"02089804",
			213 => x"00000369",
			214 => x"041a5004",
			215 => x"00b40369",
			216 => x"00000369",
			217 => x"feae0369",
			218 => x"0415af18",
			219 => x"0413e90c",
			220 => x"09005d08",
			221 => x"09004604",
			222 => x"fe7703cd",
			223 => x"feda03cd",
			224 => x"fe5503cd",
			225 => x"05066a04",
			226 => x"fe5703cd",
			227 => x"02112d04",
			228 => x"037d03cd",
			229 => x"fe6b03cd",
			230 => x"0f05850c",
			231 => x"09002504",
			232 => x"fe5a03cd",
			233 => x"0c056304",
			234 => x"fe9e03cd",
			235 => x"037103cd",
			236 => x"09001f08",
			237 => x"00083104",
			238 => x"ffcd03cd",
			239 => x"feeb03cd",
			240 => x"0303f504",
			241 => x"028c03cd",
			242 => x"038903cd",
			243 => x"04116204",
			244 => x"feb10401",
			245 => x"02087e04",
			246 => x"00000401",
			247 => x"041a3210",
			248 => x"0f07570c",
			249 => x"09001f04",
			250 => x"00000401",
			251 => x"0505df04",
			252 => x"00000401",
			253 => x"01020401",
			254 => x"00000401",
			255 => x"00000401",
			256 => x"040e6304",
			257 => x"fe810445",
			258 => x"0c059b0c",
			259 => x"0004a004",
			260 => x"00000445",
			261 => x"06014504",
			262 => x"ff730445",
			263 => x"00000445",
			264 => x"06016310",
			265 => x"0008120c",
			266 => x"0f058504",
			267 => x"00000445",
			268 => x"020a4604",
			269 => x"011e0445",
			270 => x"00000445",
			271 => x"00000445",
			272 => x"00000445",
			273 => x"0415af18",
			274 => x"040e6304",
			275 => x"fe6704a9",
			276 => x"0a030d0c",
			277 => x"0c054504",
			278 => x"fee204a9",
			279 => x"0f082204",
			280 => x"01f604a9",
			281 => x"ffb504a9",
			282 => x"0414ff04",
			283 => x"fe9b04a9",
			284 => x"ffee04a9",
			285 => x"0007f60c",
			286 => x"0303e504",
			287 => x"ff4204a9",
			288 => x"0f058504",
			289 => x"000004a9",
			290 => x"019904a9",
			291 => x"06014e04",
			292 => x"fe7b04a9",
			293 => x"0a040c08",
			294 => x"0208ad04",
			295 => x"000004a9",
			296 => x"017d04a9",
			297 => x"fee704a9",
			298 => x"0415af18",
			299 => x"01003614",
			300 => x"01001a08",
			301 => x"0a030404",
			302 => x"00000515",
			303 => x"fed50515",
			304 => x"0a032104",
			305 => x"ffb50515",
			306 => x"01001d04",
			307 => x"00000515",
			308 => x"004c0515",
			309 => x"fe680515",
			310 => x"02089310",
			311 => x"0007c20c",
			312 => x"0a037208",
			313 => x"0a036304",
			314 => x"ff860515",
			315 => x"00000515",
			316 => x"00a70515",
			317 => x"fe7f0515",
			318 => x"0303e504",
			319 => x"ff8b0515",
			320 => x"041a3204",
			321 => x"01920515",
			322 => x"0f05b604",
			323 => x"ff970515",
			324 => x"00650515",
			325 => x"09003928",
			326 => x"02087c0c",
			327 => x"09002808",
			328 => x"01001a04",
			329 => x"fe7a0579",
			330 => x"00000579",
			331 => x"00000579",
			332 => x"01001614",
			333 => x"06014908",
			334 => x"0007e504",
			335 => x"00000579",
			336 => x"fed80579",
			337 => x"0705a304",
			338 => x"ff570579",
			339 => x"00082604",
			340 => x"012d0579",
			341 => x"00000579",
			342 => x"0505df04",
			343 => x"00000579",
			344 => x"01800579",
			345 => x"0006f108",
			346 => x"01002104",
			347 => x"00000579",
			348 => x"fe750579",
			349 => x"00000579",
			350 => x"040e6304",
			351 => x"fe6b05c5",
			352 => x"07056108",
			353 => x"0416b604",
			354 => x"fe7205c5",
			355 => x"000005c5",
			356 => x"06016314",
			357 => x"0007e508",
			358 => x"02085204",
			359 => x"000005c5",
			360 => x"019705c5",
			361 => x"06014e04",
			362 => x"feae05c5",
			363 => x"0208ad04",
			364 => x"000005c5",
			365 => x"012c05c5",
			366 => x"04195404",
			367 => x"ff0505c5",
			368 => x"000005c5",
			369 => x"040e6304",
			370 => x"fe760609",
			371 => x"0d060304",
			372 => x"ff030609",
			373 => x"09002514",
			374 => x"06014d08",
			375 => x"0007a904",
			376 => x"00000609",
			377 => x"fef50609",
			378 => x"02087e04",
			379 => x"00000609",
			380 => x"00084404",
			381 => x"00d10609",
			382 => x"00000609",
			383 => x"0900a804",
			384 => x"01590609",
			385 => x"ffd30609",
			386 => x"0415af10",
			387 => x"0100360c",
			388 => x"0505f904",
			389 => x"fe64065d",
			390 => x"00062204",
			391 => x"03e7065d",
			392 => x"01b1065d",
			393 => x"fe62065d",
			394 => x"0303e504",
			395 => x"fe64065d",
			396 => x"0a040c14",
			397 => x"09001e04",
			398 => x"fe6e065d",
			399 => x"02085b04",
			400 => x"ff7e065d",
			401 => x"041a5008",
			402 => x"01002304",
			403 => x"01e7065d",
			404 => x"0124065d",
			405 => x"005b065d",
			406 => x"fe7d065d",
			407 => x"00069710",
			408 => x"0100450c",
			409 => x"0505f904",
			410 => x"fe6906c1",
			411 => x"0e03e704",
			412 => x"017506c1",
			413 => x"02fc06c1",
			414 => x"fe6406c1",
			415 => x"0303e504",
			416 => x"fe7506c1",
			417 => x"0900210c",
			418 => x"06014e04",
			419 => x"fe2506c1",
			420 => x"0a03fd04",
			421 => x"01d206c1",
			422 => x"ffee06c1",
			423 => x"0008120c",
			424 => x"0100bc08",
			425 => x"02086e04",
			426 => x"002306c1",
			427 => x"01b006c1",
			428 => x"ff6206c1",
			429 => x"06015704",
			430 => x"feab06c1",
			431 => x"015006c1",
			432 => x"09003924",
			433 => x"0f05d21c",
			434 => x"06014908",
			435 => x"09002604",
			436 => x"ff3f0725",
			437 => x"00000725",
			438 => x"06016310",
			439 => x"0008260c",
			440 => x"02087c04",
			441 => x"00000725",
			442 => x"03043504",
			443 => x"00ce0725",
			444 => x"00000725",
			445 => x"00000725",
			446 => x"00000725",
			447 => x"0505df04",
			448 => x"00000725",
			449 => x"011d0725",
			450 => x"06011804",
			451 => x"00000725",
			452 => x"0804f508",
			453 => x"01002304",
			454 => x"00000725",
			455 => x"fe8a0725",
			456 => x"00000725",
			457 => x"01002328",
			458 => x"0f05da20",
			459 => x"0601490c",
			460 => x"0f05d208",
			461 => x"0c05a404",
			462 => x"ffb70789",
			463 => x"00000789",
			464 => x"00000789",
			465 => x"06016310",
			466 => x"02087c04",
			467 => x"00000789",
			468 => x"041a6b08",
			469 => x"0506a704",
			470 => x"00a50789",
			471 => x"00000789",
			472 => x"00000789",
			473 => x"00000789",
			474 => x"0505df04",
			475 => x"00000789",
			476 => x"00d30789",
			477 => x"0416b608",
			478 => x"06011804",
			479 => x"00000789",
			480 => x"fe8e0789",
			481 => x"00000789",
			482 => x"040e6304",
			483 => x"fe6a07cd",
			484 => x"0d05f704",
			485 => x"fe6107cd",
			486 => x"06017118",
			487 => x"0007e50c",
			488 => x"02085204",
			489 => x"000007cd",
			490 => x"01007104",
			491 => x"01a107cd",
			492 => x"000007cd",
			493 => x"06014e04",
			494 => x"fe7e07cd",
			495 => x"0208ad04",
			496 => x"ff5407cd",
			497 => x"014e07cd",
			498 => x"fec407cd",
			499 => x"0415af14",
			500 => x"040e6304",
			501 => x"fe650831",
			502 => x"0a030d0c",
			503 => x"0c054504",
			504 => x"fea30831",
			505 => x"0e05e004",
			506 => x"028a0831",
			507 => x"ff260831",
			508 => x"feab0831",
			509 => x"0303e504",
			510 => x"fe870831",
			511 => x"06016c18",
			512 => x"09002310",
			513 => x"06014e08",
			514 => x"06014904",
			515 => x"fe1d0831",
			516 => x"00000831",
			517 => x"0a040504",
			518 => x"019a0831",
			519 => x"00000831",
			520 => x"08057c04",
			521 => x"01a20831",
			522 => x"00390831",
			523 => x"ffec0831",
			524 => x"0006970c",
			525 => x"09004f08",
			526 => x"07056104",
			527 => x"fe80089d",
			528 => x"01ca089d",
			529 => x"fe66089d",
			530 => x"0303f50c",
			531 => x"0007e508",
			532 => x"0303e504",
			533 => x"ffa2089d",
			534 => x"0100089d",
			535 => x"fe91089d",
			536 => x"0601921c",
			537 => x"09001f08",
			538 => x"0a03f204",
			539 => x"ff62089d",
			540 => x"002f089d",
			541 => x"02087c08",
			542 => x"01001604",
			543 => x"ffb5089d",
			544 => x"0059089d",
			545 => x"0007f604",
			546 => x"019e089d",
			547 => x"09002304",
			548 => x"0072089d",
			549 => x"0143089d",
			550 => x"fe17089d",
			551 => x"0415af20",
			552 => x"0413e914",
			553 => x"01003610",
			554 => x"0900550c",
			555 => x"09002d04",
			556 => x"fe5d0911",
			557 => x"09002e04",
			558 => x"ff670911",
			559 => x"fe970911",
			560 => x"00000911",
			561 => x"fe580911",
			562 => x"05066a04",
			563 => x"fe5a0911",
			564 => x"0100bc04",
			565 => x"02f60911",
			566 => x"fe710911",
			567 => x"0303e504",
			568 => x"fe5b0911",
			569 => x"00082614",
			570 => x"09001f04",
			571 => x"ffad0911",
			572 => x"0f058504",
			573 => x"01c00911",
			574 => x"07055d04",
			575 => x"03e50911",
			576 => x"0f059f04",
			577 => x"036b0911",
			578 => x"02fb0911",
			579 => x"fe7b0911",
			580 => x"0415af14",
			581 => x"09004f10",
			582 => x"0e03bd08",
			583 => x"0e036804",
			584 => x"fe82098d",
			585 => x"0000098d",
			586 => x"00049c04",
			587 => x"0000098d",
			588 => x"01c8098d",
			589 => x"fe66098d",
			590 => x"0303f50c",
			591 => x"0007e508",
			592 => x"0303e504",
			593 => x"ff29098d",
			594 => x"0117098d",
			595 => x"fe85098d",
			596 => x"0100231c",
			597 => x"09001f08",
			598 => x"0a03f204",
			599 => x"ff48098d",
			600 => x"0046098d",
			601 => x"02087c08",
			602 => x"01001604",
			603 => x"ff99098d",
			604 => x"0072098d",
			605 => x"041a5008",
			606 => x"041a0104",
			607 => x"01a0098d",
			608 => x"00fc098d",
			609 => x"0000098d",
			610 => x"ff8b098d",
			611 => x"040e6304",
			612 => x"fe7509fb",
			613 => x"0c059b1c",
			614 => x"03041d0c",
			615 => x"0705d208",
			616 => x"01001204",
			617 => x"000009fb",
			618 => x"fefd09fb",
			619 => x"000009fb",
			620 => x"0900390c",
			621 => x"0505df04",
			622 => x"000009fb",
			623 => x"0506a604",
			624 => x"009909fb",
			625 => x"000009fb",
			626 => x"000009fb",
			627 => x"01007314",
			628 => x"01001610",
			629 => x"06014904",
			630 => x"ffab09fb",
			631 => x"06016008",
			632 => x"0303e504",
			633 => x"000009fb",
			634 => x"009609fb",
			635 => x"000009fb",
			636 => x"014f09fb",
			637 => x"000009fb",
			638 => x"000009fd",
			639 => x"00000a01",
			640 => x"00000a05",
			641 => x"00000a09",
			642 => x"00000a0d",
			643 => x"00000a11",
			644 => x"00000a15",
			645 => x"00000a19",
			646 => x"00000a1d",
			647 => x"00000a21",
			648 => x"00000a25",
			649 => x"00000a29",
			650 => x"00000a2d",
			651 => x"00000a31",
			652 => x"00000a35",
			653 => x"00000a39",
			654 => x"00000a3d",
			655 => x"00000a41",
			656 => x"00000a45",
			657 => x"00000a49",
			658 => x"00000a4d",
			659 => x"00000a51",
			660 => x"00000a55",
			661 => x"00000a59",
			662 => x"00000a5d",
			663 => x"00000a61",
			664 => x"00000a65",
			665 => x"00000a69",
			666 => x"00000a6d",
			667 => x"00000a71",
			668 => x"00000a75",
			669 => x"00000a79",
			670 => x"00000a7d",
			671 => x"00000a81",
			672 => x"00000a85",
			673 => x"00000a89",
			674 => x"00000a8d",
			675 => x"00000a91",
			676 => x"0705a404",
			677 => x"ff410a9d",
			678 => x"00000a9d",
			679 => x"040e6304",
			680 => x"ffac0aa9",
			681 => x"00000aa9",
			682 => x"01004504",
			683 => x"00000ab5",
			684 => x"ffb50ab5",
			685 => x"09004f04",
			686 => x"00000ac1",
			687 => x"ffd60ac1",
			688 => x"01002304",
			689 => x"00000acd",
			690 => x"ffe20acd",
			691 => x"0705a404",
			692 => x"ffe70ad9",
			693 => x"00000ad9",
			694 => x"040e6304",
			695 => x"ff410aed",
			696 => x"0007e504",
			697 => x"00010aed",
			698 => x"00000aed",
			699 => x"040e6304",
			700 => x"ff880b01",
			701 => x"06017504",
			702 => x"00080b01",
			703 => x"00000b01",
			704 => x"0c059b08",
			705 => x"0d069204",
			706 => x"ffde0b15",
			707 => x"00000b15",
			708 => x"00000b15",
			709 => x"09004f08",
			710 => x"0007f604",
			711 => x"001d0b31",
			712 => x"00000b31",
			713 => x"04116204",
			714 => x"ffc80b31",
			715 => x"00000b31",
			716 => x"0100470c",
			717 => x"0007e508",
			718 => x"00049c04",
			719 => x"00000b4d",
			720 => x"00110b4d",
			721 => x"00000b4d",
			722 => x"ff4b0b4d",
			723 => x"0705a90c",
			724 => x"06012d04",
			725 => x"00000b69",
			726 => x"0418f304",
			727 => x"ff930b69",
			728 => x"00000b69",
			729 => x"00000b69",
			730 => x"0d06770c",
			731 => x"0c059b08",
			732 => x"0b05d604",
			733 => x"ffd90b85",
			734 => x"00000b85",
			735 => x"00000b85",
			736 => x"00000b85",
			737 => x"0705d20c",
			738 => x"0e032004",
			739 => x"00000ba1",
			740 => x"02096604",
			741 => x"ffe60ba1",
			742 => x"00000ba1",
			743 => x"00000ba1",
			744 => x"0705a90c",
			745 => x"06012d04",
			746 => x"00000bcd",
			747 => x"0418f304",
			748 => x"ff8b0bcd",
			749 => x"00000bcd",
			750 => x"02087e04",
			751 => x"00000bcd",
			752 => x"020a5004",
			753 => x"001a0bcd",
			754 => x"00000bcd",
			755 => x"01004510",
			756 => x"0f05c304",
			757 => x"00000bf1",
			758 => x"0c050b04",
			759 => x"00000bf1",
			760 => x"09002204",
			761 => x"00000bf1",
			762 => x"005b0bf1",
			763 => x"ff070bf1",
			764 => x"0208a404",
			765 => x"ffdc0c15",
			766 => x"0100470c",
			767 => x"01001204",
			768 => x"00000c15",
			769 => x"0e030004",
			770 => x"00000c15",
			771 => x"000e0c15",
			772 => x"00000c15",
			773 => x"0705d210",
			774 => x"0e032004",
			775 => x"00000c39",
			776 => x"0600ff04",
			777 => x"00000c39",
			778 => x"0c05bc04",
			779 => x"ffd60c39",
			780 => x"00000c39",
			781 => x"00000c39",
			782 => x"07056108",
			783 => x"0416b604",
			784 => x"feec0c65",
			785 => x"00000c65",
			786 => x"0601640c",
			787 => x"09002304",
			788 => x"00000c65",
			789 => x"0900a804",
			790 => x"00730c65",
			791 => x"00000c65",
			792 => x"00000c65",
			793 => x"09003914",
			794 => x"0f058504",
			795 => x"00000c99",
			796 => x"08056f0c",
			797 => x"0b061b08",
			798 => x"0505df04",
			799 => x"00000c99",
			800 => x"007f0c99",
			801 => x"00000c99",
			802 => x"00000c99",
			803 => x"0705d104",
			804 => x"fed30c99",
			805 => x"00000c99",
			806 => x"04116204",
			807 => x"febf0cc5",
			808 => x"06014904",
			809 => x"00000cc5",
			810 => x"0a040c0c",
			811 => x"0f070f08",
			812 => x"0f057204",
			813 => x"00000cc5",
			814 => x"00ca0cc5",
			815 => x"00000cc5",
			816 => x"00000cc5",
			817 => x"0416b60c",
			818 => x"01002308",
			819 => x"0c058104",
			820 => x"ffde0d09",
			821 => x"00000d09",
			822 => x"fe7b0d09",
			823 => x"02088b08",
			824 => x"09002504",
			825 => x"feed0d09",
			826 => x"00000d09",
			827 => x"0303e504",
			828 => x"00000d09",
			829 => x"041a6b08",
			830 => x"09001f04",
			831 => x"00000d09",
			832 => x"01690d09",
			833 => x"00000d09",
			834 => x"0705a308",
			835 => x"0418f304",
			836 => x"fe990d45",
			837 => x"00000d45",
			838 => x"01007314",
			839 => x"09002510",
			840 => x"0e032608",
			841 => x"0303e504",
			842 => x"00000d45",
			843 => x"00010d45",
			844 => x"03040e04",
			845 => x"00000d45",
			846 => x"ffc00d45",
			847 => x"00c90d45",
			848 => x"ffaa0d45",
			849 => x"0c052704",
			850 => x"fee00d81",
			851 => x"06016410",
			852 => x"0f058504",
			853 => x"00000d81",
			854 => x"041a0108",
			855 => x"01006104",
			856 => x"00be0d81",
			857 => x"00000d81",
			858 => x"00000d81",
			859 => x"05060804",
			860 => x"00000d81",
			861 => x"0418f304",
			862 => x"ffe40d81",
			863 => x"00000d81",
			864 => x"0415af0c",
			865 => x"01004508",
			866 => x"0505f904",
			867 => x"fe6b0dcd",
			868 => x"026c0dcd",
			869 => x"fe640dcd",
			870 => x"0303e504",
			871 => x"fe750dcd",
			872 => x"0900210c",
			873 => x"06014e04",
			874 => x"fe3c0dcd",
			875 => x"0a03fd04",
			876 => x"01bc0dcd",
			877 => x"00000dcd",
			878 => x"041a6b08",
			879 => x"00083104",
			880 => x"01a70dcd",
			881 => x"00000dcd",
			882 => x"00000dcd",
			883 => x"040e6304",
			884 => x"fe830e11",
			885 => x"0c059b10",
			886 => x"0004a004",
			887 => x"00000e11",
			888 => x"0418d408",
			889 => x"0705d204",
			890 => x"ff750e11",
			891 => x"00000e11",
			892 => x"00000e11",
			893 => x"03073b0c",
			894 => x"02089804",
			895 => x"00000e11",
			896 => x"041a5004",
			897 => x"01150e11",
			898 => x"00000e11",
			899 => x"00000e11",
			900 => x"0415af14",
			901 => x"01003608",
			902 => x"05066a04",
			903 => x"fe5e0e6d",
			904 => x"03fa0e6d",
			905 => x"01004708",
			906 => x"01004304",
			907 => x"fe610e6d",
			908 => x"fecf0e6d",
			909 => x"fe5b0e6d",
			910 => x"0f057204",
			911 => x"fe620e6d",
			912 => x"041a6b10",
			913 => x"0505f604",
			914 => x"00000e6d",
			915 => x"09001f04",
			916 => x"00310e6d",
			917 => x"00082604",
			918 => x"02660e6d",
			919 => x"ff210e6d",
			920 => x"06014b04",
			921 => x"fda60e6d",
			922 => x"00ee0e6d",
			923 => x"0416b610",
			924 => x"040f7004",
			925 => x"fe6c0ec9",
			926 => x"0705a404",
			927 => x"fe8b0ec9",
			928 => x"0900a804",
			929 => x"011a0ec9",
			930 => x"ff3a0ec9",
			931 => x"02088b08",
			932 => x"09002504",
			933 => x"fea30ec9",
			934 => x"00000ec9",
			935 => x"01001614",
			936 => x"06014908",
			937 => x"0a03dc04",
			938 => x"00000ec9",
			939 => x"fefd0ec9",
			940 => x"0705a304",
			941 => x"ff720ec9",
			942 => x"00082604",
			943 => x"011e0ec9",
			944 => x"00000ec9",
			945 => x"01790ec9",
			946 => x"09003924",
			947 => x"0f05d21c",
			948 => x"0601490c",
			949 => x"01001808",
			950 => x"09002a04",
			951 => x"fef70f35",
			952 => x"00000f35",
			953 => x"00000f35",
			954 => x"0a04020c",
			955 => x"02087c04",
			956 => x"00000f35",
			957 => x"0506a604",
			958 => x"00d90f35",
			959 => x"00000f35",
			960 => x"00000f35",
			961 => x"0505df04",
			962 => x"00000f35",
			963 => x"01330f35",
			964 => x"00053e08",
			965 => x"01003204",
			966 => x"00000f35",
			967 => x"fe780f35",
			968 => x"0c059c04",
			969 => x"ff2f0f35",
			970 => x"01007304",
			971 => x"007c0f35",
			972 => x"00000f35",
			973 => x"09003924",
			974 => x"0f05d21c",
			975 => x"06014908",
			976 => x"09002604",
			977 => x"ff290f99",
			978 => x"00000f99",
			979 => x"0601630c",
			980 => x"00082608",
			981 => x"02087c04",
			982 => x"00000f99",
			983 => x"00d30f99",
			984 => x"00000f99",
			985 => x"01001604",
			986 => x"fff80f99",
			987 => x"00000f99",
			988 => x"0505df04",
			989 => x"00000f99",
			990 => x"01280f99",
			991 => x"06011804",
			992 => x"00000f99",
			993 => x"0804f508",
			994 => x"01002304",
			995 => x"00000f99",
			996 => x"fe850f99",
			997 => x"00000f99",
			998 => x"04129904",
			999 => x"fe980fe5",
			1000 => x"0c059b10",
			1001 => x"03041d0c",
			1002 => x"01001504",
			1003 => x"00000fe5",
			1004 => x"0705d204",
			1005 => x"ff780fe5",
			1006 => x"00000fe5",
			1007 => x"00000fe5",
			1008 => x"02087e04",
			1009 => x"00000fe5",
			1010 => x"01001204",
			1011 => x"00000fe5",
			1012 => x"01007308",
			1013 => x"00081204",
			1014 => x"00d20fe5",
			1015 => x"00000fe5",
			1016 => x"00000fe5",
			1017 => x"0416b610",
			1018 => x"04116204",
			1019 => x"fe721041",
			1020 => x"0705a104",
			1021 => x"fec81041",
			1022 => x"01007904",
			1023 => x"00ae1041",
			1024 => x"00001041",
			1025 => x"0f058508",
			1026 => x"09002504",
			1027 => x"ff2e1041",
			1028 => x"00001041",
			1029 => x"041a6b14",
			1030 => x"0b059304",
			1031 => x"00001041",
			1032 => x"0b061b0c",
			1033 => x"0a040208",
			1034 => x"09002004",
			1035 => x"00001041",
			1036 => x"01571041",
			1037 => x"00001041",
			1038 => x"00001041",
			1039 => x"00001041",
			1040 => x"0415af24",
			1041 => x"0413e918",
			1042 => x"01003614",
			1043 => x"0900550c",
			1044 => x"09002d04",
			1045 => x"fe6110ad",
			1046 => x"09002e04",
			1047 => x"ff8010ad",
			1048 => x"fea210ad",
			1049 => x"00048504",
			1050 => x"fed410ad",
			1051 => x"010210ad",
			1052 => x"fe5a10ad",
			1053 => x"05066a04",
			1054 => x"fe5d10ad",
			1055 => x"0100bc04",
			1056 => x"029c10ad",
			1057 => x"fe7810ad",
			1058 => x"0f057204",
			1059 => x"fe5f10ad",
			1060 => x"0008260c",
			1061 => x"0303e504",
			1062 => x"fe7d10ad",
			1063 => x"01001204",
			1064 => x"017310ad",
			1065 => x"02a410ad",
			1066 => x"fe8c10ad",
			1067 => x"0415af14",
			1068 => x"040e6304",
			1069 => x"fe651111",
			1070 => x"0a030d0c",
			1071 => x"0c054504",
			1072 => x"fe921111",
			1073 => x"0e05e004",
			1074 => x"031f1111",
			1075 => x"fef91111",
			1076 => x"fea01111",
			1077 => x"0303e504",
			1078 => x"fe791111",
			1079 => x"09002310",
			1080 => x"06014a04",
			1081 => x"fdd61111",
			1082 => x"0208a408",
			1083 => x"0419b104",
			1084 => x"00001111",
			1085 => x"ffc81111",
			1086 => x"01b31111",
			1087 => x"020a5008",
			1088 => x"08057c04",
			1089 => x"01a81111",
			1090 => x"00531111",
			1091 => x"fffe1111",
			1092 => x"0415af10",
			1093 => x"0100360c",
			1094 => x"0505f904",
			1095 => x"fe66116d",
			1096 => x"0414a404",
			1097 => x"036c116d",
			1098 => x"019c116d",
			1099 => x"fe63116d",
			1100 => x"0303e504",
			1101 => x"fe66116d",
			1102 => x"09001f08",
			1103 => x"06014e04",
			1104 => x"fe68116d",
			1105 => x"0130116d",
			1106 => x"041a6b10",
			1107 => x"0a04100c",
			1108 => x"02085b04",
			1109 => x"ffbf116d",
			1110 => x"09003904",
			1111 => x"01d8116d",
			1112 => x"0105116d",
			1113 => x"fead116d",
			1114 => x"ff90116d",
			1115 => x"040e6304",
			1116 => x"fe6a11b9",
			1117 => x"07056108",
			1118 => x"0d05f704",
			1119 => x"fe7211b9",
			1120 => x"000011b9",
			1121 => x"06017018",
			1122 => x"0007e50c",
			1123 => x"02085204",
			1124 => x"000011b9",
			1125 => x"01009004",
			1126 => x"019c11b9",
			1127 => x"000011b9",
			1128 => x"06014e04",
			1129 => x"fe9611b9",
			1130 => x"0208ad04",
			1131 => x"ff6f11b9",
			1132 => x"014211b9",
			1133 => x"fed911b9",
			1134 => x"040e6304",
			1135 => x"fe8611fd",
			1136 => x"02085204",
			1137 => x"ffc611fd",
			1138 => x"06016314",
			1139 => x"041a0110",
			1140 => x"07054504",
			1141 => x"000011fd",
			1142 => x"01005808",
			1143 => x"0f058504",
			1144 => x"000011fd",
			1145 => x"012d11fd",
			1146 => x"000011fd",
			1147 => x"000011fd",
			1148 => x"04192604",
			1149 => x"ffe811fd",
			1150 => x"000011fd",
			1151 => x"0006a01c",
			1152 => x"00068610",
			1153 => x"0100320c",
			1154 => x"0505f904",
			1155 => x"fe511271",
			1156 => x"00060d04",
			1157 => x"09cf1271",
			1158 => x"063c1271",
			1159 => x"fe4f1271",
			1160 => x"03044604",
			1161 => x"fe591271",
			1162 => x"0100b404",
			1163 => x"06531271",
			1164 => x"fe721271",
			1165 => x"0303e504",
			1166 => x"fe541271",
			1167 => x"0a040914",
			1168 => x"0f057204",
			1169 => x"fe9c1271",
			1170 => x"0008260c",
			1171 => x"06017308",
			1172 => x"0d062b04",
			1173 => x"089f1271",
			1174 => x"06221271",
			1175 => x"00581271",
			1176 => x"fecc1271",
			1177 => x"0e031804",
			1178 => x"003d1271",
			1179 => x"fe671271",
			1180 => x"040e6304",
			1181 => x"fe6e12cd",
			1182 => x"02085208",
			1183 => x"0c05a204",
			1184 => x"febc12cd",
			1185 => x"000012cd",
			1186 => x"06016318",
			1187 => x"0007e50c",
			1188 => x"07053204",
			1189 => x"000012cd",
			1190 => x"0900a804",
			1191 => x"018b12cd",
			1192 => x"000012cd",
			1193 => x"06014e04",
			1194 => x"ff0d12cd",
			1195 => x"0208ad04",
			1196 => x"000012cd",
			1197 => x"010212cd",
			1198 => x"06017504",
			1199 => x"000012cd",
			1200 => x"07055d04",
			1201 => x"000012cd",
			1202 => x"ff0412cd",
			1203 => x"0415af24",
			1204 => x"01003620",
			1205 => x"09002d08",
			1206 => x"0a030404",
			1207 => x"00001359",
			1208 => x"feed1359",
			1209 => x"08041e0c",
			1210 => x"0a02c608",
			1211 => x"0a02ac04",
			1212 => x"ffd51359",
			1213 => x"00111359",
			1214 => x"ffc21359",
			1215 => x"08048f08",
			1216 => x"0a032104",
			1217 => x"00001359",
			1218 => x"00571359",
			1219 => x"00001359",
			1220 => x"fe691359",
			1221 => x"0208930c",
			1222 => x"09002504",
			1223 => x"feb11359",
			1224 => x"0a036304",
			1225 => x"00001359",
			1226 => x"00991359",
			1227 => x"041a320c",
			1228 => x"06016608",
			1229 => x"09001f04",
			1230 => x"00001359",
			1231 => x"01901359",
			1232 => x"00001359",
			1233 => x"06014a04",
			1234 => x"ff701359",
			1235 => x"0208d604",
			1236 => x"00001359",
			1237 => x"009d1359",
			1238 => x"04129904",
			1239 => x"fe9d13b5",
			1240 => x"0c059b14",
			1241 => x"0e034a10",
			1242 => x"0e032004",
			1243 => x"000013b5",
			1244 => x"0d069208",
			1245 => x"0705e504",
			1246 => x"ff8913b5",
			1247 => x"000013b5",
			1248 => x"000013b5",
			1249 => x"000013b5",
			1250 => x"06014904",
			1251 => x"000013b5",
			1252 => x"06016310",
			1253 => x"09001f04",
			1254 => x"000013b5",
			1255 => x"0f057204",
			1256 => x"000013b5",
			1257 => x"0f06ea04",
			1258 => x"00be13b5",
			1259 => x"000013b5",
			1260 => x"000013b5",
			1261 => x"040e6304",
			1262 => x"fe701413",
			1263 => x"02085208",
			1264 => x"0c05a204",
			1265 => x"fedf1413",
			1266 => x"00001413",
			1267 => x"01004720",
			1268 => x"01001614",
			1269 => x"0007e508",
			1270 => x"0e031804",
			1271 => x"00001413",
			1272 => x"00a81413",
			1273 => x"0e034308",
			1274 => x"0d066d04",
			1275 => x"00001413",
			1276 => x"005e1413",
			1277 => x"ff4c1413",
			1278 => x"0505df04",
			1279 => x"00001413",
			1280 => x"00085504",
			1281 => x"017e1413",
			1282 => x"00001413",
			1283 => x"ff3e1413",
			1284 => x"00001415",
			1285 => x"00001419",
			1286 => x"0000141d",
			1287 => x"00001421",
			1288 => x"00001425",
			1289 => x"00001429",
			1290 => x"0000142d",
			1291 => x"00001431",
			1292 => x"00001435",
			1293 => x"00001439",
			1294 => x"0000143d",
			1295 => x"00001441",
			1296 => x"00001445",
			1297 => x"00001449",
			1298 => x"0000144d",
			1299 => x"00001451",
			1300 => x"00001455",
			1301 => x"00001459",
			1302 => x"0000145d",
			1303 => x"00001461",
			1304 => x"00001465",
			1305 => x"00001469",
			1306 => x"0000146d",
			1307 => x"00001471",
			1308 => x"00001475",
			1309 => x"00001479",
			1310 => x"0000147d",
			1311 => x"00001481",
			1312 => x"00001485",
			1313 => x"00001489",
			1314 => x"0000148d",
			1315 => x"00001491",
			1316 => x"00001495",
			1317 => x"00001499",
			1318 => x"0000149d",
			1319 => x"000014a1",
			1320 => x"000014a5",
			1321 => x"000014a9",
			1322 => x"040e6304",
			1323 => x"ff5414b5",
			1324 => x"000014b5",
			1325 => x"07054504",
			1326 => x"ffb214c1",
			1327 => x"000014c1",
			1328 => x"0705a404",
			1329 => x"ffa614cd",
			1330 => x"000014cd",
			1331 => x"09004f04",
			1332 => x"000014d9",
			1333 => x"ffd914d9",
			1334 => x"09003904",
			1335 => x"000014e5",
			1336 => x"ffe514e5",
			1337 => x"0705a404",
			1338 => x"ffe914f1",
			1339 => x"000014f1",
			1340 => x"01003608",
			1341 => x"02087e04",
			1342 => x"00001505",
			1343 => x"00081505",
			1344 => x"ff501505",
			1345 => x"09004f04",
			1346 => x"00001519",
			1347 => x"04116204",
			1348 => x"ffaa1519",
			1349 => x"00001519",
			1350 => x"0b056508",
			1351 => x"0e032004",
			1352 => x"00001535",
			1353 => x"ff781535",
			1354 => x"06016004",
			1355 => x"00081535",
			1356 => x"00001535",
			1357 => x"09004f08",
			1358 => x"0007f604",
			1359 => x"00161551",
			1360 => x"00001551",
			1361 => x"04116204",
			1362 => x"ffcd1551",
			1363 => x"00001551",
			1364 => x"0100360c",
			1365 => x"06014904",
			1366 => x"0000156d",
			1367 => x"02087e04",
			1368 => x"0000156d",
			1369 => x"0034156d",
			1370 => x"ff62156d",
			1371 => x"0705a404",
			1372 => x"ff961589",
			1373 => x"02087e04",
			1374 => x"00001589",
			1375 => x"020a2004",
			1376 => x"002d1589",
			1377 => x"00001589",
			1378 => x"0d06770c",
			1379 => x"0c059b08",
			1380 => x"0b05d604",
			1381 => x"ffdc15a5",
			1382 => x"000015a5",
			1383 => x"000015a5",
			1384 => x"000015a5",
			1385 => x"0c059b0c",
			1386 => x"0d069208",
			1387 => x"0705d204",
			1388 => x"ffde15c1",
			1389 => x"000015c1",
			1390 => x"000015c1",
			1391 => x"000015c1",
			1392 => x"07054504",
			1393 => x"fecd15e5",
			1394 => x"01005a0c",
			1395 => x"0f058504",
			1396 => x"000015e5",
			1397 => x"0007e504",
			1398 => x"00a815e5",
			1399 => x"000015e5",
			1400 => x"000015e5",
			1401 => x"0208a404",
			1402 => x"ffd61609",
			1403 => x"0100470c",
			1404 => x"09001f04",
			1405 => x"00001609",
			1406 => x"0e030004",
			1407 => x"00001609",
			1408 => x"001c1609",
			1409 => x"00001609",
			1410 => x"0705a904",
			1411 => x"ffc7162d",
			1412 => x"0100790c",
			1413 => x"09001f04",
			1414 => x"0000162d",
			1415 => x"0d065104",
			1416 => x"0000162d",
			1417 => x"001a162d",
			1418 => x"0000162d",
			1419 => x"0c059b10",
			1420 => x"0e031004",
			1421 => x"00001651",
			1422 => x"0d069208",
			1423 => x"0705d204",
			1424 => x"ffc61651",
			1425 => x"00001651",
			1426 => x"00001651",
			1427 => x"00001651",
			1428 => x"07056108",
			1429 => x"04192604",
			1430 => x"ff15167d",
			1431 => x"0000167d",
			1432 => x"0601630c",
			1433 => x"06014904",
			1434 => x"0000167d",
			1435 => x"06016004",
			1436 => x"0038167d",
			1437 => x"0000167d",
			1438 => x"0000167d",
			1439 => x"07056108",
			1440 => x"04192604",
			1441 => x"ff0a16b1",
			1442 => x"000016b1",
			1443 => x"06016310",
			1444 => x"09002304",
			1445 => x"000016b1",
			1446 => x"01007308",
			1447 => x"0e030804",
			1448 => x"000016b1",
			1449 => x"006316b1",
			1450 => x"000016b1",
			1451 => x"000016b1",
			1452 => x"0705a904",
			1453 => x"ffc116dd",
			1454 => x"01007910",
			1455 => x"02087e04",
			1456 => x"000016dd",
			1457 => x"041a3208",
			1458 => x"09001f04",
			1459 => x"000016dd",
			1460 => x"005516dd",
			1461 => x"000016dd",
			1462 => x"000016dd",
			1463 => x"0100361c",
			1464 => x"0d06470c",
			1465 => x"03041d08",
			1466 => x"0b05b804",
			1467 => x"ff541721",
			1468 => x"00001721",
			1469 => x"00001721",
			1470 => x"02087e08",
			1471 => x"09002704",
			1472 => x"ffff1721",
			1473 => x"00001721",
			1474 => x"00080104",
			1475 => x"00fe1721",
			1476 => x"00001721",
			1477 => x"00069704",
			1478 => x"fe8c1721",
			1479 => x"00001721",
			1480 => x"040e6304",
			1481 => x"fea8175d",
			1482 => x"0c059b0c",
			1483 => x"03041d08",
			1484 => x"0705e504",
			1485 => x"ff99175d",
			1486 => x"0000175d",
			1487 => x"0000175d",
			1488 => x"0100730c",
			1489 => x"02089804",
			1490 => x"0000175d",
			1491 => x"041a5004",
			1492 => x"00c1175d",
			1493 => x"0000175d",
			1494 => x"0000175d",
			1495 => x"07056108",
			1496 => x"0c054c04",
			1497 => x"fea71799",
			1498 => x"00001799",
			1499 => x"01007114",
			1500 => x"0007ba04",
			1501 => x"00cf1799",
			1502 => x"06014d04",
			1503 => x"ffd51799",
			1504 => x"06016808",
			1505 => x"0c056204",
			1506 => x"00001799",
			1507 => x"003e1799",
			1508 => x"00001799",
			1509 => x"ffba1799",
			1510 => x"040e6304",
			1511 => x"fe7e17cd",
			1512 => x"06017514",
			1513 => x"02084b04",
			1514 => x"ff8917cd",
			1515 => x"0007f60c",
			1516 => x"07054704",
			1517 => x"000017cd",
			1518 => x"01005804",
			1519 => x"013f17cd",
			1520 => x"000017cd",
			1521 => x"000017cd",
			1522 => x"ff3317cd",
			1523 => x"0416b610",
			1524 => x"040f7004",
			1525 => x"fe6d1829",
			1526 => x"0705a404",
			1527 => x"fe9c1829",
			1528 => x"0900a804",
			1529 => x"01051829",
			1530 => x"ff521829",
			1531 => x"0f05d218",
			1532 => x"06014908",
			1533 => x"09002604",
			1534 => x"fe8c1829",
			1535 => x"00001829",
			1536 => x"06016308",
			1537 => x"0f058504",
			1538 => x"00001829",
			1539 => x"012e1829",
			1540 => x"0705d004",
			1541 => x"ff591829",
			1542 => x"00001829",
			1543 => x"09002204",
			1544 => x"00001829",
			1545 => x"016f1829",
			1546 => x"0415af18",
			1547 => x"040e6304",
			1548 => x"fe671885",
			1549 => x"0a030d0c",
			1550 => x"0c054504",
			1551 => x"fed31885",
			1552 => x"0f082204",
			1553 => x"02261885",
			1554 => x"ff9f1885",
			1555 => x"04151804",
			1556 => x"fe981885",
			1557 => x"fff91885",
			1558 => x"0f057204",
			1559 => x"febe1885",
			1560 => x"0007f608",
			1561 => x"0b056504",
			1562 => x"00001885",
			1563 => x"01981885",
			1564 => x"06014e04",
			1565 => x"fe661885",
			1566 => x"0a040c04",
			1567 => x"017b1885",
			1568 => x"ff4a1885",
			1569 => x"0415f31c",
			1570 => x"0415af14",
			1571 => x"0413e908",
			1572 => x"01004704",
			1573 => x"d39118f9",
			1574 => x"d37718f9",
			1575 => x"05066a04",
			1576 => x"d37818f9",
			1577 => x"0100b404",
			1578 => x"eb6f18f9",
			1579 => x"d38518f9",
			1580 => x"02089804",
			1581 => x"d38b18f9",
			1582 => x"ead018f9",
			1583 => x"0f05850c",
			1584 => x"0007cf08",
			1585 => x"02084d04",
			1586 => x"d3a918f9",
			1587 => x"e5e218f9",
			1588 => x"d37918f9",
			1589 => x"00082610",
			1590 => x"0f059f08",
			1591 => x"0007f604",
			1592 => x"ea3518f9",
			1593 => x"d5ac18f9",
			1594 => x"05062604",
			1595 => x"e29618f9",
			1596 => x"ec4e18f9",
			1597 => x"d3ae18f9",
			1598 => x"00069710",
			1599 => x"040e6304",
			1600 => x"fe68195d",
			1601 => x"07056104",
			1602 => x"fe91195d",
			1603 => x"01007304",
			1604 => x"01c3195d",
			1605 => x"fea5195d",
			1606 => x"09002310",
			1607 => x"06014a04",
			1608 => x"fe8e195d",
			1609 => x"00082608",
			1610 => x"0303e504",
			1611 => x"0000195d",
			1612 => x"015d195d",
			1613 => x"ff47195d",
			1614 => x"0a040c10",
			1615 => x"0415af04",
			1616 => x"0000195d",
			1617 => x"00081208",
			1618 => x"0303e504",
			1619 => x"0000195d",
			1620 => x"0197195d",
			1621 => x"0000195d",
			1622 => x"ff66195d",
			1623 => x"0415af10",
			1624 => x"0100470c",
			1625 => x"0705a404",
			1626 => x"fe6019b9",
			1627 => x"00061504",
			1628 => x"066619b9",
			1629 => x"01dd19b9",
			1630 => x"fe5e19b9",
			1631 => x"0303e504",
			1632 => x"fe6519b9",
			1633 => x"041a6b14",
			1634 => x"0f058508",
			1635 => x"04194504",
			1636 => x"017719b9",
			1637 => x"fe9519b9",
			1638 => x"01001204",
			1639 => x"015919b9",
			1640 => x"020a5004",
			1641 => x"021719b9",
			1642 => x"016719b9",
			1643 => x"06014a04",
			1644 => x"fdd519b9",
			1645 => x"007919b9",
			1646 => x"0415af18",
			1647 => x"01003614",
			1648 => x"01002a08",
			1649 => x"0a035704",
			1650 => x"ff451a2d",
			1651 => x"00001a2d",
			1652 => x"08037a04",
			1653 => x"00001a2d",
			1654 => x"0a02c604",
			1655 => x"00451a2d",
			1656 => x"00001a2d",
			1657 => x"fe681a2d",
			1658 => x"02089310",
			1659 => x"0007c20c",
			1660 => x"0a037208",
			1661 => x"0a036304",
			1662 => x"ff991a2d",
			1663 => x"00001a2d",
			1664 => x"00911a2d",
			1665 => x"fe921a2d",
			1666 => x"041a3208",
			1667 => x"06016604",
			1668 => x"018f1a2d",
			1669 => x"00001a2d",
			1670 => x"06014a04",
			1671 => x"ff601a2d",
			1672 => x"0208d604",
			1673 => x"00001a2d",
			1674 => x"00b71a2d",
			1675 => x"09003920",
			1676 => x"0f058508",
			1677 => x"01001c04",
			1678 => x"ff2c1a89",
			1679 => x"00001a89",
			1680 => x"0303e504",
			1681 => x"00001a89",
			1682 => x"09001f04",
			1683 => x"00001a89",
			1684 => x"0b061b0c",
			1685 => x"00081208",
			1686 => x"0a040104",
			1687 => x"014b1a89",
			1688 => x"00001a89",
			1689 => x"00001a89",
			1690 => x"00001a89",
			1691 => x"0006f10c",
			1692 => x"06011804",
			1693 => x"00001a89",
			1694 => x"01002304",
			1695 => x"00001a89",
			1696 => x"fe7c1a89",
			1697 => x"00001a89",
			1698 => x"0415af14",
			1699 => x"01003608",
			1700 => x"05066a04",
			1701 => x"fe601aed",
			1702 => x"03ac1aed",
			1703 => x"01004708",
			1704 => x"01004304",
			1705 => x"fe641aed",
			1706 => x"fede1aed",
			1707 => x"fe5c1aed",
			1708 => x"0303e504",
			1709 => x"fe621aed",
			1710 => x"041a6b14",
			1711 => x"0f057204",
			1712 => x"feb61aed",
			1713 => x"09001f04",
			1714 => x"00741aed",
			1715 => x"0f058504",
			1716 => x"01561aed",
			1717 => x"0f059f04",
			1718 => x"02951aed",
			1719 => x"02351aed",
			1720 => x"06014a04",
			1721 => x"fdad1aed",
			1722 => x"008c1aed",
			1723 => x"00069714",
			1724 => x"09005d08",
			1725 => x"0505f904",
			1726 => x"fe721b51",
			1727 => x"02041b51",
			1728 => x"00053e04",
			1729 => x"fe651b51",
			1730 => x"0f070f04",
			1731 => x"02551b51",
			1732 => x"fe781b51",
			1733 => x"0303e504",
			1734 => x"fe861b51",
			1735 => x"06019218",
			1736 => x"09002310",
			1737 => x"06014e08",
			1738 => x"06014904",
			1739 => x"fdfa1b51",
			1740 => x"00001b51",
			1741 => x"0a040504",
			1742 => x"01a61b51",
			1743 => x"00001b51",
			1744 => x"08057c04",
			1745 => x"01a51b51",
			1746 => x"00441b51",
			1747 => x"fdc51b51",
			1748 => x"0415af10",
			1749 => x"0100450c",
			1750 => x"0505f904",
			1751 => x"fe691bad",
			1752 => x"0e03e704",
			1753 => x"01751bad",
			1754 => x"03341bad",
			1755 => x"fe631bad",
			1756 => x"0303e504",
			1757 => x"fe6d1bad",
			1758 => x"09001f08",
			1759 => x"06014e04",
			1760 => x"fe971bad",
			1761 => x"00f91bad",
			1762 => x"041a6b10",
			1763 => x"0f057204",
			1764 => x"ff3a1bad",
			1765 => x"041a3204",
			1766 => x"01b31bad",
			1767 => x"0f05da04",
			1768 => x"ffd71bad",
			1769 => x"01921bad",
			1770 => x"ffff1bad",
			1771 => x"0415af20",
			1772 => x"09004f1c",
			1773 => x"09003608",
			1774 => x"09003004",
			1775 => x"febb1c29",
			1776 => x"00001c29",
			1777 => x"01002108",
			1778 => x"0004bc04",
			1779 => x"01991c29",
			1780 => x"00001c29",
			1781 => x"0411a308",
			1782 => x"01002d04",
			1783 => x"ff3d1c29",
			1784 => x"00001c29",
			1785 => x"00951c29",
			1786 => x"fe661c29",
			1787 => x"0303f50c",
			1788 => x"0007e508",
			1789 => x"0303e504",
			1790 => x"ff551c29",
			1791 => x"00e81c29",
			1792 => x"fe9d1c29",
			1793 => x"020a4610",
			1794 => x"041a0108",
			1795 => x"02087c04",
			1796 => x"00001c29",
			1797 => x"01991c29",
			1798 => x"06014a04",
			1799 => x"fe6e1c29",
			1800 => x"01621c29",
			1801 => x"ff971c29",
			1802 => x"00069710",
			1803 => x"0100360c",
			1804 => x"0505f904",
			1805 => x"fe631c8d",
			1806 => x"00062204",
			1807 => x"04801c8d",
			1808 => x"01db1c8d",
			1809 => x"fe601c8d",
			1810 => x"0303e504",
			1811 => x"fe621c8d",
			1812 => x"06017818",
			1813 => x"09001f08",
			1814 => x"06014e04",
			1815 => x"fe511c8d",
			1816 => x"017c1c8d",
			1817 => x"0008260c",
			1818 => x"02085b04",
			1819 => x"ffa41c8d",
			1820 => x"00081204",
			1821 => x"01fd1c8d",
			1822 => x"016a1c8d",
			1823 => x"fed51c8d",
			1824 => x"08052704",
			1825 => x"fe551c8d",
			1826 => x"00001c8d",
			1827 => x"0415af10",
			1828 => x"0100470c",
			1829 => x"05066a04",
			1830 => x"fe651cf1",
			1831 => x"04141b04",
			1832 => x"03e01cf1",
			1833 => x"019c1cf1",
			1834 => x"fe621cf1",
			1835 => x"0303e504",
			1836 => x"fe691cf1",
			1837 => x"09001f08",
			1838 => x"0c05b904",
			1839 => x"fe5f1cf1",
			1840 => x"00001cf1",
			1841 => x"0a040c14",
			1842 => x"041a010c",
			1843 => x"02086c04",
			1844 => x"00af1cf1",
			1845 => x"020a4604",
			1846 => x"01cf1cf1",
			1847 => x"00b11cf1",
			1848 => x"06014d04",
			1849 => x"fe011cf1",
			1850 => x"01d41cf1",
			1851 => x"fea91cf1",
			1852 => x"040e6304",
			1853 => x"fe6f1d4d",
			1854 => x"02084b08",
			1855 => x"03043504",
			1856 => x"fece1d4d",
			1857 => x"00001d4d",
			1858 => x"06016318",
			1859 => x"0007e50c",
			1860 => x"07053204",
			1861 => x"00001d4d",
			1862 => x"01007304",
			1863 => x"01851d4d",
			1864 => x"00001d4d",
			1865 => x"06014e04",
			1866 => x"ff251d4d",
			1867 => x"0208ad04",
			1868 => x"00001d4d",
			1869 => x"00f11d4d",
			1870 => x"06017504",
			1871 => x"00001d4d",
			1872 => x"07055d04",
			1873 => x"00001d4d",
			1874 => x"ff1b1d4d",
			1875 => x"0415af10",
			1876 => x"0100470c",
			1877 => x"05066a04",
			1878 => x"fe671db1",
			1879 => x"0b061904",
			1880 => x"01ab1db1",
			1881 => x"034e1db1",
			1882 => x"fe631db1",
			1883 => x"0303e504",
			1884 => x"fe6f1db1",
			1885 => x"09001f08",
			1886 => x"0c05b904",
			1887 => x"fe8b1db1",
			1888 => x"00001db1",
			1889 => x"0a040c14",
			1890 => x"0f057204",
			1891 => x"ff451db1",
			1892 => x"041a0108",
			1893 => x"020a4604",
			1894 => x"01ba1db1",
			1895 => x"00701db1",
			1896 => x"06014d04",
			1897 => x"fe5d1db1",
			1898 => x"01be1db1",
			1899 => x"feda1db1",
			1900 => x"0415af28",
			1901 => x"0413e91c",
			1902 => x"01004718",
			1903 => x"09007b14",
			1904 => x"040e6304",
			1905 => x"fe541e35",
			1906 => x"09004608",
			1907 => x"040eab04",
			1908 => x"00311e35",
			1909 => x"fe641e35",
			1910 => x"040f7004",
			1911 => x"fe8d1e35",
			1912 => x"039e1e35",
			1913 => x"010d1e35",
			1914 => x"fe521e35",
			1915 => x"05066a04",
			1916 => x"fe541e35",
			1917 => x"0100b404",
			1918 => x"045e1e35",
			1919 => x"fe641e35",
			1920 => x"0f057204",
			1921 => x"fe581e35",
			1922 => x"09001f08",
			1923 => x"06014a04",
			1924 => x"fe3f1e35",
			1925 => x"00001e35",
			1926 => x"0008260c",
			1927 => x"00081208",
			1928 => x"0b056904",
			1929 => x"02ee1e35",
			1930 => x"04671e35",
			1931 => x"02e41e35",
			1932 => x"fe9d1e35",
			1933 => x"0415af24",
			1934 => x"04116204",
			1935 => x"fe641ebb",
			1936 => x"0a030d08",
			1937 => x"07057504",
			1938 => x"fe991ebb",
			1939 => x"03771ebb",
			1940 => x"0414ff10",
			1941 => x"0804240c",
			1942 => x"0a032304",
			1943 => x"febb1ebb",
			1944 => x"0a032704",
			1945 => x"01411ebb",
			1946 => x"00001ebb",
			1947 => x"fe7f1ebb",
			1948 => x"03045e04",
			1949 => x"fe7e1ebb",
			1950 => x"016c1ebb",
			1951 => x"0303e504",
			1952 => x"fe6b1ebb",
			1953 => x"0a040c18",
			1954 => x"0f057204",
			1955 => x"ff0e1ebb",
			1956 => x"041a010c",
			1957 => x"020a4608",
			1958 => x"02088b04",
			1959 => x"01401ebb",
			1960 => x"01c41ebb",
			1961 => x"008e1ebb",
			1962 => x"06014a04",
			1963 => x"fd471ebb",
			1964 => x"01c31ebb",
			1965 => x"fead1ebb",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(638, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(1284, initial_addr_3'length));
	end generate gen_rom_1;

	gen_rom_2: if SELECT_ROM = 2 generate
		bank <= (
			0 => x"00000005",
			1 => x"00000009",
			2 => x"0000000d",
			3 => x"0c060f04",
			4 => x"00000021",
			5 => x"0c064d04",
			6 => x"00070021",
			7 => x"00000021",
			8 => x"0b071008",
			9 => x"0b06bc04",
			10 => x"00000035",
			11 => x"fff30035",
			12 => x"00000035",
			13 => x"0b06dd04",
			14 => x"00000049",
			15 => x"0b076304",
			16 => x"000a0049",
			17 => x"00000049",
			18 => x"00032408",
			19 => x"0c05d704",
			20 => x"00000065",
			21 => x"001d0065",
			22 => x"0c063404",
			23 => x"ffd40065",
			24 => x"00000065",
			25 => x"0507e708",
			26 => x"0506f104",
			27 => x"00000081",
			28 => x"00120081",
			29 => x"05081f04",
			30 => x"fff40081",
			31 => x"00000081",
			32 => x"0b06dd04",
			33 => x"0000009d",
			34 => x"02092808",
			35 => x"0208ce04",
			36 => x"0000009d",
			37 => x"002b009d",
			38 => x"0000009d",
			39 => x"0209200c",
			40 => x"00030c08",
			41 => x"0207c504",
			42 => x"000000c1",
			43 => x"002800c1",
			44 => x"000000c1",
			45 => x"02097b04",
			46 => x"fff100c1",
			47 => x"000000c1",
			48 => x"0003240c",
			49 => x"0207c504",
			50 => x"000000e5",
			51 => x"02097804",
			52 => x"000c00e5",
			53 => x"000000e5",
			54 => x"020a5004",
			55 => x"fff800e5",
			56 => x"000000e5",
			57 => x"00030c0c",
			58 => x"02092808",
			59 => x"0207c504",
			60 => x"00000111",
			61 => x"001b0111",
			62 => x"00000111",
			63 => x"02099d04",
			64 => x"ffde0111",
			65 => x"020a2d04",
			66 => x"00050111",
			67 => x"00000111",
			68 => x"00037810",
			69 => x"09017d04",
			70 => x"00000135",
			71 => x"040ac908",
			72 => x"04094504",
			73 => x"00000135",
			74 => x"00100135",
			75 => x"00000135",
			76 => x"00000135",
			77 => x"040a2810",
			78 => x"07064604",
			79 => x"00000161",
			80 => x"04094504",
			81 => x"00000161",
			82 => x"0c05f204",
			83 => x"00000161",
			84 => x"003e0161",
			85 => x"0c063404",
			86 => x"ffd70161",
			87 => x"00000161",
			88 => x"06013e08",
			89 => x"0c05f204",
			90 => x"0000018d",
			91 => x"004e018d",
			92 => x"0c06320c",
			93 => x"04097204",
			94 => x"0000018d",
			95 => x"06016f04",
			96 => x"ffd1018d",
			97 => x"0000018d",
			98 => x"0000018d",
			99 => x"00030c08",
			100 => x"0b063c04",
			101 => x"000001c1",
			102 => x"000901c1",
			103 => x"0b06d208",
			104 => x"0b06bc04",
			105 => x"000001c1",
			106 => x"ffc601c1",
			107 => x"0b071e08",
			108 => x"0b06dd04",
			109 => x"000001c1",
			110 => x"001f01c1",
			111 => x"000001c1",
			112 => x"00030c08",
			113 => x"0b063c04",
			114 => x"000001fd",
			115 => x"000901fd",
			116 => x"0b06d208",
			117 => x"0b06bc04",
			118 => x"000001fd",
			119 => x"ffbd01fd",
			120 => x"0b071e08",
			121 => x"0b06dd04",
			122 => x"000001fd",
			123 => x"002201fd",
			124 => x"0b073304",
			125 => x"fffd01fd",
			126 => x"000001fd",
			127 => x"0b06dd08",
			128 => x"0901dd04",
			129 => x"ffe80231",
			130 => x"00000231",
			131 => x"07064604",
			132 => x"00000231",
			133 => x"07066c0c",
			134 => x"09017a04",
			135 => x"00000231",
			136 => x"09021f04",
			137 => x"005c0231",
			138 => x"00000231",
			139 => x"00000231",
			140 => x"0e098714",
			141 => x"0b072010",
			142 => x"0408db04",
			143 => x"0000025d",
			144 => x"06016208",
			145 => x"07068804",
			146 => x"ffd9025d",
			147 => x"0000025d",
			148 => x"0000025d",
			149 => x"0000025d",
			150 => x"0000025d",
			151 => x"040a3a14",
			152 => x"08025a04",
			153 => x"00000299",
			154 => x"0c05f604",
			155 => x"00000299",
			156 => x"0c065008",
			157 => x"00035304",
			158 => x"004d0299",
			159 => x"00000299",
			160 => x"00000299",
			161 => x"01014908",
			162 => x"0c06e504",
			163 => x"ffdc0299",
			164 => x"00000299",
			165 => x"00000299",
			166 => x"0e093310",
			167 => x"04091d04",
			168 => x"000002dd",
			169 => x"0a01ec04",
			170 => x"ffc102dd",
			171 => x"0a01f704",
			172 => x"000402dd",
			173 => x"ffef02dd",
			174 => x"040a3a10",
			175 => x"0101360c",
			176 => x"0309ef08",
			177 => x"03097804",
			178 => x"000002dd",
			179 => x"009402dd",
			180 => x"000002dd",
			181 => x"000002dd",
			182 => x"000002dd",
			183 => x"040a281c",
			184 => x"0e094014",
			185 => x"00030c0c",
			186 => x"0002ee04",
			187 => x"00000331",
			188 => x"0100e504",
			189 => x"00000331",
			190 => x"00410331",
			191 => x"0b06d204",
			192 => x"ffad0331",
			193 => x"00000331",
			194 => x"03097804",
			195 => x"00000331",
			196 => x"00c60331",
			197 => x"0901fc0c",
			198 => x"07072608",
			199 => x"08029904",
			200 => x"00000331",
			201 => x"ffaa0331",
			202 => x"00000331",
			203 => x"00000331",
			204 => x"040a3a18",
			205 => x"09018304",
			206 => x"0000036d",
			207 => x"01013610",
			208 => x"07063d04",
			209 => x"0000036d",
			210 => x"00035308",
			211 => x"0b06a504",
			212 => x"0000036d",
			213 => x"008a036d",
			214 => x"0000036d",
			215 => x"0000036d",
			216 => x"06018804",
			217 => x"fff4036d",
			218 => x"0000036d",
			219 => x"0e093308",
			220 => x"0d075504",
			221 => x"000003a9",
			222 => x"fffa03a9",
			223 => x"0d089a14",
			224 => x"09018304",
			225 => x"000003a9",
			226 => x"0e0a860c",
			227 => x"0d080e04",
			228 => x"000003a9",
			229 => x"09021b04",
			230 => x"003003a9",
			231 => x"000003a9",
			232 => x"000003a9",
			233 => x"000003a9",
			234 => x"0100f108",
			235 => x"0801cb04",
			236 => x"000003e5",
			237 => x"ffe103e5",
			238 => x"0f0ab614",
			239 => x"0e092404",
			240 => x"000003e5",
			241 => x"09018704",
			242 => x"000003e5",
			243 => x"01014e08",
			244 => x"0802fb04",
			245 => x"003b03e5",
			246 => x"000003e5",
			247 => x"000003e5",
			248 => x"000003e5",
			249 => x"040a2818",
			250 => x"0100e704",
			251 => x"00000429",
			252 => x"0309ef10",
			253 => x"0003530c",
			254 => x"0f090d04",
			255 => x"00000429",
			256 => x"03090f04",
			257 => x"00000429",
			258 => x"00320429",
			259 => x"00000429",
			260 => x"00000429",
			261 => x"01012e08",
			262 => x"030a6904",
			263 => x"fff70429",
			264 => x"00000429",
			265 => x"00000429",
			266 => x"0c05d804",
			267 => x"0000045d",
			268 => x"05082114",
			269 => x"00037810",
			270 => x"0d087f0c",
			271 => x"0d080b04",
			272 => x"0000045d",
			273 => x"07068604",
			274 => x"004b045d",
			275 => x"0000045d",
			276 => x"0000045d",
			277 => x"0000045d",
			278 => x"0000045d",
			279 => x"0c063018",
			280 => x"04091d04",
			281 => x"00000491",
			282 => x"0901dd10",
			283 => x"0c05da04",
			284 => x"00000491",
			285 => x"07062c04",
			286 => x"00000491",
			287 => x"01012a04",
			288 => x"ffa60491",
			289 => x"00000491",
			290 => x"00000491",
			291 => x"00000491",
			292 => x"040a0110",
			293 => x"0a01ec04",
			294 => x"000004e5",
			295 => x"0d081704",
			296 => x"000004e5",
			297 => x"0309d804",
			298 => x"004504e5",
			299 => x"000004e5",
			300 => x"0901d908",
			301 => x"0c063a04",
			302 => x"ff8504e5",
			303 => x"000004e5",
			304 => x"0c064d10",
			305 => x"0e098704",
			306 => x"000004e5",
			307 => x"01015508",
			308 => x"00039a04",
			309 => x"005304e5",
			310 => x"000004e5",
			311 => x"000004e5",
			312 => x"000004e5",
			313 => x"0003020c",
			314 => x"08025a04",
			315 => x"00000541",
			316 => x"09017d04",
			317 => x"00000541",
			318 => x"00140541",
			319 => x"06018810",
			320 => x"0b07330c",
			321 => x"02093a04",
			322 => x"00000541",
			323 => x"08026f04",
			324 => x"00000541",
			325 => x"ff6d0541",
			326 => x"00000541",
			327 => x"00039a10",
			328 => x"0901fc04",
			329 => x"00000541",
			330 => x"09022808",
			331 => x"0b075f04",
			332 => x"003b0541",
			333 => x"00000541",
			334 => x"00000541",
			335 => x"00000541",
			336 => x"06017718",
			337 => x"0b073314",
			338 => x"0209780c",
			339 => x"0e093308",
			340 => x"0e088e04",
			341 => x"0000059d",
			342 => x"ffec059d",
			343 => x"0000059d",
			344 => x"0b06bc04",
			345 => x"0000059d",
			346 => x"ff8c059d",
			347 => x"0000059d",
			348 => x"0b074414",
			349 => x"0901dd04",
			350 => x"0000059d",
			351 => x"0a027b0c",
			352 => x"0e09a204",
			353 => x"0000059d",
			354 => x"0f0ac304",
			355 => x"0065059d",
			356 => x"0000059d",
			357 => x"0000059d",
			358 => x"0000059d",
			359 => x"0b06dd10",
			360 => x"0e094008",
			361 => x"03097804",
			362 => x"ffc405f1",
			363 => x"000005f1",
			364 => x"0901ee04",
			365 => x"000405f1",
			366 => x"000005f1",
			367 => x"07064604",
			368 => x"000005f1",
			369 => x"040a2814",
			370 => x"0002dd04",
			371 => x"000005f1",
			372 => x"04094504",
			373 => x"000005f1",
			374 => x"0100e704",
			375 => x"000005f1",
			376 => x"0f091f04",
			377 => x"000005f1",
			378 => x"008005f1",
			379 => x"000005f1",
			380 => x"0003701c",
			381 => x"0c05d804",
			382 => x"00000635",
			383 => x"0d087f14",
			384 => x"0d080b04",
			385 => x"00000635",
			386 => x"0a01e904",
			387 => x"00000635",
			388 => x"0b06bf04",
			389 => x"00000635",
			390 => x"0b071e04",
			391 => x"005d0635",
			392 => x"00000635",
			393 => x"00000635",
			394 => x"06018d04",
			395 => x"fff60635",
			396 => x"00000635",
			397 => x"040a2824",
			398 => x"0e09401c",
			399 => x"00030c14",
			400 => x"08025f10",
			401 => x"0d086d0c",
			402 => x"0f08bf04",
			403 => x"00000691",
			404 => x"0d080a04",
			405 => x"00000691",
			406 => x"ffc30691",
			407 => x"00000691",
			408 => x"00520691",
			409 => x"0b06d204",
			410 => x"ff9f0691",
			411 => x"00000691",
			412 => x"03097804",
			413 => x"00000691",
			414 => x"00df0691",
			415 => x"06018808",
			416 => x"0c068904",
			417 => x"ff9e0691",
			418 => x"00000691",
			419 => x"00000691",
			420 => x"05082124",
			421 => x"0507c70c",
			422 => x"0002e604",
			423 => x"000006f5",
			424 => x"02099d04",
			425 => x"ffae06f5",
			426 => x"000006f5",
			427 => x"0c062e14",
			428 => x"06014104",
			429 => x"000006f5",
			430 => x"020a2d0c",
			431 => x"01014308",
			432 => x"00037d04",
			433 => x"00b706f5",
			434 => x"000006f5",
			435 => x"000006f5",
			436 => x"000006f5",
			437 => x"000006f5",
			438 => x"0b07330c",
			439 => x"0e0a3908",
			440 => x"0b06fe04",
			441 => x"000006f5",
			442 => x"ffba06f5",
			443 => x"000006f5",
			444 => x"000006f5",
			445 => x"04098710",
			446 => x"08025a04",
			447 => x"00000759",
			448 => x"0f096008",
			449 => x"0e089604",
			450 => x"00000759",
			451 => x"00330759",
			452 => x"00000759",
			453 => x"06018818",
			454 => x"0b073314",
			455 => x"00030204",
			456 => x"00000759",
			457 => x"0601800c",
			458 => x"0b06bc04",
			459 => x"00000759",
			460 => x"08026f04",
			461 => x"00000759",
			462 => x"ff6a0759",
			463 => x"00000759",
			464 => x"00000759",
			465 => x"00039a08",
			466 => x"01015404",
			467 => x"00220759",
			468 => x"00000759",
			469 => x"00000759",
			470 => x"04091d04",
			471 => x"00000795",
			472 => x"05081f18",
			473 => x"0e098714",
			474 => x"0b071010",
			475 => x"0c05de04",
			476 => x"00000795",
			477 => x"0b06bc04",
			478 => x"00000795",
			479 => x"0309b004",
			480 => x"ff7c0795",
			481 => x"00000795",
			482 => x"00000795",
			483 => x"00000795",
			484 => x"00000795",
			485 => x"0e09871c",
			486 => x"0b072018",
			487 => x"0507e704",
			488 => x"000007d1",
			489 => x"0100e804",
			490 => x"000007d1",
			491 => x"05081f0c",
			492 => x"0a021d08",
			493 => x"07068504",
			494 => x"ff9d07d1",
			495 => x"000007d1",
			496 => x"000007d1",
			497 => x"000007d1",
			498 => x"000007d1",
			499 => x"000007d1",
			500 => x"09017d04",
			501 => x"0000080d",
			502 => x"00037018",
			503 => x"0d087f14",
			504 => x"0d080b04",
			505 => x"0000080d",
			506 => x"0b06bd04",
			507 => x"0000080d",
			508 => x"0a01e404",
			509 => x"0000080d",
			510 => x"0c05d904",
			511 => x"0000080d",
			512 => x"004e080d",
			513 => x"0000080d",
			514 => x"0000080d",
			515 => x"0003891c",
			516 => x"09017a04",
			517 => x"00000849",
			518 => x"07064604",
			519 => x"00000849",
			520 => x"0002e604",
			521 => x"00000849",
			522 => x"0101540c",
			523 => x"0c05dc04",
			524 => x"00000849",
			525 => x"04094504",
			526 => x"00000849",
			527 => x"00630849",
			528 => x"00000849",
			529 => x"00000849",
			530 => x"0100f314",
			531 => x"02092004",
			532 => x"000008a5",
			533 => x"0d086604",
			534 => x"000008a5",
			535 => x"05084d08",
			536 => x"0e092404",
			537 => x"000008a5",
			538 => x"ffa108a5",
			539 => x"000008a5",
			540 => x"00037d18",
			541 => x"0c05f304",
			542 => x"000008a5",
			543 => x"0e093304",
			544 => x"000008a5",
			545 => x"01013d0c",
			546 => x"020a2d08",
			547 => x"0507bb04",
			548 => x"000008a5",
			549 => x"008f08a5",
			550 => x"000008a5",
			551 => x"000008a5",
			552 => x"000008a5",
			553 => x"0409db18",
			554 => x"0f08f904",
			555 => x"00000919",
			556 => x"0309b010",
			557 => x"0a01f204",
			558 => x"00000919",
			559 => x"07064404",
			560 => x"00000919",
			561 => x"0a022804",
			562 => x"00a90919",
			563 => x"00000919",
			564 => x"00000919",
			565 => x"0309d810",
			566 => x"0c05da04",
			567 => x"00000919",
			568 => x"0507ab04",
			569 => x"00000919",
			570 => x"0507f604",
			571 => x"ff890919",
			572 => x"00000919",
			573 => x"01011704",
			574 => x"00000919",
			575 => x"020aa80c",
			576 => x"01015408",
			577 => x"0f0ab604",
			578 => x"00230919",
			579 => x"00000919",
			580 => x"00000919",
			581 => x"00000919",
			582 => x"0b06dd10",
			583 => x"04097204",
			584 => x"00000995",
			585 => x"0e098708",
			586 => x"0507f404",
			587 => x"ff6c0995",
			588 => x"00000995",
			589 => x"00000995",
			590 => x"06014510",
			591 => x"0b06fc04",
			592 => x"00000995",
			593 => x"05082e08",
			594 => x"0c061004",
			595 => x"00000995",
			596 => x"ff680995",
			597 => x"00000995",
			598 => x"040a3a08",
			599 => x"07064604",
			600 => x"00000995",
			601 => x"00c10995",
			602 => x"0901f808",
			603 => x"0b075f04",
			604 => x"ff770995",
			605 => x"00000995",
			606 => x"0101580c",
			607 => x"0d08b308",
			608 => x"0309ef04",
			609 => x"00000995",
			610 => x"00820995",
			611 => x"00000995",
			612 => x"00000995",
			613 => x"0c06132c",
			614 => x"04095910",
			615 => x"0c05d704",
			616 => x"00000a19",
			617 => x"07066c08",
			618 => x"07061304",
			619 => x"00000a19",
			620 => x"00310a19",
			621 => x"00000a19",
			622 => x"0901dd0c",
			623 => x"0507d804",
			624 => x"00000a19",
			625 => x"0e092404",
			626 => x"00000a19",
			627 => x"ff660a19",
			628 => x"0101360c",
			629 => x"0e096204",
			630 => x"00000a19",
			631 => x"0a025904",
			632 => x"003f0a19",
			633 => x"00000a19",
			634 => x"00000a19",
			635 => x"0b070e04",
			636 => x"00000a19",
			637 => x"01015010",
			638 => x"07066e04",
			639 => x"00000a19",
			640 => x"0f0ab208",
			641 => x"00039e04",
			642 => x"00b80a19",
			643 => x"00000a19",
			644 => x"00000a19",
			645 => x"00000a19",
			646 => x"06013e10",
			647 => x"07061304",
			648 => x"00000a95",
			649 => x"07068308",
			650 => x"02092804",
			651 => x"00580a95",
			652 => x"00000a95",
			653 => x"00000a95",
			654 => x"07067024",
			655 => x"0901c310",
			656 => x"0507e704",
			657 => x"00000a95",
			658 => x"0d087208",
			659 => x"0d083804",
			660 => x"00000a95",
			661 => x"ff680a95",
			662 => x"00000a95",
			663 => x"0a025710",
			664 => x"0a021704",
			665 => x"00000a95",
			666 => x"020a2d08",
			667 => x"02091104",
			668 => x"00000a95",
			669 => x"00290a95",
			670 => x"00000a95",
			671 => x"00000a95",
			672 => x"0309ef08",
			673 => x"0802c304",
			674 => x"00600a95",
			675 => x"00000a95",
			676 => x"00000a95",
			677 => x"0c063230",
			678 => x"06018824",
			679 => x"0409db18",
			680 => x"02095110",
			681 => x"0208fe04",
			682 => x"00000b19",
			683 => x"0a021d08",
			684 => x"0f090d04",
			685 => x"00000b19",
			686 => x"ffc00b19",
			687 => x"00000b19",
			688 => x"06014d04",
			689 => x"00000b19",
			690 => x"004e0b19",
			691 => x"07064104",
			692 => x"00000b19",
			693 => x"06015f04",
			694 => x"00000b19",
			695 => x"ff5d0b19",
			696 => x"00038508",
			697 => x"030a1204",
			698 => x"00000b19",
			699 => x"00480b19",
			700 => x"00000b19",
			701 => x"020a8c10",
			702 => x"08025a04",
			703 => x"00000b19",
			704 => x"0706cb08",
			705 => x"01014b04",
			706 => x"008b0b19",
			707 => x"00000b19",
			708 => x"00000b19",
			709 => x"00000b19",
			710 => x"040a0138",
			711 => x"0c061124",
			712 => x"07064010",
			713 => x"07062b04",
			714 => x"00000bb5",
			715 => x"0a021d08",
			716 => x"0408ea04",
			717 => x"00000bb5",
			718 => x"ff9b0bb5",
			719 => x"00000bb5",
			720 => x"06013904",
			721 => x"00000bb5",
			722 => x"0409ed0c",
			723 => x"05082108",
			724 => x"0a01ec04",
			725 => x"00000bb5",
			726 => x"00cb0bb5",
			727 => x"00000bb5",
			728 => x"00000bb5",
			729 => x"0507f40c",
			730 => x"0901c308",
			731 => x"04090804",
			732 => x"00000bb5",
			733 => x"ff6a0bb5",
			734 => x"00000bb5",
			735 => x"0208fe04",
			736 => x"00000bb5",
			737 => x"003f0bb5",
			738 => x"0601770c",
			739 => x"0c063408",
			740 => x"00033504",
			741 => x"00000bb5",
			742 => x"ff570bb5",
			743 => x"00000bb5",
			744 => x"00037008",
			745 => x"0706a104",
			746 => x"00600bb5",
			747 => x"00000bb5",
			748 => x"00000bb5",
			749 => x"040a3a30",
			750 => x"0b071028",
			751 => x"0d084b14",
			752 => x"0d080b04",
			753 => x"00000c29",
			754 => x"09017a04",
			755 => x"00000c29",
			756 => x"0901d708",
			757 => x"0a01e404",
			758 => x"00000c29",
			759 => x"00880c29",
			760 => x"00000c29",
			761 => x"08029110",
			762 => x"0d086d0c",
			763 => x"09017a04",
			764 => x"00000c29",
			765 => x"0208dd04",
			766 => x"00000c29",
			767 => x"ffa90c29",
			768 => x"00000c29",
			769 => x"00000c29",
			770 => x"0309ef04",
			771 => x"005f0c29",
			772 => x"00000c29",
			773 => x"0c063408",
			774 => x"030a8104",
			775 => x"ffae0c29",
			776 => x"00000c29",
			777 => x"00000c29",
			778 => x"0b06dd14",
			779 => x"00030c0c",
			780 => x"0c061208",
			781 => x"0c05ba04",
			782 => x"00000cc5",
			783 => x"001c0cc5",
			784 => x"00000cc5",
			785 => x"0e098704",
			786 => x"ff860cc5",
			787 => x"00000cc5",
			788 => x"06014114",
			789 => x"0e092410",
			790 => x"0d083e04",
			791 => x"00000cc5",
			792 => x"0c05f304",
			793 => x"00000cc5",
			794 => x"0e08cb04",
			795 => x"00000cc5",
			796 => x"ff640cc5",
			797 => x"00000cc5",
			798 => x"040a3a0c",
			799 => x"09017d04",
			800 => x"00000cc5",
			801 => x"07064604",
			802 => x"00000cc5",
			803 => x"00b80cc5",
			804 => x"0901fc0c",
			805 => x"0b075f08",
			806 => x"0901f804",
			807 => x"ff900cc5",
			808 => x"00000cc5",
			809 => x"00000cc5",
			810 => x"0101580c",
			811 => x"0d08b308",
			812 => x"00039a04",
			813 => x"007b0cc5",
			814 => x"00000cc5",
			815 => x"00000cc5",
			816 => x"00000cc5",
			817 => x"0003242c",
			818 => x"0e097724",
			819 => x"0c05d704",
			820 => x"00000d61",
			821 => x"0a01f210",
			822 => x"09018008",
			823 => x"03096804",
			824 => x"005a0d61",
			825 => x"00000d61",
			826 => x"0208c904",
			827 => x"00000d61",
			828 => x"ffe30d61",
			829 => x"0507b804",
			830 => x"00000d61",
			831 => x"07063d04",
			832 => x"00000d61",
			833 => x"0309c004",
			834 => x"00ed0d61",
			835 => x"00000d61",
			836 => x"0c062e04",
			837 => x"ffe60d61",
			838 => x"00000d61",
			839 => x"06017710",
			840 => x"040a0108",
			841 => x"0409c704",
			842 => x"fff00d61",
			843 => x"00000d61",
			844 => x"0c063404",
			845 => x"ff0b0d61",
			846 => x"00000d61",
			847 => x"0c063a10",
			848 => x"040b220c",
			849 => x"0c05f604",
			850 => x"00000d61",
			851 => x"0a027704",
			852 => x"00360d61",
			853 => x"00000d61",
			854 => x"00000d61",
			855 => x"00000d61",
			856 => x"00039a28",
			857 => x"0c05ba04",
			858 => x"fe2d0db5",
			859 => x"05088620",
			860 => x"0e0a2a14",
			861 => x"09017a08",
			862 => x"02080004",
			863 => x"01b90db5",
			864 => x"fe620db5",
			865 => x"00037d08",
			866 => x"0c063204",
			867 => x"00a10db5",
			868 => x"01af0db5",
			869 => x"fe820db5",
			870 => x"00039208",
			871 => x"0802e204",
			872 => x"00600db5",
			873 => x"02780db5",
			874 => x"04890db5",
			875 => x"fe8e0db5",
			876 => x"fe660db5",
			877 => x"0409a020",
			878 => x"0c05d704",
			879 => x"00000e61",
			880 => x"07066c0c",
			881 => x"01011108",
			882 => x"0100eb04",
			883 => x"00000e61",
			884 => x"00f00e61",
			885 => x"00000e61",
			886 => x"0002e608",
			887 => x"0002dd04",
			888 => x"00000e61",
			889 => x"ffb70e61",
			890 => x"0002ee04",
			891 => x"00000e61",
			892 => x"00460e61",
			893 => x"03097810",
			894 => x"0c06130c",
			895 => x"07065908",
			896 => x"0e096204",
			897 => x"fee70e61",
			898 => x"00000e61",
			899 => x"00000e61",
			900 => x"00000e61",
			901 => x"02099508",
			902 => x"0100f304",
			903 => x"00000e61",
			904 => x"00e40e61",
			905 => x"0e09870c",
			906 => x"0c061208",
			907 => x"07064104",
			908 => x"00000e61",
			909 => x"ff100e61",
			910 => x"00000e61",
			911 => x"0209c104",
			912 => x"009b0e61",
			913 => x"01012e08",
			914 => x"0706c904",
			915 => x"ff5b0e61",
			916 => x"00000e61",
			917 => x"01014504",
			918 => x"00420e61",
			919 => x"ffc40e61",
			920 => x"00039a28",
			921 => x"0c05ba04",
			922 => x"fe2e0eb5",
			923 => x"0d08f420",
			924 => x"0e0a2a18",
			925 => x"09017a08",
			926 => x"0a01b604",
			927 => x"01f00eb5",
			928 => x"fe5c0eb5",
			929 => x"0c063208",
			930 => x"0d088d04",
			931 => x"00c00eb5",
			932 => x"fefe0eb5",
			933 => x"01014504",
			934 => x"01c10eb5",
			935 => x"ff8f0eb5",
			936 => x"00039204",
			937 => x"026d0eb5",
			938 => x"04e60eb5",
			939 => x"fe790eb5",
			940 => x"fe660eb5",
			941 => x"040abb3c",
			942 => x"09017a10",
			943 => x"0b07010c",
			944 => x"0600ef08",
			945 => x"0801be04",
			946 => x"fe7e0f51",
			947 => x"01ef0f51",
			948 => x"fe610f51",
			949 => x"00000f51",
			950 => x"0d07fd08",
			951 => x"06015604",
			952 => x"00f10f51",
			953 => x"fe720f51",
			954 => x"0d08da1c",
			955 => x"0e09fd10",
			956 => x"040a3a08",
			957 => x"0a01e904",
			958 => x"00bd0f51",
			959 => x"02120f51",
			960 => x"0e09a204",
			961 => x"fd940f51",
			962 => x"01d90f51",
			963 => x"07066e08",
			964 => x"0802e004",
			965 => x"02f00f51",
			966 => x"00000f51",
			967 => x"03f30f51",
			968 => x"0c06a604",
			969 => x"fe410f51",
			970 => x"00c20f51",
			971 => x"040b2210",
			972 => x"06019404",
			973 => x"fe680f51",
			974 => x"05081f04",
			975 => x"fe8c0f51",
			976 => x"01015b04",
			977 => x"033f0f51",
			978 => x"fec10f51",
			979 => x"fe610f51",
			980 => x"00036340",
			981 => x"06016230",
			982 => x"01010f24",
			983 => x"03095810",
			984 => x"06013804",
			985 => x"00000fdd",
			986 => x"04098708",
			987 => x"0a01e404",
			988 => x"00000fdd",
			989 => x"00940fdd",
			990 => x"00000fdd",
			991 => x"0c06320c",
			992 => x"06013e04",
			993 => x"00000fdd",
			994 => x"01010604",
			995 => x"ff940fdd",
			996 => x"00000fdd",
			997 => x"0f093d04",
			998 => x"00000fdd",
			999 => x"005e0fdd",
			1000 => x"0a021708",
			1001 => x"07062b04",
			1002 => x"00000fdd",
			1003 => x"ff4f0fdd",
			1004 => x"00000fdd",
			1005 => x"0901b804",
			1006 => x"00000fdd",
			1007 => x"0c05f304",
			1008 => x"00000fdd",
			1009 => x"03094f04",
			1010 => x"00000fdd",
			1011 => x"01100fdd",
			1012 => x"06018c04",
			1013 => x"ff2d0fdd",
			1014 => x"00000fdd",
			1015 => x"0f092a0c",
			1016 => x"04091d04",
			1017 => x"00001089",
			1018 => x"08025a04",
			1019 => x"ff3f1089",
			1020 => x"00001089",
			1021 => x"040a3a20",
			1022 => x"0a021714",
			1023 => x"05081f0c",
			1024 => x"02092004",
			1025 => x"00001089",
			1026 => x"0507e704",
			1027 => x"00001089",
			1028 => x"ff5f1089",
			1029 => x"0100eb04",
			1030 => x"00001089",
			1031 => x"008b1089",
			1032 => x"00035308",
			1033 => x"0d080e04",
			1034 => x"00001089",
			1035 => x"010e1089",
			1036 => x"00001089",
			1037 => x"0209e80c",
			1038 => x"06018008",
			1039 => x"07062e04",
			1040 => x"00001089",
			1041 => x"ff2a1089",
			1042 => x"00001089",
			1043 => x"00037d10",
			1044 => x"07064004",
			1045 => x"00001089",
			1046 => x"040ac908",
			1047 => x"01014b04",
			1048 => x"009d1089",
			1049 => x"00001089",
			1050 => x"00001089",
			1051 => x"06019404",
			1052 => x"ffb41089",
			1053 => x"040b2208",
			1054 => x"09020e04",
			1055 => x"00001089",
			1056 => x"00371089",
			1057 => x"00001089",
			1058 => x"0409a030",
			1059 => x"01010f24",
			1060 => x"03098720",
			1061 => x"0a01e910",
			1062 => x"03091a0c",
			1063 => x"0307f404",
			1064 => x"0000114d",
			1065 => x"0507e604",
			1066 => x"002b114d",
			1067 => x"0000114d",
			1068 => x"0000114d",
			1069 => x"07062804",
			1070 => x"0000114d",
			1071 => x"0100e704",
			1072 => x"0000114d",
			1073 => x"0002d504",
			1074 => x"0000114d",
			1075 => x"00d4114d",
			1076 => x"0000114d",
			1077 => x"0b06cd08",
			1078 => x"0a021704",
			1079 => x"ffc8114d",
			1080 => x"0000114d",
			1081 => x"0000114d",
			1082 => x"06018820",
			1083 => x"040a0114",
			1084 => x"0a021d0c",
			1085 => x"0b070e08",
			1086 => x"0507d804",
			1087 => x"0000114d",
			1088 => x"ff4d114d",
			1089 => x"0000114d",
			1090 => x"03095804",
			1091 => x"0000114d",
			1092 => x"0068114d",
			1093 => x"0b074408",
			1094 => x"06017704",
			1095 => x"fefa114d",
			1096 => x"0000114d",
			1097 => x"0000114d",
			1098 => x"0901fc04",
			1099 => x"0000114d",
			1100 => x"00039a0c",
			1101 => x"0b074408",
			1102 => x"0b06dd04",
			1103 => x"0000114d",
			1104 => x"006e114d",
			1105 => x"0000114d",
			1106 => x"0000114d",
			1107 => x"0c05f61c",
			1108 => x"0e098710",
			1109 => x"0003240c",
			1110 => x"0a021708",
			1111 => x"08026f04",
			1112 => x"000011f9",
			1113 => x"ffa811f9",
			1114 => x"000011f9",
			1115 => x"fedb11f9",
			1116 => x"00037808",
			1117 => x"0901dd04",
			1118 => x"000011f9",
			1119 => x"004611f9",
			1120 => x"000011f9",
			1121 => x"00038538",
			1122 => x"0e09331c",
			1123 => x"0507f610",
			1124 => x"04091d04",
			1125 => x"000011f9",
			1126 => x"0b06bd04",
			1127 => x"000011f9",
			1128 => x"0507f404",
			1129 => x"ff6d11f9",
			1130 => x"000011f9",
			1131 => x"0a01e904",
			1132 => x"000011f9",
			1133 => x"02092804",
			1134 => x"009411f9",
			1135 => x"000011f9",
			1136 => x"0100f308",
			1137 => x"0309c004",
			1138 => x"000011f9",
			1139 => x"ffff11f9",
			1140 => x"01013d08",
			1141 => x"00036304",
			1142 => x"010211f9",
			1143 => x"000011f9",
			1144 => x"0507ea04",
			1145 => x"fff411f9",
			1146 => x"05084d04",
			1147 => x"004711f9",
			1148 => x"000011f9",
			1149 => x"ffcc11f9",
			1150 => x"0f092a0c",
			1151 => x"04091d04",
			1152 => x"000012ad",
			1153 => x"08025a04",
			1154 => x"ff5012ad",
			1155 => x"000012ad",
			1156 => x"040a3a20",
			1157 => x"06016214",
			1158 => x"0b06ec08",
			1159 => x"0507e704",
			1160 => x"000012ad",
			1161 => x"ff4312ad",
			1162 => x"0002e604",
			1163 => x"000012ad",
			1164 => x"0d085704",
			1165 => x"000012ad",
			1166 => x"009712ad",
			1167 => x"00035308",
			1168 => x"0d080e04",
			1169 => x"000012ad",
			1170 => x"00f312ad",
			1171 => x"000012ad",
			1172 => x"0209e810",
			1173 => x"0601800c",
			1174 => x"07062e04",
			1175 => x"000012ad",
			1176 => x"0b06cf04",
			1177 => x"000012ad",
			1178 => x"ff3312ad",
			1179 => x"000012ad",
			1180 => x"00037d10",
			1181 => x"07064004",
			1182 => x"000012ad",
			1183 => x"040ac908",
			1184 => x"01014b04",
			1185 => x"009612ad",
			1186 => x"000012ad",
			1187 => x"000012ad",
			1188 => x"06019404",
			1189 => x"ffbf12ad",
			1190 => x"020aa808",
			1191 => x"01014904",
			1192 => x"000012ad",
			1193 => x"002b12ad",
			1194 => x"000012ad",
			1195 => x"00038944",
			1196 => x"0100e710",
			1197 => x"0600ef08",
			1198 => x"09010a04",
			1199 => x"feba1349",
			1200 => x"02181349",
			1201 => x"09017a04",
			1202 => x"fe5b1349",
			1203 => x"00001349",
			1204 => x"0d08da2c",
			1205 => x"07064014",
			1206 => x"00035b10",
			1207 => x"0c05f608",
			1208 => x"02091904",
			1209 => x"00d61349",
			1210 => x"fef51349",
			1211 => x"0b06a504",
			1212 => x"00001349",
			1213 => x"019e1349",
			1214 => x"fe641349",
			1215 => x"030a1210",
			1216 => x"00036308",
			1217 => x"01013904",
			1218 => x"014b1349",
			1219 => x"ff6b1349",
			1220 => x"0b06e004",
			1221 => x"fe361349",
			1222 => x"00001349",
			1223 => x"06018d04",
			1224 => x"01be1349",
			1225 => x"02991349",
			1226 => x"07072404",
			1227 => x"fe711349",
			1228 => x"00cc1349",
			1229 => x"00039608",
			1230 => x"06019404",
			1231 => x"fe751349",
			1232 => x"02671349",
			1233 => x"fe651349",
			1234 => x"00038940",
			1235 => x"030a1230",
			1236 => x"00035328",
			1237 => x"06016f20",
			1238 => x"02093a10",
			1239 => x"0100eb08",
			1240 => x"0002cc04",
			1241 => x"000013d5",
			1242 => x"ff2813d5",
			1243 => x"0b070e04",
			1244 => x"00ab13d5",
			1245 => x"ffea13d5",
			1246 => x"0c061308",
			1247 => x"0c05de04",
			1248 => x"000013d5",
			1249 => x"ff2e13d5",
			1250 => x"01010204",
			1251 => x"ffbd13d5",
			1252 => x"00e313d5",
			1253 => x"03097804",
			1254 => x"000013d5",
			1255 => x"016513d5",
			1256 => x"0309ef04",
			1257 => x"fea113d5",
			1258 => x"000013d5",
			1259 => x"020a2d04",
			1260 => x"013413d5",
			1261 => x"0d088d04",
			1262 => x"004b13d5",
			1263 => x"020a5b04",
			1264 => x"ffb313d5",
			1265 => x"000013d5",
			1266 => x"09021504",
			1267 => x"fe8d13d5",
			1268 => x"000013d5",
			1269 => x"040abb3c",
			1270 => x"09017a10",
			1271 => x"0e09070c",
			1272 => x"0600ef08",
			1273 => x"0600ee04",
			1274 => x"fe6f14b9",
			1275 => x"01b514b9",
			1276 => x"fe5d14b9",
			1277 => x"016d14b9",
			1278 => x"0d080e0c",
			1279 => x"01010f08",
			1280 => x"04098704",
			1281 => x"035114b9",
			1282 => x"feea14b9",
			1283 => x"fe5a14b9",
			1284 => x"01014518",
			1285 => x"0a01e408",
			1286 => x"0507e604",
			1287 => x"021014b9",
			1288 => x"fe6614b9",
			1289 => x"040a9508",
			1290 => x"0100e704",
			1291 => x"000014b9",
			1292 => x"036b14b9",
			1293 => x"030a1204",
			1294 => x"febc14b9",
			1295 => x"078614b9",
			1296 => x"0c061204",
			1297 => x"00e114b9",
			1298 => x"fe6e14b9",
			1299 => x"040af718",
			1300 => x"06019410",
			1301 => x"06019108",
			1302 => x"040ac204",
			1303 => x"fef314b9",
			1304 => x"fe5c14b9",
			1305 => x"040ae204",
			1306 => x"00ff14b9",
			1307 => x"feb414b9",
			1308 => x"030a4904",
			1309 => x"fe8514b9",
			1310 => x"066514b9",
			1311 => x"040b221c",
			1312 => x"040b1c10",
			1313 => x"0802f804",
			1314 => x"fe5e14b9",
			1315 => x"08030208",
			1316 => x"0802fb04",
			1317 => x"00d214b9",
			1318 => x"fffa14b9",
			1319 => x"fe6514b9",
			1320 => x"0802f104",
			1321 => x"fe8014b9",
			1322 => x"01013a04",
			1323 => x"fe9a14b9",
			1324 => x"046e14b9",
			1325 => x"fe5c14b9",
			1326 => x"00037044",
			1327 => x"03094f1c",
			1328 => x"0901800c",
			1329 => x"09017a04",
			1330 => x"c96a15ad",
			1331 => x"0a01e404",
			1332 => x"c9c015ad",
			1333 => x"d32215ad",
			1334 => x"00030208",
			1335 => x"0c061704",
			1336 => x"f60915ad",
			1337 => x"e51015ad",
			1338 => x"0d081704",
			1339 => x"c96515ad",
			1340 => x"dd1915ad",
			1341 => x"0d081808",
			1342 => x"0d080e04",
			1343 => x"c98415ad",
			1344 => x"d52215ad",
			1345 => x"09018010",
			1346 => x"06014108",
			1347 => x"08025a04",
			1348 => x"c98a15ad",
			1349 => x"d42f15ad",
			1350 => x"07066e04",
			1351 => x"cffe15ad",
			1352 => x"e89515ad",
			1353 => x"0101450c",
			1354 => x"040a9508",
			1355 => x"08025f04",
			1356 => x"e70115ad",
			1357 => x"f4de15ad",
			1358 => x"e0d515ad",
			1359 => x"c9a815ad",
			1360 => x"00037d18",
			1361 => x"0802db14",
			1362 => x"0601880c",
			1363 => x"06018304",
			1364 => x"c96c15ad",
			1365 => x"040aa904",
			1366 => x"cd2b15ad",
			1367 => x"c9d315ad",
			1368 => x"01015304",
			1369 => x"d52215ad",
			1370 => x"c9db15ad",
			1371 => x"e90c15ad",
			1372 => x"00039518",
			1373 => x"06019914",
			1374 => x"0802e90c",
			1375 => x"0802e504",
			1376 => x"c96215ad",
			1377 => x"040ae204",
			1378 => x"cd2b15ad",
			1379 => x"c97c15ad",
			1380 => x"01015904",
			1381 => x"d91d15ad",
			1382 => x"c9fb15ad",
			1383 => x"ed0715ad",
			1384 => x"00039a04",
			1385 => x"c9a915ad",
			1386 => x"c96015ad",
			1387 => x"0901dd50",
			1388 => x"0003243c",
			1389 => x"0507e718",
			1390 => x"08025a10",
			1391 => x"0901900c",
			1392 => x"0c05f204",
			1393 => x"000016a9",
			1394 => x"03093704",
			1395 => x"004416a9",
			1396 => x"000016a9",
			1397 => x"ffa816a9",
			1398 => x"0507b804",
			1399 => x"000016a9",
			1400 => x"00fc16a9",
			1401 => x"0507f60c",
			1402 => x"0f096808",
			1403 => x"06014104",
			1404 => x"000016a9",
			1405 => x"000616a9",
			1406 => x"ff1416a9",
			1407 => x"0100f110",
			1408 => x"03096808",
			1409 => x"09018004",
			1410 => x"008b16a9",
			1411 => x"000016a9",
			1412 => x"07068504",
			1413 => x"ff6716a9",
			1414 => x"000016a9",
			1415 => x"08028704",
			1416 => x"007716a9",
			1417 => x"000016a9",
			1418 => x"0c05fa08",
			1419 => x"01012a04",
			1420 => x"fefa16a9",
			1421 => x"000016a9",
			1422 => x"01010204",
			1423 => x"fff516a9",
			1424 => x"0901cc04",
			1425 => x"004f16a9",
			1426 => x"000016a9",
			1427 => x"00036810",
			1428 => x"06016f04",
			1429 => x"000016a9",
			1430 => x"03098704",
			1431 => x"000016a9",
			1432 => x"05083004",
			1433 => x"010a16a9",
			1434 => x"000016a9",
			1435 => x"0e0a1b0c",
			1436 => x"0c05f404",
			1437 => x"000016a9",
			1438 => x"030a5c04",
			1439 => x"ff7716a9",
			1440 => x"000016a9",
			1441 => x"0f0ac310",
			1442 => x"06018d04",
			1443 => x"000016a9",
			1444 => x"05080104",
			1445 => x"000016a9",
			1446 => x"0a027704",
			1447 => x"00da16a9",
			1448 => x"000016a9",
			1449 => x"000016a9",
			1450 => x"0c05d80c",
			1451 => x"0e098708",
			1452 => x"0507c704",
			1453 => x"ff0c1775",
			1454 => x"00001775",
			1455 => x"00001775",
			1456 => x"0c061a30",
			1457 => x"05081220",
			1458 => x"0901db0c",
			1459 => x"00034608",
			1460 => x"07068304",
			1461 => x"00e01775",
			1462 => x"00001775",
			1463 => x"00001775",
			1464 => x"06017008",
			1465 => x"0901e804",
			1466 => x"ff621775",
			1467 => x"00001775",
			1468 => x"00037d08",
			1469 => x"06018904",
			1470 => x"00d31775",
			1471 => x"00001775",
			1472 => x"00001775",
			1473 => x"09019c08",
			1474 => x"03097804",
			1475 => x"00001775",
			1476 => x"ff901775",
			1477 => x"00039604",
			1478 => x"006f1775",
			1479 => x"00001775",
			1480 => x"05080f08",
			1481 => x"07066d04",
			1482 => x"ff661775",
			1483 => x"00001775",
			1484 => x"0c063214",
			1485 => x"0c062e0c",
			1486 => x"05083e08",
			1487 => x"0d087f04",
			1488 => x"00321775",
			1489 => x"00001775",
			1490 => x"00001775",
			1491 => x"020a4604",
			1492 => x"ffbb1775",
			1493 => x"00001775",
			1494 => x"020a8c0c",
			1495 => x"0f093d04",
			1496 => x"00001775",
			1497 => x"040af704",
			1498 => x"00af1775",
			1499 => x"00001775",
			1500 => x"00001775",
			1501 => x"0c05f624",
			1502 => x"0409720c",
			1503 => x"0e078e04",
			1504 => x"00001871",
			1505 => x"02090004",
			1506 => x"00101871",
			1507 => x"00001871",
			1508 => x"0901e30c",
			1509 => x"00032408",
			1510 => x"00030c04",
			1511 => x"ff671871",
			1512 => x"00001871",
			1513 => x"feb71871",
			1514 => x"00037808",
			1515 => x"0e098704",
			1516 => x"00001871",
			1517 => x"00681871",
			1518 => x"00001871",
			1519 => x"06013e18",
			1520 => x"02090010",
			1521 => x"03092e0c",
			1522 => x"0308bf04",
			1523 => x"00001871",
			1524 => x"0d083f04",
			1525 => x"00211871",
			1526 => x"00001871",
			1527 => x"fff31871",
			1528 => x"0d086d04",
			1529 => x"00001871",
			1530 => x"00e51871",
			1531 => x"0c05f810",
			1532 => x"0601890c",
			1533 => x"00038108",
			1534 => x"0d07fd04",
			1535 => x"00001871",
			1536 => x"00de1871",
			1537 => x"00001871",
			1538 => x"00001871",
			1539 => x"0507f414",
			1540 => x"0901a108",
			1541 => x"09017d04",
			1542 => x"00001871",
			1543 => x"00041871",
			1544 => x"0a021704",
			1545 => x"fedd1871",
			1546 => x"0901f004",
			1547 => x"00071871",
			1548 => x"ff9a1871",
			1549 => x"0100ff10",
			1550 => x"06015208",
			1551 => x"0c063204",
			1552 => x"ffe91871",
			1553 => x"00a01871",
			1554 => x"0309ef04",
			1555 => x"00001871",
			1556 => x"ff5c1871",
			1557 => x"00037808",
			1558 => x"030a7804",
			1559 => x"00f91871",
			1560 => x"00001871",
			1561 => x"0e0a2a04",
			1562 => x"ff731871",
			1563 => x"00211871",
			1564 => x"0c05dc18",
			1565 => x"00034614",
			1566 => x"02093a0c",
			1567 => x"0c05d708",
			1568 => x"07064304",
			1569 => x"ff71195d",
			1570 => x"0000195d",
			1571 => x"0000195d",
			1572 => x"0d081704",
			1573 => x"0000195d",
			1574 => x"00d6195d",
			1575 => x"fe88195d",
			1576 => x"0c061338",
			1577 => x"0508122c",
			1578 => x"01013d20",
			1579 => x"0d082210",
			1580 => x"0507ad08",
			1581 => x"00033e04",
			1582 => x"0100195d",
			1583 => x"0000195d",
			1584 => x"0507ba04",
			1585 => x"feda195d",
			1586 => x"0000195d",
			1587 => x"0d085908",
			1588 => x"06013d04",
			1589 => x"0000195d",
			1590 => x"0133195d",
			1591 => x"0507f404",
			1592 => x"ff7b195d",
			1593 => x"0034195d",
			1594 => x"0d085708",
			1595 => x"0c05f404",
			1596 => x"0000195d",
			1597 => x"ff34195d",
			1598 => x"0000195d",
			1599 => x"03097804",
			1600 => x"0000195d",
			1601 => x"09019c04",
			1602 => x"fec8195d",
			1603 => x"0000195d",
			1604 => x"0209000c",
			1605 => x"0100ef08",
			1606 => x"04090804",
			1607 => x"0000195d",
			1608 => x"ffc0195d",
			1609 => x"0000195d",
			1610 => x"0c064d10",
			1611 => x"0902290c",
			1612 => x"0100e704",
			1613 => x"0000195d",
			1614 => x"00039a04",
			1615 => x"0135195d",
			1616 => x"0000195d",
			1617 => x"0000195d",
			1618 => x"0802b708",
			1619 => x"07068504",
			1620 => x"0000195d",
			1621 => x"00a2195d",
			1622 => x"ffc9195d",
			1623 => x"0901dd50",
			1624 => x"0409db40",
			1625 => x"0507ea20",
			1626 => x"0d082514",
			1627 => x"01010f08",
			1628 => x"0c05d704",
			1629 => x"00001a69",
			1630 => x"00081a69",
			1631 => x"0a021d08",
			1632 => x"0c05db04",
			1633 => x"00001a69",
			1634 => x"ff691a69",
			1635 => x"00001a69",
			1636 => x"06013d04",
			1637 => x"00001a69",
			1638 => x"0208d004",
			1639 => x"00001a69",
			1640 => x"00c71a69",
			1641 => x"07065b0c",
			1642 => x"06015208",
			1643 => x"03092e04",
			1644 => x"00001a69",
			1645 => x"ff281a69",
			1646 => x"00001a69",
			1647 => x"07066c08",
			1648 => x"02090904",
			1649 => x"00001a69",
			1650 => x"006a1a69",
			1651 => x"03094f04",
			1652 => x"00001a69",
			1653 => x"07068504",
			1654 => x"ffb01a69",
			1655 => x"00001a69",
			1656 => x"0c064d0c",
			1657 => x"0901d908",
			1658 => x"08028704",
			1659 => x"00001a69",
			1660 => x"feed1a69",
			1661 => x"00001a69",
			1662 => x"00001a69",
			1663 => x"07065818",
			1664 => x"06016f04",
			1665 => x"00001a69",
			1666 => x"020a2d10",
			1667 => x"03099604",
			1668 => x"00001a69",
			1669 => x"0a025b08",
			1670 => x"0d081704",
			1671 => x"00001a69",
			1672 => x"00ee1a69",
			1673 => x"00001a69",
			1674 => x"00001a69",
			1675 => x"0e0a1b0c",
			1676 => x"040a0104",
			1677 => x"00001a69",
			1678 => x"030a5c04",
			1679 => x"ffc91a69",
			1680 => x"00001a69",
			1681 => x"0f0ac310",
			1682 => x"05080f04",
			1683 => x"00001a69",
			1684 => x"0706b708",
			1685 => x"0c064d04",
			1686 => x"004e1a69",
			1687 => x"00001a69",
			1688 => x"00001a69",
			1689 => x"00001a69",
			1690 => x"00039a40",
			1691 => x"0c05d50c",
			1692 => x"07064104",
			1693 => x"fe601aed",
			1694 => x"06013904",
			1695 => x"00001aed",
			1696 => x"00211aed",
			1697 => x"0a026d30",
			1698 => x"0003531c",
			1699 => x"06016610",
			1700 => x"00032408",
			1701 => x"0b071004",
			1702 => x"00751aed",
			1703 => x"01a11aed",
			1704 => x"0c061004",
			1705 => x"fd941aed",
			1706 => x"ffa11aed",
			1707 => x"0e096208",
			1708 => x"01012504",
			1709 => x"01421aed",
			1710 => x"fe9e1aed",
			1711 => x"01d61aed",
			1712 => x"0309d804",
			1713 => x"fdeb1aed",
			1714 => x"01014508",
			1715 => x"00038904",
			1716 => x"017e1aed",
			1717 => x"ff151aed",
			1718 => x"0a026504",
			1719 => x"feb11aed",
			1720 => x"00171aed",
			1721 => x"034b1aed",
			1722 => x"fe691aed",
			1723 => x"0c05d808",
			1724 => x"00034604",
			1725 => x"00001bb9",
			1726 => x"ff021bb9",
			1727 => x"0c061a30",
			1728 => x"0b071e28",
			1729 => x"07064018",
			1730 => x"07062c0c",
			1731 => x"00035308",
			1732 => x"07061304",
			1733 => x"00001bb9",
			1734 => x"00ae1bb9",
			1735 => x"00001bb9",
			1736 => x"0a021d08",
			1737 => x"0f091f04",
			1738 => x"00001bb9",
			1739 => x"ff261bb9",
			1740 => x"00001bb9",
			1741 => x"0003890c",
			1742 => x"06013d04",
			1743 => x"00001bb9",
			1744 => x"0100e804",
			1745 => x"00001bb9",
			1746 => x"01021bb9",
			1747 => x"00001bb9",
			1748 => x"09019c04",
			1749 => x"ff981bb9",
			1750 => x"00001bb9",
			1751 => x"0b070e0c",
			1752 => x"06018d08",
			1753 => x"0c063204",
			1754 => x"ff2f1bb9",
			1755 => x"00001bb9",
			1756 => x"00001bb9",
			1757 => x"0d08b310",
			1758 => x"07066e04",
			1759 => x"00001bb9",
			1760 => x"0c065008",
			1761 => x"0003aa04",
			1762 => x"00e11bb9",
			1763 => x"00001bb9",
			1764 => x"00001bb9",
			1765 => x"0706b708",
			1766 => x"09022104",
			1767 => x"ff801bb9",
			1768 => x"00001bb9",
			1769 => x"01012308",
			1770 => x"0b079304",
			1771 => x"00411bb9",
			1772 => x"00001bb9",
			1773 => x"00001bb9",
			1774 => x"00039a44",
			1775 => x"0c05d50c",
			1776 => x"07064104",
			1777 => x"fe581c45",
			1778 => x"06013904",
			1779 => x"00001c45",
			1780 => x"00281c45",
			1781 => x"0a026d34",
			1782 => x"0d089a20",
			1783 => x"0b06ee10",
			1784 => x"00035308",
			1785 => x"0d084b04",
			1786 => x"01341c45",
			1787 => x"ff4b1c45",
			1788 => x"0d084a04",
			1789 => x"fe351c45",
			1790 => x"011d1c45",
			1791 => x"0002dd08",
			1792 => x"06014104",
			1793 => x"fe261c45",
			1794 => x"00551c45",
			1795 => x"03097804",
			1796 => x"02361c45",
			1797 => x"00e81c45",
			1798 => x"040a2808",
			1799 => x"07068604",
			1800 => x"00001c45",
			1801 => x"01751c45",
			1802 => x"07072508",
			1803 => x"0a026404",
			1804 => x"fe371c45",
			1805 => x"fff11c45",
			1806 => x"00841c45",
			1807 => x"03c91c45",
			1808 => x"fe681c45",
			1809 => x"07063f10",
			1810 => x"0002ee04",
			1811 => x"00001d39",
			1812 => x"03098708",
			1813 => x"0c061004",
			1814 => x"febb1d39",
			1815 => x"00001d39",
			1816 => x"00001d39",
			1817 => x"07067048",
			1818 => x"0507e724",
			1819 => x"0e08d608",
			1820 => x"01010f04",
			1821 => x"00001d39",
			1822 => x"ff351d39",
			1823 => x"0101260c",
			1824 => x"00034b08",
			1825 => x"0a01e404",
			1826 => x"00001d39",
			1827 => x"00f41d39",
			1828 => x"00001d39",
			1829 => x"0309b008",
			1830 => x"040a0104",
			1831 => x"00001d39",
			1832 => x"ff461d39",
			1833 => x"0a025704",
			1834 => x"00ca1d39",
			1835 => x"00001d39",
			1836 => x"0f094514",
			1837 => x"0e09070c",
			1838 => x"0a01ec08",
			1839 => x"03092204",
			1840 => x"00001d39",
			1841 => x"ffaf1d39",
			1842 => x"00001d39",
			1843 => x"03097804",
			1844 => x"00ba1d39",
			1845 => x"00001d39",
			1846 => x"0c06300c",
			1847 => x"0c05da04",
			1848 => x"00001d39",
			1849 => x"07064404",
			1850 => x"00001d39",
			1851 => x"ff301d39",
			1852 => x"00001d39",
			1853 => x"0309ef10",
			1854 => x"0002dd04",
			1855 => x"00001d39",
			1856 => x"040a5b08",
			1857 => x"07067104",
			1858 => x"00001d39",
			1859 => x"012a1d39",
			1860 => x"00001d39",
			1861 => x"01010604",
			1862 => x"ff9c1d39",
			1863 => x"020a8c0c",
			1864 => x"01015608",
			1865 => x"030a3904",
			1866 => x"00001d39",
			1867 => x"00b91d39",
			1868 => x"00001d39",
			1869 => x"00001d39",
			1870 => x"07063f10",
			1871 => x"04097204",
			1872 => x"00001e35",
			1873 => x"02095708",
			1874 => x"0c05f904",
			1875 => x"fee31e35",
			1876 => x"00001e35",
			1877 => x"00001e35",
			1878 => x"06016640",
			1879 => x"0409c730",
			1880 => x"0a01f21c",
			1881 => x"0100e90c",
			1882 => x"06013e08",
			1883 => x"0c061004",
			1884 => x"00001e35",
			1885 => x"00811e35",
			1886 => x"00001e35",
			1887 => x"06014008",
			1888 => x"0e08cb04",
			1889 => x"00001e35",
			1890 => x"ff2e1e35",
			1891 => x"03092204",
			1892 => x"ffbb1e35",
			1893 => x"00461e35",
			1894 => x"0b06d20c",
			1895 => x"0f095608",
			1896 => x"0100fc04",
			1897 => x"00001e35",
			1898 => x"00171e35",
			1899 => x"ffc21e35",
			1900 => x"0100ed04",
			1901 => x"00001e35",
			1902 => x"00fc1e35",
			1903 => x"0706a10c",
			1904 => x"0507ea04",
			1905 => x"00001e35",
			1906 => x"0c063a04",
			1907 => x"fee91e35",
			1908 => x"00001e35",
			1909 => x"00011e35",
			1910 => x"00035310",
			1911 => x"0101380c",
			1912 => x"0c05f304",
			1913 => x"00001e35",
			1914 => x"03094f04",
			1915 => x"00001e35",
			1916 => x"01151e35",
			1917 => x"00001e35",
			1918 => x"01013808",
			1919 => x"0c06e504",
			1920 => x"ff7e1e35",
			1921 => x"00001e35",
			1922 => x"0101450c",
			1923 => x"0a026708",
			1924 => x"0507d904",
			1925 => x"00001e35",
			1926 => x"00c21e35",
			1927 => x"00001e35",
			1928 => x"0a026504",
			1929 => x"ff741e35",
			1930 => x"040b2204",
			1931 => x"00721e35",
			1932 => x"00001e35",
			1933 => x"09017a10",
			1934 => x"0801cb0c",
			1935 => x"0406a304",
			1936 => x"00001f11",
			1937 => x"0a017904",
			1938 => x"00101f11",
			1939 => x"00001f11",
			1940 => x"fe6f1f11",
			1941 => x"0c065054",
			1942 => x"0c05f630",
			1943 => x"0507f41c",
			1944 => x"0901f210",
			1945 => x"07063f08",
			1946 => x"0a020804",
			1947 => x"007a1f11",
			1948 => x"feca1f11",
			1949 => x"0b06ed04",
			1950 => x"01691f11",
			1951 => x"ffa71f11",
			1952 => x"0b06dc04",
			1953 => x"fdee1f11",
			1954 => x"01014104",
			1955 => x"00551f11",
			1956 => x"00001f11",
			1957 => x"0b070110",
			1958 => x"06017408",
			1959 => x"0e090704",
			1960 => x"00001f11",
			1961 => x"fe371f11",
			1962 => x"01014504",
			1963 => x"00001f11",
			1964 => x"ffa81f11",
			1965 => x"00001f11",
			1966 => x"0100e908",
			1967 => x"03094f04",
			1968 => x"02271f11",
			1969 => x"003b1f11",
			1970 => x"0601400c",
			1971 => x"09017d04",
			1972 => x"00ab1f11",
			1973 => x"09018304",
			1974 => x"febf1f11",
			1975 => x"00931f11",
			1976 => x"02092008",
			1977 => x"01011704",
			1978 => x"015d1f11",
			1979 => x"00001f11",
			1980 => x"0e093304",
			1981 => x"feff1f11",
			1982 => x"00a11f11",
			1983 => x"09019604",
			1984 => x"f9761f11",
			1985 => x"020a2d04",
			1986 => x"00aa1f11",
			1987 => x"feec1f11",
			1988 => x"0c05d810",
			1989 => x"0003460c",
			1990 => x"0b06bb04",
			1991 => x"00002015",
			1992 => x"08024e04",
			1993 => x"00002015",
			1994 => x"00a02015",
			1995 => x"fe672015",
			1996 => x"02093a30",
			1997 => x"01010f24",
			1998 => x"03096818",
			1999 => x"0002dd0c",
			2000 => x"0b06ed08",
			2001 => x"04091d04",
			2002 => x"00ef2015",
			2003 => x"00002015",
			2004 => x"ff512015",
			2005 => x"0a01e904",
			2006 => x"00002015",
			2007 => x"09017604",
			2008 => x"00002015",
			2009 => x"01852015",
			2010 => x"08025f08",
			2011 => x"0002ee04",
			2012 => x"ff552015",
			2013 => x"00002015",
			2014 => x"00d52015",
			2015 => x"0e08e104",
			2016 => x"febc2015",
			2017 => x"03094004",
			2018 => x"00002015",
			2019 => x"006a2015",
			2020 => x"0e09872c",
			2021 => x"0409db18",
			2022 => x"0a021710",
			2023 => x"07068308",
			2024 => x"0f096004",
			2025 => x"00002015",
			2026 => x"fed52015",
			2027 => x"0b071004",
			2028 => x"00002015",
			2029 => x"004f2015",
			2030 => x"0901d904",
			2031 => x"01182015",
			2032 => x"00002015",
			2033 => x"0309b00c",
			2034 => x"0c05da04",
			2035 => x"00002015",
			2036 => x"06017704",
			2037 => x"fe6e2015",
			2038 => x"00002015",
			2039 => x"06017404",
			2040 => x"00032015",
			2041 => x"00002015",
			2042 => x"040a3a04",
			2043 => x"01382015",
			2044 => x"0309ef04",
			2045 => x"feef2015",
			2046 => x"0b071e08",
			2047 => x"01014504",
			2048 => x"01322015",
			2049 => x"00002015",
			2050 => x"07072504",
			2051 => x"ff1a2015",
			2052 => x"00002015",
			2053 => x"09017a08",
			2054 => x"0600ef04",
			2055 => x"00002109",
			2056 => x"fe822109",
			2057 => x"0901dd48",
			2058 => x"00030c28",
			2059 => x"0002e618",
			2060 => x"0d084b08",
			2061 => x"0d083e04",
			2062 => x"01042109",
			2063 => x"00002109",
			2064 => x"0f092a08",
			2065 => x"08025a04",
			2066 => x"fe942109",
			2067 => x"00002109",
			2068 => x"02091904",
			2069 => x"00312109",
			2070 => x"ff382109",
			2071 => x"0208d004",
			2072 => x"ff9d2109",
			2073 => x"0f099508",
			2074 => x"07064004",
			2075 => x"00002109",
			2076 => x"01202109",
			2077 => x"00002109",
			2078 => x"0c066a18",
			2079 => x"040a2810",
			2080 => x"0b06dd08",
			2081 => x"0a021704",
			2082 => x"fe812109",
			2083 => x"ffe92109",
			2084 => x"0100ff04",
			2085 => x"ff7c2109",
			2086 => x"00de2109",
			2087 => x"0c064d04",
			2088 => x"fe972109",
			2089 => x"00002109",
			2090 => x"040b4204",
			2091 => x"00cb2109",
			2092 => x"00002109",
			2093 => x"00037814",
			2094 => x"06016f08",
			2095 => x"0901df04",
			2096 => x"00002109",
			2097 => x"ff4c2109",
			2098 => x"0e096204",
			2099 => x"00002109",
			2100 => x"0706b404",
			2101 => x"01462109",
			2102 => x"00002109",
			2103 => x"0e0a1b04",
			2104 => x"feca2109",
			2105 => x"06018d08",
			2106 => x"0a025704",
			2107 => x"00002109",
			2108 => x"ff982109",
			2109 => x"0f0ac308",
			2110 => x"0b072f04",
			2111 => x"00fe2109",
			2112 => x"00002109",
			2113 => x"ffef2109",
			2114 => x"00039a70",
			2115 => x"0706704c",
			2116 => x"07066e38",
			2117 => x"0507e418",
			2118 => x"0101260c",
			2119 => x"03097808",
			2120 => x"01010f04",
			2121 => x"007a21ed",
			2122 => x"febf21ed",
			2123 => x"018e21ed",
			2124 => x"0507ca04",
			2125 => x"fe1221ed",
			2126 => x"0c05f804",
			2127 => x"005d21ed",
			2128 => x"ff1421ed",
			2129 => x"0c05f610",
			2130 => x"0507ea08",
			2131 => x"0100ef04",
			2132 => x"000021ed",
			2133 => x"00e121ed",
			2134 => x"0d083f04",
			2135 => x"000021ed",
			2136 => x"fed621ed",
			2137 => x"0100ef08",
			2138 => x"05082104",
			2139 => x"005221ed",
			2140 => x"fef621ed",
			2141 => x"00037d04",
			2142 => x"019821ed",
			2143 => x"ff2121ed",
			2144 => x"06014104",
			2145 => x"000021ed",
			2146 => x"06016708",
			2147 => x"03096804",
			2148 => x"000021ed",
			2149 => x"fe4621ed",
			2150 => x"0901e804",
			2151 => x"000021ed",
			2152 => x"ffb221ed",
			2153 => x"0c065018",
			2154 => x"0d08b310",
			2155 => x"0002dd04",
			2156 => x"000021ed",
			2157 => x"0b070e08",
			2158 => x"0b06fe04",
			2159 => x"013121ed",
			2160 => x"000021ed",
			2161 => x"01a921ed",
			2162 => x"05089404",
			2163 => x"ff6121ed",
			2164 => x"000021ed",
			2165 => x"0901a104",
			2166 => x"fdef21ed",
			2167 => x"01014504",
			2168 => x"008321ed",
			2169 => x"ffc421ed",
			2170 => x"fe7421ed",
			2171 => x"0c05d508",
			2172 => x"07064104",
			2173 => x"fe7622e9",
			2174 => x"000022e9",
			2175 => x"06013e20",
			2176 => x"0d086d1c",
			2177 => x"0b06dc0c",
			2178 => x"0c05f204",
			2179 => x"000022e9",
			2180 => x"0d083e04",
			2181 => x"00fd22e9",
			2182 => x"000022e9",
			2183 => x"07065b08",
			2184 => x"0d083804",
			2185 => x"000022e9",
			2186 => x"ff2022e9",
			2187 => x"0100eb04",
			2188 => x"000022e9",
			2189 => x"007b22e9",
			2190 => x"018822e9",
			2191 => x"0507e428",
			2192 => x"01012614",
			2193 => x"0e094010",
			2194 => x"01010f08",
			2195 => x"0802b304",
			2196 => x"010222e9",
			2197 => x"ffa422e9",
			2198 => x"0c05f504",
			2199 => x"000022e9",
			2200 => x"fe7722e9",
			2201 => x"018122e9",
			2202 => x"0d08380c",
			2203 => x"07062a04",
			2204 => x"000022e9",
			2205 => x"0a023004",
			2206 => x"000022e9",
			2207 => x"fe3022e9",
			2208 => x"0a026d04",
			2209 => x"003822e9",
			2210 => x"000022e9",
			2211 => x"0507ea14",
			2212 => x"0101410c",
			2213 => x"0d085908",
			2214 => x"020a2d04",
			2215 => x"018322e9",
			2216 => x"000022e9",
			2217 => x"000022e9",
			2218 => x"07065504",
			2219 => x"000022e9",
			2220 => x"ff9422e9",
			2221 => x"0c064d10",
			2222 => x"07067008",
			2223 => x"07066c04",
			2224 => x"004922e9",
			2225 => x"ff2f22e9",
			2226 => x"0d08b304",
			2227 => x"012c22e9",
			2228 => x"ffc022e9",
			2229 => x"0b072004",
			2230 => x"fe5822e9",
			2231 => x"06017804",
			2232 => x"00d222e9",
			2233 => x"ff0322e9",
			2234 => x"0c05d408",
			2235 => x"07064204",
			2236 => x"fe7123d5",
			2237 => x"000023d5",
			2238 => x"0c065060",
			2239 => x"0c061334",
			2240 => x"0706581c",
			2241 => x"07064010",
			2242 => x"07062b08",
			2243 => x"00035304",
			2244 => x"00c323d5",
			2245 => x"000023d5",
			2246 => x"0a021d04",
			2247 => x"fe8e23d5",
			2248 => x"000023d5",
			2249 => x"08024e04",
			2250 => x"ff9a23d5",
			2251 => x"00037d04",
			2252 => x"014a23d5",
			2253 => x"fffb23d5",
			2254 => x"0f091508",
			2255 => x"0a01e404",
			2256 => x"000023d5",
			2257 => x"018e23d5",
			2258 => x"0c05db08",
			2259 => x"0d084c04",
			2260 => x"fdbf23d5",
			2261 => x"000023d5",
			2262 => x"06014204",
			2263 => x"fe9f23d5",
			2264 => x"ffc423d5",
			2265 => x"0d083f10",
			2266 => x"0c061a0c",
			2267 => x"00034b08",
			2268 => x"0100eb04",
			2269 => x"000023d5",
			2270 => x"00fa23d5",
			2271 => x"000023d5",
			2272 => x"febb23d5",
			2273 => x"0d088d10",
			2274 => x"06014108",
			2275 => x"06013a04",
			2276 => x"013623d5",
			2277 => x"ffd923d5",
			2278 => x"00039604",
			2279 => x"017923d5",
			2280 => x"000023d5",
			2281 => x"07066f04",
			2282 => x"ff0823d5",
			2283 => x"0d08b304",
			2284 => x"00f923d5",
			2285 => x"ffec23d5",
			2286 => x"0b072004",
			2287 => x"fc3e23d5",
			2288 => x"06017404",
			2289 => x"00a423d5",
			2290 => x"0706a104",
			2291 => x"000023d5",
			2292 => x"fed323d5",
			2293 => x"00039a80",
			2294 => x"0100f140",
			2295 => x"07066c24",
			2296 => x"07065a18",
			2297 => x"03092e10",
			2298 => x"0c05f208",
			2299 => x"07064304",
			2300 => x"fea024db",
			2301 => x"000024db",
			2302 => x"09017a04",
			2303 => x"004024db",
			2304 => x"029924db",
			2305 => x"0507e604",
			2306 => x"000024db",
			2307 => x"fe9224db",
			2308 => x"0002dd08",
			2309 => x"03092e04",
			2310 => x"000024db",
			2311 => x"ffbe24db",
			2312 => x"027124db",
			2313 => x"03094f0c",
			2314 => x"07067208",
			2315 => x"0208dd04",
			2316 => x"002424db",
			2317 => x"000024db",
			2318 => x"038624db",
			2319 => x"0002e604",
			2320 => x"fdaf24db",
			2321 => x"07066e04",
			2322 => x"fdd324db",
			2323 => x"02095704",
			2324 => x"014f24db",
			2325 => x"feed24db",
			2326 => x"07065b20",
			2327 => x"0c062e1c",
			2328 => x"0003530c",
			2329 => x"01013a08",
			2330 => x"0507ba04",
			2331 => x"ffb824db",
			2332 => x"013124db",
			2333 => x"fe4324db",
			2334 => x"06017c08",
			2335 => x"0c061004",
			2336 => x"fe1724db",
			2337 => x"000024db",
			2338 => x"0507e404",
			2339 => x"feb324db",
			2340 => x"013b24db",
			2341 => x"fe3524db",
			2342 => x"0d08da18",
			2343 => x"09018708",
			2344 => x"02093a04",
			2345 => x"00a824db",
			2346 => x"ffcd24db",
			2347 => x"0b06dc08",
			2348 => x"00035304",
			2349 => x"011824db",
			2350 => x"ffc124db",
			2351 => x"00039504",
			2352 => x"018624db",
			2353 => x"030e24db",
			2354 => x"07072504",
			2355 => x"fea224db",
			2356 => x"005024db",
			2357 => x"fe6924db",
			2358 => x"000024dd",
			2359 => x"000024e1",
			2360 => x"000024e5",
			2361 => x"0c060f04",
			2362 => x"000024f9",
			2363 => x"0c064d04",
			2364 => x"000824f9",
			2365 => x"000024f9",
			2366 => x"0c05d804",
			2367 => x"0000250d",
			2368 => x"00037804",
			2369 => x"0011250d",
			2370 => x"0000250d",
			2371 => x"00030c08",
			2372 => x"00022e04",
			2373 => x"00002521",
			2374 => x"00072521",
			2375 => x"00002521",
			2376 => x"0507e708",
			2377 => x"0506f104",
			2378 => x"0000253d",
			2379 => x"0015253d",
			2380 => x"05081f04",
			2381 => x"fff2253d",
			2382 => x"0000253d",
			2383 => x"040a2808",
			2384 => x"0207c504",
			2385 => x"00002559",
			2386 => x"000b2559",
			2387 => x"020a5004",
			2388 => x"fff42559",
			2389 => x"00002559",
			2390 => x"0e09870c",
			2391 => x"07065b08",
			2392 => x"0901b204",
			2393 => x"ffcb257d",
			2394 => x"0000257d",
			2395 => x"0000257d",
			2396 => x"020a2d04",
			2397 => x"0036257d",
			2398 => x"0000257d",
			2399 => x"0c06320c",
			2400 => x"0c05f404",
			2401 => x"000025a1",
			2402 => x"0c061304",
			2403 => x"ffef25a1",
			2404 => x"000025a1",
			2405 => x"0c064d04",
			2406 => x"000125a1",
			2407 => x"000025a1",
			2408 => x"0003240c",
			2409 => x"02090904",
			2410 => x"000025cd",
			2411 => x"0c05f304",
			2412 => x"000025cd",
			2413 => x"004625cd",
			2414 => x"0c063408",
			2415 => x"020a8c04",
			2416 => x"ffc725cd",
			2417 => x"000025cd",
			2418 => x"000025cd",
			2419 => x"04091d04",
			2420 => x"000025f1",
			2421 => x"0b07330c",
			2422 => x"0e0a1b08",
			2423 => x"030a3904",
			2424 => x"ffab25f1",
			2425 => x"000025f1",
			2426 => x"000025f1",
			2427 => x"000025f1",
			2428 => x"040a2810",
			2429 => x"0507ba04",
			2430 => x"00002615",
			2431 => x"05081208",
			2432 => x"0408c304",
			2433 => x"00002615",
			2434 => x"001f2615",
			2435 => x"00002615",
			2436 => x"00002615",
			2437 => x"0c063210",
			2438 => x"06013a04",
			2439 => x"00002641",
			2440 => x"06017708",
			2441 => x"0b06bc04",
			2442 => x"00002641",
			2443 => x"ffb82641",
			2444 => x"00002641",
			2445 => x"0c064d04",
			2446 => x"00022641",
			2447 => x"00002641",
			2448 => x"06013e08",
			2449 => x"0c05f204",
			2450 => x"0000266d",
			2451 => x"0043266d",
			2452 => x"0c06320c",
			2453 => x"04097204",
			2454 => x"0000266d",
			2455 => x"06016f04",
			2456 => x"ffd5266d",
			2457 => x"0000266d",
			2458 => x"0000266d",
			2459 => x"0209200c",
			2460 => x"00030c08",
			2461 => x"0207c504",
			2462 => x"000026a1",
			2463 => x"002a26a1",
			2464 => x"000026a1",
			2465 => x"02097b04",
			2466 => x"ffe326a1",
			2467 => x"00036308",
			2468 => x"00031a04",
			2469 => x"000026a1",
			2470 => x"001e26a1",
			2471 => x"000026a1",
			2472 => x"040a3a14",
			2473 => x"0a01ec04",
			2474 => x"000026d5",
			2475 => x"0101240c",
			2476 => x"09017a04",
			2477 => x"000026d5",
			2478 => x"0e08cb04",
			2479 => x"000026d5",
			2480 => x"004b26d5",
			2481 => x"000026d5",
			2482 => x"09020e04",
			2483 => x"ffd326d5",
			2484 => x"000026d5",
			2485 => x"00037014",
			2486 => x"0c05d804",
			2487 => x"00002701",
			2488 => x"0d087f0c",
			2489 => x"0d080b04",
			2490 => x"00002701",
			2491 => x"0a01e904",
			2492 => x"00002701",
			2493 => x"00402701",
			2494 => x"00002701",
			2495 => x"00002701",
			2496 => x"05082114",
			2497 => x"0c05f204",
			2498 => x"0000272d",
			2499 => x"0003850c",
			2500 => x"0c062e08",
			2501 => x"0d087404",
			2502 => x"0069272d",
			2503 => x"0000272d",
			2504 => x"0000272d",
			2505 => x"0000272d",
			2506 => x"0000272d",
			2507 => x"0100f30c",
			2508 => x"02092004",
			2509 => x"00002769",
			2510 => x"0d086604",
			2511 => x"00002769",
			2512 => x"ffaf2769",
			2513 => x"0c05f304",
			2514 => x"00002769",
			2515 => x"020a930c",
			2516 => x"01015208",
			2517 => x"0d083f04",
			2518 => x"00002769",
			2519 => x"005b2769",
			2520 => x"00002769",
			2521 => x"00002769",
			2522 => x"0507ba08",
			2523 => x"0e098704",
			2524 => x"ffc327ad",
			2525 => x"000027ad",
			2526 => x"0507e710",
			2527 => x"020a2d0c",
			2528 => x"0e08cb04",
			2529 => x"000027ad",
			2530 => x"0208db04",
			2531 => x"000027ad",
			2532 => x"005727ad",
			2533 => x"000027ad",
			2534 => x"07067004",
			2535 => x"ffed27ad",
			2536 => x"0706cb04",
			2537 => x"001a27ad",
			2538 => x"000027ad",
			2539 => x"00030c10",
			2540 => x"0901a90c",
			2541 => x"04095908",
			2542 => x"0b063c04",
			2543 => x"00002801",
			2544 => x"002d2801",
			2545 => x"00002801",
			2546 => x"00002801",
			2547 => x"0901dd0c",
			2548 => x"0b073308",
			2549 => x"0b06bc04",
			2550 => x"00002801",
			2551 => x"ffaa2801",
			2552 => x"00002801",
			2553 => x"00037d0c",
			2554 => x"0b06d204",
			2555 => x"00002801",
			2556 => x"0b073304",
			2557 => x"00402801",
			2558 => x"00002801",
			2559 => x"00002801",
			2560 => x"040a3a18",
			2561 => x"09018304",
			2562 => x"0000283d",
			2563 => x"01013610",
			2564 => x"07063d04",
			2565 => x"0000283d",
			2566 => x"0b06a504",
			2567 => x"0000283d",
			2568 => x"0a023e04",
			2569 => x"007e283d",
			2570 => x"0000283d",
			2571 => x"0000283d",
			2572 => x"0901f804",
			2573 => x"fff5283d",
			2574 => x"0000283d",
			2575 => x"0e093308",
			2576 => x"0d075504",
			2577 => x"00002879",
			2578 => x"fffb2879",
			2579 => x"0d089a14",
			2580 => x"09018304",
			2581 => x"00002879",
			2582 => x"0e0a860c",
			2583 => x"0d080e04",
			2584 => x"00002879",
			2585 => x"09021b04",
			2586 => x"002e2879",
			2587 => x"00002879",
			2588 => x"00002879",
			2589 => x"00002879",
			2590 => x"0100f108",
			2591 => x"0a017904",
			2592 => x"000028b5",
			2593 => x"ffea28b5",
			2594 => x"0f0ab614",
			2595 => x"01015010",
			2596 => x"09018704",
			2597 => x"000028b5",
			2598 => x"0a01f204",
			2599 => x"000028b5",
			2600 => x"0a027404",
			2601 => x"002928b5",
			2602 => x"000028b5",
			2603 => x"000028b5",
			2604 => x"000028b5",
			2605 => x"0601771c",
			2606 => x"0409c710",
			2607 => x"0c061208",
			2608 => x"0c05d704",
			2609 => x"00002911",
			2610 => x"004b2911",
			2611 => x"0c063204",
			2612 => x"ffc62911",
			2613 => x"00002911",
			2614 => x"0b073308",
			2615 => x"0a020004",
			2616 => x"00002911",
			2617 => x"ff6f2911",
			2618 => x"00002911",
			2619 => x"00037d10",
			2620 => x"05084d0c",
			2621 => x"0c05dc04",
			2622 => x"00002911",
			2623 => x"0e097704",
			2624 => x"00002911",
			2625 => x"00932911",
			2626 => x"00002911",
			2627 => x"00002911",
			2628 => x"040a3a18",
			2629 => x"0309ef14",
			2630 => x"0c05d904",
			2631 => x"00002945",
			2632 => x"0c062e0c",
			2633 => x"07066c08",
			2634 => x"00032404",
			2635 => x"006d2945",
			2636 => x"00002945",
			2637 => x"00002945",
			2638 => x"00002945",
			2639 => x"00002945",
			2640 => x"00002945",
			2641 => x"0003851c",
			2642 => x"0e093308",
			2643 => x"04091d04",
			2644 => x"00002981",
			2645 => x"fff42981",
			2646 => x"0d083104",
			2647 => x"00002981",
			2648 => x"0508300c",
			2649 => x"0c05dc04",
			2650 => x"00002981",
			2651 => x"09018304",
			2652 => x"00002981",
			2653 => x"00942981",
			2654 => x"00002981",
			2655 => x"00002981",
			2656 => x"0f092a0c",
			2657 => x"08025a08",
			2658 => x"07064404",
			2659 => x"000029dd",
			2660 => x"ff9629dd",
			2661 => x"000029dd",
			2662 => x"0c061410",
			2663 => x"0a021d08",
			2664 => x"06013e04",
			2665 => x"000029dd",
			2666 => x"ffe329dd",
			2667 => x"0a025704",
			2668 => x"001229dd",
			2669 => x"000029dd",
			2670 => x"0c064d10",
			2671 => x"0d08b30c",
			2672 => x"0e08fd04",
			2673 => x"000029dd",
			2674 => x"0a027704",
			2675 => x"008f29dd",
			2676 => x"000029dd",
			2677 => x"000029dd",
			2678 => x"000029dd",
			2679 => x"040a0124",
			2680 => x"0c061110",
			2681 => x"0c05f604",
			2682 => x"00002a49",
			2683 => x"0a01df04",
			2684 => x"00002a49",
			2685 => x"0b06a504",
			2686 => x"00002a49",
			2687 => x"00682a49",
			2688 => x"0b071010",
			2689 => x"00031a0c",
			2690 => x"0c063208",
			2691 => x"0208c904",
			2692 => x"00002a49",
			2693 => x"ff9e2a49",
			2694 => x"00002a49",
			2695 => x"00002a49",
			2696 => x"002a2a49",
			2697 => x"0209e80c",
			2698 => x"00033504",
			2699 => x"00002a49",
			2700 => x"0b06cc04",
			2701 => x"00002a49",
			2702 => x"ffa22a49",
			2703 => x"020a2d04",
			2704 => x"00042a49",
			2705 => x"00002a49",
			2706 => x"040a3a20",
			2707 => x"08025a08",
			2708 => x"0100e904",
			2709 => x"00002a9d",
			2710 => x"ffff2a9d",
			2711 => x"07064004",
			2712 => x"00002a9d",
			2713 => x"06014104",
			2714 => x"00002a9d",
			2715 => x"0c06500c",
			2716 => x"06015f08",
			2717 => x"00032404",
			2718 => x"00892a9d",
			2719 => x"00002a9d",
			2720 => x"00002a9d",
			2721 => x"00002a9d",
			2722 => x"06019408",
			2723 => x"0c066a04",
			2724 => x"ffa62a9d",
			2725 => x"00002a9d",
			2726 => x"00002a9d",
			2727 => x"040a3a1c",
			2728 => x"0a01ec04",
			2729 => x"00002ae9",
			2730 => x"0c05f604",
			2731 => x"00002ae9",
			2732 => x"0c065010",
			2733 => x"0e08cb04",
			2734 => x"00002ae9",
			2735 => x"09017d04",
			2736 => x"00002ae9",
			2737 => x"0d080104",
			2738 => x"00002ae9",
			2739 => x"007a2ae9",
			2740 => x"00002ae9",
			2741 => x"06018c08",
			2742 => x"0c06c504",
			2743 => x"ffbc2ae9",
			2744 => x"00002ae9",
			2745 => x"00002ae9",
			2746 => x"0c06321c",
			2747 => x"0901fc18",
			2748 => x"0b06bc04",
			2749 => x"00002b2d",
			2750 => x"0100e804",
			2751 => x"00002b2d",
			2752 => x"0f08f004",
			2753 => x"00002b2d",
			2754 => x"0802b308",
			2755 => x"07062b04",
			2756 => x"00002b2d",
			2757 => x"ffa42b2d",
			2758 => x"00002b2d",
			2759 => x"00002b2d",
			2760 => x"0c064d04",
			2761 => x"00012b2d",
			2762 => x"00002b2d",
			2763 => x"0901f824",
			2764 => x"0b06cc14",
			2765 => x"0b063c04",
			2766 => x"00002b99",
			2767 => x"0101340c",
			2768 => x"0f0a0308",
			2769 => x"0e078e04",
			2770 => x"00002b99",
			2771 => x"001d2b99",
			2772 => x"00002b99",
			2773 => x"00002b99",
			2774 => x"0b06ec0c",
			2775 => x"0f08f004",
			2776 => x"00002b99",
			2777 => x"0e09a204",
			2778 => x"ffa72b99",
			2779 => x"00002b99",
			2780 => x"00002b99",
			2781 => x"0b074410",
			2782 => x"0507d904",
			2783 => x"00002b99",
			2784 => x"0f0ac308",
			2785 => x"020aa804",
			2786 => x"00512b99",
			2787 => x"00002b99",
			2788 => x"00002b99",
			2789 => x"00002b99",
			2790 => x"05082124",
			2791 => x"0507c70c",
			2792 => x"0002e604",
			2793 => x"00002bfd",
			2794 => x"06016f04",
			2795 => x"ffb42bfd",
			2796 => x"00002bfd",
			2797 => x"0c062e14",
			2798 => x"06014104",
			2799 => x"00002bfd",
			2800 => x"020a2d0c",
			2801 => x"08025304",
			2802 => x"00002bfd",
			2803 => x"0a025704",
			2804 => x"00a62bfd",
			2805 => x"00002bfd",
			2806 => x"00002bfd",
			2807 => x"00002bfd",
			2808 => x"0b07330c",
			2809 => x"0e0a3908",
			2810 => x"0309ef04",
			2811 => x"00002bfd",
			2812 => x"ffa62bfd",
			2813 => x"00002bfd",
			2814 => x"00002bfd",
			2815 => x"0d084b1c",
			2816 => x"00035314",
			2817 => x"09017a04",
			2818 => x"00002c79",
			2819 => x"07063f04",
			2820 => x"00002c79",
			2821 => x"0b06f008",
			2822 => x"0d080104",
			2823 => x"00002c79",
			2824 => x"00d62c79",
			2825 => x"00002c79",
			2826 => x"0d084a04",
			2827 => x"ffeb2c79",
			2828 => x"00002c79",
			2829 => x"06014910",
			2830 => x"0a01ec04",
			2831 => x"00002c79",
			2832 => x"0b06ec04",
			2833 => x"00002c79",
			2834 => x"02095704",
			2835 => x"004c2c79",
			2836 => x"00002c79",
			2837 => x"0a022808",
			2838 => x"07068304",
			2839 => x"ff792c79",
			2840 => x"00002c79",
			2841 => x"00037808",
			2842 => x"020a4604",
			2843 => x"00262c79",
			2844 => x"00002c79",
			2845 => x"00002c79",
			2846 => x"04091d04",
			2847 => x"00002cb5",
			2848 => x"0b06ef18",
			2849 => x"0e0a1b14",
			2850 => x"0b06cc04",
			2851 => x"00002cb5",
			2852 => x"07062c04",
			2853 => x"00002cb5",
			2854 => x"05081308",
			2855 => x"07067204",
			2856 => x"ff9a2cb5",
			2857 => x"00002cb5",
			2858 => x"00002cb5",
			2859 => x"00002cb5",
			2860 => x"00002cb5",
			2861 => x"09017d04",
			2862 => x"00002cf1",
			2863 => x"00039a18",
			2864 => x"0c05f604",
			2865 => x"00002cf1",
			2866 => x"05088610",
			2867 => x"0a01e404",
			2868 => x"00002cf1",
			2869 => x"01015508",
			2870 => x"0b06a504",
			2871 => x"00002cf1",
			2872 => x"004a2cf1",
			2873 => x"00002cf1",
			2874 => x"00002cf1",
			2875 => x"00002cf1",
			2876 => x"0003891c",
			2877 => x"0c05bc04",
			2878 => x"00002d2d",
			2879 => x"09017a04",
			2880 => x"00002d2d",
			2881 => x"07064604",
			2882 => x"00002d2d",
			2883 => x"02090004",
			2884 => x"00002d2d",
			2885 => x"01015408",
			2886 => x"030a8a04",
			2887 => x"00582d2d",
			2888 => x"00002d2d",
			2889 => x"00002d2d",
			2890 => x"00002d2d",
			2891 => x"04091d04",
			2892 => x"00002d79",
			2893 => x"05081f1c",
			2894 => x"0e098714",
			2895 => x"0b071010",
			2896 => x"0b06bc04",
			2897 => x"00002d79",
			2898 => x"0c05de04",
			2899 => x"00002d79",
			2900 => x"0309b004",
			2901 => x"ff8c2d79",
			2902 => x"00002d79",
			2903 => x"00002d79",
			2904 => x"0a025704",
			2905 => x"001c2d79",
			2906 => x"00002d79",
			2907 => x"0309a304",
			2908 => x"00022d79",
			2909 => x"00002d79",
			2910 => x"0003241c",
			2911 => x"01010f10",
			2912 => x"07061304",
			2913 => x"00002e05",
			2914 => x"0f096808",
			2915 => x"03098704",
			2916 => x"007a2e05",
			2917 => x"00002e05",
			2918 => x"00002e05",
			2919 => x"0a021708",
			2920 => x"07062b04",
			2921 => x"00002e05",
			2922 => x"ff9f2e05",
			2923 => x"00002e05",
			2924 => x"0901dd10",
			2925 => x"0706f60c",
			2926 => x"0409ed08",
			2927 => x"0409c704",
			2928 => x"fffe2e05",
			2929 => x"00002e05",
			2930 => x"ff432e05",
			2931 => x"00002e05",
			2932 => x"0d083f10",
			2933 => x"0507bc04",
			2934 => x"00002e05",
			2935 => x"0e097704",
			2936 => x"00002e05",
			2937 => x"0507e404",
			2938 => x"ffd92e05",
			2939 => x"00002e05",
			2940 => x"0d08b308",
			2941 => x"0e0aa404",
			2942 => x"003d2e05",
			2943 => x"00002e05",
			2944 => x"00002e05",
			2945 => x"0c061328",
			2946 => x"04091d08",
			2947 => x"0100aa04",
			2948 => x"00002e81",
			2949 => x"00072e81",
			2950 => x"0901c310",
			2951 => x"0706700c",
			2952 => x"06013e04",
			2953 => x"00002e81",
			2954 => x"0b06cc04",
			2955 => x"00002e81",
			2956 => x"ff952e81",
			2957 => x"00002e81",
			2958 => x"01013d0c",
			2959 => x"07065808",
			2960 => x"07061704",
			2961 => x"00002e81",
			2962 => x"00262e81",
			2963 => x"00002e81",
			2964 => x"00002e81",
			2965 => x"0002dd04",
			2966 => x"00002e81",
			2967 => x"06014e08",
			2968 => x"0c061604",
			2969 => x"00002e81",
			2970 => x"00942e81",
			2971 => x"01010204",
			2972 => x"ffcf2e81",
			2973 => x"01015204",
			2974 => x"00492e81",
			2975 => x"00002e81",
			2976 => x"0e09872c",
			2977 => x"00030c1c",
			2978 => x"03097814",
			2979 => x"09017a04",
			2980 => x"00002efd",
			2981 => x"06014a0c",
			2982 => x"0100e704",
			2983 => x"00002efd",
			2984 => x"0002dd04",
			2985 => x"00002efd",
			2986 => x"00912efd",
			2987 => x"00002efd",
			2988 => x"08026404",
			2989 => x"fffe2efd",
			2990 => x"00002efd",
			2991 => x"0507ac04",
			2992 => x"00002efd",
			2993 => x"0d088d08",
			2994 => x"0b06bc04",
			2995 => x"00002efd",
			2996 => x"ffad2efd",
			2997 => x"00002efd",
			2998 => x"00037d10",
			2999 => x"040ac90c",
			3000 => x"08029e04",
			3001 => x"00002efd",
			3002 => x"01014b04",
			3003 => x"00762efd",
			3004 => x"00002efd",
			3005 => x"00002efd",
			3006 => x"00002efd",
			3007 => x"0c06132c",
			3008 => x"04095910",
			3009 => x"0c05d704",
			3010 => x"00002f81",
			3011 => x"07066c08",
			3012 => x"07061304",
			3013 => x"00002f81",
			3014 => x"002a2f81",
			3015 => x"00002f81",
			3016 => x"0901dd0c",
			3017 => x"0b06bc04",
			3018 => x"00002f81",
			3019 => x"0e092404",
			3020 => x"00002f81",
			3021 => x"ff7d2f81",
			3022 => x"0101360c",
			3023 => x"0e096204",
			3024 => x"00002f81",
			3025 => x"0a025904",
			3026 => x"00392f81",
			3027 => x"00002f81",
			3028 => x"00002f81",
			3029 => x"0e093304",
			3030 => x"00002f81",
			3031 => x"01015010",
			3032 => x"0100ed04",
			3033 => x"00002f81",
			3034 => x"00039d08",
			3035 => x"0d090f04",
			3036 => x"00b22f81",
			3037 => x"00002f81",
			3038 => x"00002f81",
			3039 => x"00002f81",
			3040 => x"040a0134",
			3041 => x"0d084b18",
			3042 => x"07063f04",
			3043 => x"00003015",
			3044 => x"09017a04",
			3045 => x"00003015",
			3046 => x"0b06f00c",
			3047 => x"0a01e404",
			3048 => x"00003015",
			3049 => x"0d080b04",
			3050 => x"00003015",
			3051 => x"00ae3015",
			3052 => x"00003015",
			3053 => x"0b06f00c",
			3054 => x"0309b008",
			3055 => x"0f08f004",
			3056 => x"00003015",
			3057 => x"ffcc3015",
			3058 => x"00003015",
			3059 => x"03098708",
			3060 => x"0f092a04",
			3061 => x"00003015",
			3062 => x"00773015",
			3063 => x"02097b04",
			3064 => x"ffff3015",
			3065 => x"00003015",
			3066 => x"0309d80c",
			3067 => x"0e09a208",
			3068 => x"00033504",
			3069 => x"00003015",
			3070 => x"ff5d3015",
			3071 => x"00003015",
			3072 => x"00037008",
			3073 => x"00033e04",
			3074 => x"00003015",
			3075 => x"005b3015",
			3076 => x"00003015",
			3077 => x"00032420",
			3078 => x"0d08180c",
			3079 => x"01010f08",
			3080 => x"0100aa04",
			3081 => x"000030a9",
			3082 => x"000830a9",
			3083 => x"ffd930a9",
			3084 => x"05081210",
			3085 => x"0f08f904",
			3086 => x"000030a9",
			3087 => x"09017a04",
			3088 => x"000030a9",
			3089 => x"0e095104",
			3090 => x"00c430a9",
			3091 => x"000030a9",
			3092 => x"000030a9",
			3093 => x"0101260c",
			3094 => x"0b074408",
			3095 => x"0409b304",
			3096 => x"000030a9",
			3097 => x"ff3430a9",
			3098 => x"000030a9",
			3099 => x"0507e40c",
			3100 => x"01013604",
			3101 => x"000030a9",
			3102 => x"07065b04",
			3103 => x"ff7e30a9",
			3104 => x"000030a9",
			3105 => x"0d08b310",
			3106 => x"0101590c",
			3107 => x"0b06dc04",
			3108 => x"000030a9",
			3109 => x"00039a04",
			3110 => x"00a530a9",
			3111 => x"000030a9",
			3112 => x"000030a9",
			3113 => x"000030a9",
			3114 => x"00036334",
			3115 => x"0901dd28",
			3116 => x"0209781c",
			3117 => x"08027914",
			3118 => x"0100ff0c",
			3119 => x"09018308",
			3120 => x"07065804",
			3121 => x"fff9311d",
			3122 => x"0000311d",
			3123 => x"008a311d",
			3124 => x"07065b04",
			3125 => x"ff52311d",
			3126 => x"0000311d",
			3127 => x"0d082204",
			3128 => x"0000311d",
			3129 => x"00e9311d",
			3130 => x"0b073308",
			3131 => x"0901ce04",
			3132 => x"ff33311d",
			3133 => x"0000311d",
			3134 => x"0012311d",
			3135 => x"02099d04",
			3136 => x"0000311d",
			3137 => x"03099604",
			3138 => x"0000311d",
			3139 => x"00cc311d",
			3140 => x"0e0a3904",
			3141 => x"ff23311d",
			3142 => x"0000311d",
			3143 => x"0e098734",
			3144 => x"00030c1c",
			3145 => x"03097814",
			3146 => x"09017a04",
			3147 => x"000031a1",
			3148 => x"06014a0c",
			3149 => x"0100e704",
			3150 => x"000031a1",
			3151 => x"0002dd04",
			3152 => x"000031a1",
			3153 => x"009e31a1",
			3154 => x"000031a1",
			3155 => x"08026404",
			3156 => x"fff831a1",
			3157 => x"000031a1",
			3158 => x"0507ac04",
			3159 => x"000031a1",
			3160 => x"07062b04",
			3161 => x"000031a1",
			3162 => x"0b07200c",
			3163 => x"0b06bc04",
			3164 => x"000031a1",
			3165 => x"07068304",
			3166 => x"ff9831a1",
			3167 => x"000031a1",
			3168 => x"000031a1",
			3169 => x"00037d0c",
			3170 => x"01011904",
			3171 => x"000031a1",
			3172 => x"01014b04",
			3173 => x"007231a1",
			3174 => x"000031a1",
			3175 => x"000031a1",
			3176 => x"040a9530",
			3177 => x"09017a10",
			3178 => x"0706720c",
			3179 => x"0a017908",
			3180 => x"0c057f04",
			3181 => x"fe743245",
			3182 => x"05d63245",
			3183 => x"fe623245",
			3184 => x"00743245",
			3185 => x"0d080a08",
			3186 => x"08028704",
			3187 => x"01253245",
			3188 => x"fe6d3245",
			3189 => x"030a4910",
			3190 => x"0100e804",
			3191 => x"ff9f3245",
			3192 => x"0a025f08",
			3193 => x"0a01ec04",
			3194 => x"01b23245",
			3195 => x"02553245",
			3196 => x"fee83245",
			3197 => x"040a8804",
			3198 => x"fef63245",
			3199 => x"01433245",
			3200 => x"040af718",
			3201 => x"07065504",
			3202 => x"fe5d3245",
			3203 => x"0d08b310",
			3204 => x"05081208",
			3205 => x"0d085b04",
			3206 => x"fea93245",
			3207 => x"01d33245",
			3208 => x"0f0a7c04",
			3209 => x"03533245",
			3210 => x"05a13245",
			3211 => x"fe633245",
			3212 => x"040b2208",
			3213 => x"040b1c04",
			3214 => x"fe753245",
			3215 => x"ff713245",
			3216 => x"fe603245",
			3217 => x"00038938",
			3218 => x"0901760c",
			3219 => x"0600ef08",
			3220 => x"02069d04",
			3221 => x"fe9c32c9",
			3222 => x"01bf32c9",
			3223 => x"fe6832c9",
			3224 => x"0d08b324",
			3225 => x"0507ba0c",
			3226 => x"01010b08",
			3227 => x"0c05d904",
			3228 => x"fff832c9",
			3229 => x"01af32c9",
			3230 => x"fe4132c9",
			3231 => x"06018c10",
			3232 => x"00035308",
			3233 => x"0100ed04",
			3234 => x"007c32c9",
			3235 => x"019732c9",
			3236 => x"0309d804",
			3237 => x"fd9432c9",
			3238 => x"019f32c9",
			3239 => x"020a5004",
			3240 => x"025032c9",
			3241 => x"039c32c9",
			3242 => x"020a1804",
			3243 => x"006732c9",
			3244 => x"fe6d32c9",
			3245 => x"00039508",
			3246 => x"06019404",
			3247 => x"fe6f32c9",
			3248 => x"016932c9",
			3249 => x"fe6432c9",
			3250 => x"0003893c",
			3251 => x"0100e710",
			3252 => x"0b06fe0c",
			3253 => x"0600ef08",
			3254 => x"00022e04",
			3255 => x"fe8e3355",
			3256 => x"01d13355",
			3257 => x"fe663355",
			3258 => x"00003355",
			3259 => x"0d08b324",
			3260 => x"0507ba0c",
			3261 => x"01010b08",
			3262 => x"0c05d904",
			3263 => x"00003355",
			3264 => x"01c33355",
			3265 => x"fe3e3355",
			3266 => x"06018c10",
			3267 => x"0a01e408",
			3268 => x"0308f704",
			3269 => x"014e3355",
			3270 => x"fe5c3355",
			3271 => x"00035304",
			3272 => x"01b73355",
			3273 => x"00ca3355",
			3274 => x"05082e04",
			3275 => x"043a3355",
			3276 => x"029d3355",
			3277 => x"020a1804",
			3278 => x"00663355",
			3279 => x"fe633355",
			3280 => x"00039508",
			3281 => x"06019404",
			3282 => x"fe6a3355",
			3283 => x"01a73355",
			3284 => x"fe633355",
			3285 => x"0f092a10",
			3286 => x"0a017904",
			3287 => x"000033f9",
			3288 => x"09018308",
			3289 => x"0100ef04",
			3290 => x"ff8d33f9",
			3291 => x"000033f9",
			3292 => x"000033f9",
			3293 => x"0209b724",
			3294 => x"0a021714",
			3295 => x"0b06ec08",
			3296 => x"0507e704",
			3297 => x"000033f9",
			3298 => x"ff4c33f9",
			3299 => x"09017d04",
			3300 => x"000033f9",
			3301 => x"0100eb04",
			3302 => x"000033f9",
			3303 => x"007733f9",
			3304 => x"03094f04",
			3305 => x"000033f9",
			3306 => x"0d080e04",
			3307 => x"000033f9",
			3308 => x"0a023c04",
			3309 => x"00e433f9",
			3310 => x"000033f9",
			3311 => x"0e09a204",
			3312 => x"ff9a33f9",
			3313 => x"0d08b314",
			3314 => x"00037d08",
			3315 => x"06017304",
			3316 => x"000033f9",
			3317 => x"007033f9",
			3318 => x"09020e04",
			3319 => x"ffdb33f9",
			3320 => x"030a3904",
			3321 => x"000033f9",
			3322 => x"003f33f9",
			3323 => x"0b075f04",
			3324 => x"fff533f9",
			3325 => x"000033f9",
			3326 => x"00037d3c",
			3327 => x"09017a10",
			3328 => x"0508130c",
			3329 => x"0600ef08",
			3330 => x"09010a04",
			3331 => x"fe81349d",
			3332 => x"0269349d",
			3333 => x"fe64349d",
			3334 => x"fff4349d",
			3335 => x"0d07fd08",
			3336 => x"0901b204",
			3337 => x"00ed349d",
			3338 => x"fe73349d",
			3339 => x"0d08b31c",
			3340 => x"0a01e90c",
			3341 => x"03092204",
			3342 => x"0237349d",
			3343 => x"0507ea04",
			3344 => x"0000349d",
			3345 => x"fe36349d",
			3346 => x"0c05d908",
			3347 => x"00034b04",
			3348 => x"01b0349d",
			3349 => x"fe21349d",
			3350 => x"030a1204",
			3351 => x"01d8349d",
			3352 => x"02cd349d",
			3353 => x"00035b04",
			3354 => x"002e349d",
			3355 => x"fe6e349d",
			3356 => x"00039614",
			3357 => x"0802eb0c",
			3358 => x"00038108",
			3359 => x"0802dd04",
			3360 => x"fe9d349d",
			3361 => x"02fa349d",
			3362 => x"fe65349d",
			3363 => x"06019404",
			3364 => x"000f349d",
			3365 => x"033a349d",
			3366 => x"fe61349d",
			3367 => x"040abb34",
			3368 => x"0100e70c",
			3369 => x"0600ef08",
			3370 => x"0e060f04",
			3371 => x"feae3539",
			3372 => x"02733539",
			3373 => x"fe6e3539",
			3374 => x"0d080e0c",
			3375 => x"04091d04",
			3376 => x"01bb3539",
			3377 => x"0507c704",
			3378 => x"fe4d3539",
			3379 => x"00343539",
			3380 => x"01014b18",
			3381 => x"0a01e408",
			3382 => x"0208a604",
			3383 => x"009f3539",
			3384 => x"fe793539",
			3385 => x"02092808",
			3386 => x"05082104",
			3387 => x"01c83539",
			3388 => x"007a3539",
			3389 => x"08026404",
			3390 => x"ff3f3539",
			3391 => x"013c3539",
			3392 => x"fe9b3539",
			3393 => x"01014304",
			3394 => x"fe653539",
			3395 => x"030aa114",
			3396 => x"0d086d04",
			3397 => x"fed93539",
			3398 => x"07067208",
			3399 => x"040b2404",
			3400 => x"03173539",
			3401 => x"00003539",
			3402 => x"06019d04",
			3403 => x"fee93539",
			3404 => x"00f33539",
			3405 => x"fe6b3539",
			3406 => x"00032428",
			3407 => x"0d08180c",
			3408 => x"01010f08",
			3409 => x"0100aa04",
			3410 => x"000035fd",
			3411 => x"000735fd",
			3412 => x"ffdb35fd",
			3413 => x"06014d14",
			3414 => x"0e09240c",
			3415 => x"0d086d08",
			3416 => x"0d083f04",
			3417 => x"000035fd",
			3418 => x"fff635fd",
			3419 => x"009235fd",
			3420 => x"0d087204",
			3421 => x"ffc335fd",
			3422 => x"000035fd",
			3423 => x"0100fa04",
			3424 => x"000035fd",
			3425 => x"00d535fd",
			3426 => x"06016b0c",
			3427 => x"0c063208",
			3428 => x"0409b304",
			3429 => x"000035fd",
			3430 => x"ff2935fd",
			3431 => x"000035fd",
			3432 => x"07065810",
			3433 => x"0b06bd04",
			3434 => x"000035fd",
			3435 => x"0a026208",
			3436 => x"03097804",
			3437 => x"000035fd",
			3438 => x"009035fd",
			3439 => x"000035fd",
			3440 => x"030a3910",
			3441 => x"0a023604",
			3442 => x"000035fd",
			3443 => x"0e0a3908",
			3444 => x"06017404",
			3445 => x"000035fd",
			3446 => x"ffa635fd",
			3447 => x"000035fd",
			3448 => x"040b220c",
			3449 => x"0d08b308",
			3450 => x"05080f04",
			3451 => x"000035fd",
			3452 => x"006e35fd",
			3453 => x"000035fd",
			3454 => x"000035fd",
			3455 => x"0c05f61c",
			3456 => x"0e098708",
			3457 => x"00032404",
			3458 => x"00003699",
			3459 => x"fef43699",
			3460 => x"07065810",
			3461 => x"0f0a5a0c",
			3462 => x"07062c04",
			3463 => x"00003699",
			3464 => x"00038c04",
			3465 => x"005c3699",
			3466 => x"00003699",
			3467 => x"00003699",
			3468 => x"00003699",
			3469 => x"00038530",
			3470 => x"0e093318",
			3471 => x"0d086d10",
			3472 => x"07064204",
			3473 => x"00003699",
			3474 => x"0b06bd04",
			3475 => x"00003699",
			3476 => x"07066e04",
			3477 => x"ff823699",
			3478 => x"00003699",
			3479 => x"02092804",
			3480 => x"00ce3699",
			3481 => x"00003699",
			3482 => x"0100f304",
			3483 => x"00003699",
			3484 => x"0d083808",
			3485 => x"01013604",
			3486 => x"00423699",
			3487 => x"ffb63699",
			3488 => x"05088608",
			3489 => x"01014b04",
			3490 => x"01043699",
			3491 => x"00003699",
			3492 => x"00003699",
			3493 => x"ffd83699",
			3494 => x"00038940",
			3495 => x"030a122c",
			3496 => x"00035324",
			3497 => x"06016f1c",
			3498 => x"0f096010",
			3499 => x"0002e608",
			3500 => x"0507f504",
			3501 => x"00633725",
			3502 => x"ff403725",
			3503 => x"0d082204",
			3504 => x"ff893725",
			3505 => x"00f83725",
			3506 => x"0b073308",
			3507 => x"01010604",
			3508 => x"fee93725",
			3509 => x"ffe73725",
			3510 => x"00be3725",
			3511 => x"03097804",
			3512 => x"00003725",
			3513 => x"01743725",
			3514 => x"0309ef04",
			3515 => x"fe8a3725",
			3516 => x"00003725",
			3517 => x"020a2d04",
			3518 => x"01573725",
			3519 => x"0802e008",
			3520 => x"040ac204",
			3521 => x"00003725",
			3522 => x"ff863725",
			3523 => x"01015504",
			3524 => x"00de3725",
			3525 => x"00003725",
			3526 => x"01014d04",
			3527 => x"fe863725",
			3528 => x"00003725",
			3529 => x"0003242c",
			3530 => x"0d08180c",
			3531 => x"01010f08",
			3532 => x"0100aa04",
			3533 => x"000037f1",
			3534 => x"000737f1",
			3535 => x"ffdd37f1",
			3536 => x"06014d18",
			3537 => x"0d086d0c",
			3538 => x"0208e204",
			3539 => x"000037f1",
			3540 => x"0d083f04",
			3541 => x"000037f1",
			3542 => x"ffb437f1",
			3543 => x"0a01f708",
			3544 => x"0100ef04",
			3545 => x"00ae37f1",
			3546 => x"000037f1",
			3547 => x"000037f1",
			3548 => x"02099504",
			3549 => x"00cd37f1",
			3550 => x"000037f1",
			3551 => x"06016b0c",
			3552 => x"0c063208",
			3553 => x"0507ac04",
			3554 => x"000037f1",
			3555 => x"ff2537f1",
			3556 => x"000037f1",
			3557 => x"07065810",
			3558 => x"0b06bd04",
			3559 => x"000037f1",
			3560 => x"0a026208",
			3561 => x"03097804",
			3562 => x"000037f1",
			3563 => x"008937f1",
			3564 => x"000037f1",
			3565 => x"07066d10",
			3566 => x"0901e604",
			3567 => x"000037f1",
			3568 => x"0c063208",
			3569 => x"030a8104",
			3570 => x"ffa237f1",
			3571 => x"000037f1",
			3572 => x"000037f1",
			3573 => x"0d08b30c",
			3574 => x"0901d904",
			3575 => x"000037f1",
			3576 => x"0c05fa04",
			3577 => x"000037f1",
			3578 => x"006637f1",
			3579 => x"000037f1",
			3580 => x"05080138",
			3581 => x"02099d24",
			3582 => x"00032418",
			3583 => x"0a021010",
			3584 => x"0b06cc04",
			3585 => x"000038b5",
			3586 => x"0507f608",
			3587 => x"0b06ff04",
			3588 => x"ffa038b5",
			3589 => x"000038b5",
			3590 => x"000038b5",
			3591 => x"0d081804",
			3592 => x"000038b5",
			3593 => x"009c38b5",
			3594 => x"0c05fa08",
			3595 => x"07065b04",
			3596 => x"fee138b5",
			3597 => x"000038b5",
			3598 => x"000038b5",
			3599 => x"040a3a04",
			3600 => x"005d38b5",
			3601 => x"040ab20c",
			3602 => x"07066d08",
			3603 => x"0c05d904",
			3604 => x"000038b5",
			3605 => x"ff8a38b5",
			3606 => x"000038b5",
			3607 => x"000038b5",
			3608 => x"00038524",
			3609 => x"0a01e904",
			3610 => x"000038b5",
			3611 => x"0d087f0c",
			3612 => x"09017d04",
			3613 => x"000038b5",
			3614 => x"0c05f504",
			3615 => x"000038b5",
			3616 => x"00f438b5",
			3617 => x"0c063208",
			3618 => x"09018704",
			3619 => x"ffed38b5",
			3620 => x"000038b5",
			3621 => x"020a3a08",
			3622 => x"09020a04",
			3623 => x"005738b5",
			3624 => x"000038b5",
			3625 => x"000038b5",
			3626 => x"0c061504",
			3627 => x"000038b5",
			3628 => x"ffe338b5",
			3629 => x"0901760c",
			3630 => x"0a017908",
			3631 => x"0406a304",
			3632 => x"00003961",
			3633 => x"00173961",
			3634 => x"fe6e3961",
			3635 => x"04091d10",
			3636 => x"03092e0c",
			3637 => x"0100e804",
			3638 => x"00003961",
			3639 => x"09017a04",
			3640 => x"00003961",
			3641 => x"01b93961",
			3642 => x"ffc53961",
			3643 => x"0e0a1b24",
			3644 => x"0c063218",
			3645 => x"0d08820c",
			3646 => x"030a1208",
			3647 => x"0901f404",
			3648 => x"fff63961",
			3649 => x"fedd3961",
			3650 => x"01763961",
			3651 => x"0309ef08",
			3652 => x"02096c04",
			3653 => x"ff6d3961",
			3654 => x"00733961",
			3655 => x"fe7c3961",
			3656 => x"040aa908",
			3657 => x"0100ed04",
			3658 => x"ffc43961",
			3659 => x"01703961",
			3660 => x"ff703961",
			3661 => x"0d08b310",
			3662 => x"0a027408",
			3663 => x"0b06dd04",
			3664 => x"00003961",
			3665 => x"01b33961",
			3666 => x"0d089a04",
			3667 => x"ffce3961",
			3668 => x"00003961",
			3669 => x"0b074404",
			3670 => x"00003961",
			3671 => x"fedc3961",
			3672 => x"00036348",
			3673 => x"06016230",
			3674 => x"01010f24",
			3675 => x"0f096814",
			3676 => x"09018310",
			3677 => x"0b070108",
			3678 => x"03092e04",
			3679 => x"000039fd",
			3680 => x"ffcf39fd",
			3681 => x"02090004",
			3682 => x"000039fd",
			3683 => x"006039fd",
			3684 => x"00b739fd",
			3685 => x"0b07330c",
			3686 => x"01010608",
			3687 => x"0c05f404",
			3688 => x"000039fd",
			3689 => x"ff5c39fd",
			3690 => x"000039fd",
			3691 => x"000039fd",
			3692 => x"0a021708",
			3693 => x"07062b04",
			3694 => x"000039fd",
			3695 => x"ff3639fd",
			3696 => x"000039fd",
			3697 => x"0901b804",
			3698 => x"000039fd",
			3699 => x"0c05f30c",
			3700 => x"07064408",
			3701 => x"07062604",
			3702 => x"000039fd",
			3703 => x"000b39fd",
			3704 => x"000039fd",
			3705 => x"03094f04",
			3706 => x"000039fd",
			3707 => x"011d39fd",
			3708 => x"0e0a3904",
			3709 => x"ff1639fd",
			3710 => x"000039fd",
			3711 => x"00037848",
			3712 => x"0100e920",
			3713 => x"0100e710",
			3714 => x"0a017908",
			3715 => x"0705a204",
			3716 => x"fe6e3ad9",
			3717 => x"0d7a3ad9",
			3718 => x"07067004",
			3719 => x"fe603ad9",
			3720 => x"ff6b3ad9",
			3721 => x"0d083808",
			3722 => x"0b06d204",
			3723 => x"ff083ad9",
			3724 => x"07993ad9",
			3725 => x"0b06ef04",
			3726 => x"fe713ad9",
			3727 => x"00003ad9",
			3728 => x"0d080a08",
			3729 => x"0208e204",
			3730 => x"01953ad9",
			3731 => x"fe683ad9",
			3732 => x"0d08da18",
			3733 => x"0a01e90c",
			3734 => x"03091a04",
			3735 => x"02fc3ad9",
			3736 => x"0c061504",
			3737 => x"fe503ad9",
			3738 => x"002c3ad9",
			3739 => x"0c05d504",
			3740 => x"ffe23ad9",
			3741 => x"0507bb04",
			3742 => x"01953ad9",
			3743 => x"03043ad9",
			3744 => x"00036804",
			3745 => x"00203ad9",
			3746 => x"fe873ad9",
			3747 => x"00039a24",
			3748 => x"0802eb18",
			3749 => x"0802e810",
			3750 => x"00037d0c",
			3751 => x"05084d08",
			3752 => x"0c05db04",
			3753 => x"fea33ad9",
			3754 => x"02283ad9",
			3755 => x"fe6a3ad9",
			3756 => x"fe5f3ad9",
			3757 => x"0c063004",
			3758 => x"05ec3ad9",
			3759 => x"fe833ad9",
			3760 => x"0706a108",
			3761 => x"0b070e04",
			3762 => x"01dc3ad9",
			3763 => x"06253ad9",
			3764 => x"fe9a3ad9",
			3765 => x"fe5d3ad9",
			3766 => x"00032438",
			3767 => x"0d084a14",
			3768 => x"0c05d704",
			3769 => x"00003b9d",
			3770 => x"0101210c",
			3771 => x"0b06ee08",
			3772 => x"07060204",
			3773 => x"00003b9d",
			3774 => x"00e83b9d",
			3775 => x"00003b9d",
			3776 => x"00003b9d",
			3777 => x"0c061618",
			3778 => x"0b06ec0c",
			3779 => x"0507ea04",
			3780 => x"00003b9d",
			3781 => x"0f090d04",
			3782 => x"00003b9d",
			3783 => x"ff1e3b9d",
			3784 => x"0002f608",
			3785 => x"0208fe04",
			3786 => x"00003b9d",
			3787 => x"ffcd3b9d",
			3788 => x"00263b9d",
			3789 => x"02097808",
			3790 => x"02090004",
			3791 => x"00003b9d",
			3792 => x"00cf3b9d",
			3793 => x"00003b9d",
			3794 => x"0e094004",
			3795 => x"fec63b9d",
			3796 => x"0f09b104",
			3797 => x"00be3b9d",
			3798 => x"0706410c",
			3799 => x"020a2d08",
			3800 => x"0d080e04",
			3801 => x"00003b9d",
			3802 => x"00433b9d",
			3803 => x"00003b9d",
			3804 => x"0209e808",
			3805 => x"0c05fa04",
			3806 => x"ff043b9d",
			3807 => x"00003b9d",
			3808 => x"020a2d08",
			3809 => x"0802de04",
			3810 => x"00863b9d",
			3811 => x"00003b9d",
			3812 => x"07066e04",
			3813 => x"ff783b9d",
			3814 => x"00003b9d",
			3815 => x"07063f10",
			3816 => x"04093104",
			3817 => x"00003c71",
			3818 => x"03098708",
			3819 => x"0b06cf04",
			3820 => x"fead3c71",
			3821 => x"00003c71",
			3822 => x"00003c71",
			3823 => x"0b06dd24",
			3824 => x"0b06cc10",
			3825 => x"0101340c",
			3826 => x"03094f04",
			3827 => x"00003c71",
			3828 => x"040a5b04",
			3829 => x"00d23c71",
			3830 => x"00003c71",
			3831 => x"00003c71",
			3832 => x"07064404",
			3833 => x"00003c71",
			3834 => x"0f08f004",
			3835 => x"00003c71",
			3836 => x"0c05de04",
			3837 => x"00003c71",
			3838 => x"07067004",
			3839 => x"ff193c71",
			3840 => x"00003c71",
			3841 => x"040a3a20",
			3842 => x"0706460c",
			3843 => x"0901b808",
			3844 => x"03092e04",
			3845 => x"00003c71",
			3846 => x"ffb43c71",
			3847 => x"00003c71",
			3848 => x"0100f310",
			3849 => x"0a01f708",
			3850 => x"03098704",
			3851 => x"00793c71",
			3852 => x"00003c71",
			3853 => x"07068504",
			3854 => x"ff8e3c71",
			3855 => x"00003c71",
			3856 => x"012e3c71",
			3857 => x"0e0a1b0c",
			3858 => x"0508a308",
			3859 => x"030a5c04",
			3860 => x"ff703c71",
			3861 => x"00003c71",
			3862 => x"00003c71",
			3863 => x"040af708",
			3864 => x"0d08b304",
			3865 => x"00983c71",
			3866 => x"00003c71",
			3867 => x"00003c71",
			3868 => x"01011340",
			3869 => x"0409ed38",
			3870 => x"0d083e10",
			3871 => x"0100e804",
			3872 => x"00003d4d",
			3873 => x"0d081704",
			3874 => x"00003d4d",
			3875 => x"0a01df04",
			3876 => x"00003d4d",
			3877 => x"009a3d4d",
			3878 => x"02090910",
			3879 => x"0d084b04",
			3880 => x"00003d4d",
			3881 => x"0a01f208",
			3882 => x"0208db04",
			3883 => x"00003d4d",
			3884 => x"ff5a3d4d",
			3885 => x"00003d4d",
			3886 => x"07065b0c",
			3887 => x"0e093308",
			3888 => x"0b06f004",
			3889 => x"ffc63d4d",
			3890 => x"00003d4d",
			3891 => x"00003d4d",
			3892 => x"0100e904",
			3893 => x"00003d4d",
			3894 => x"02097804",
			3895 => x"00713d4d",
			3896 => x"00003d4d",
			3897 => x"0c065004",
			3898 => x"ff463d4d",
			3899 => x"00003d4d",
			3900 => x"0a025714",
			3901 => x"0507ca04",
			3902 => x"00003d4d",
			3903 => x"0c05db04",
			3904 => x"00003d4d",
			3905 => x"040abb08",
			3906 => x"01014b04",
			3907 => x"01033d4d",
			3908 => x"00003d4d",
			3909 => x"00003d4d",
			3910 => x"0e0a1b08",
			3911 => x"07064404",
			3912 => x"00003d4d",
			3913 => x"ffbc3d4d",
			3914 => x"040af710",
			3915 => x"0c05f804",
			3916 => x"00003d4d",
			3917 => x"030a2804",
			3918 => x"00003d4d",
			3919 => x"0706a104",
			3920 => x"00753d4d",
			3921 => x"00003d4d",
			3922 => x"00003d4d",
			3923 => x"0c05dc14",
			3924 => x"00034610",
			3925 => x"02093a08",
			3926 => x"0c05d704",
			3927 => x"ff7f3e31",
			3928 => x"00003e31",
			3929 => x"0b06bb04",
			3930 => x"00003e31",
			3931 => x"00c93e31",
			3932 => x"fe8f3e31",
			3933 => x"0c061340",
			3934 => x"0d085924",
			3935 => x"01013d1c",
			3936 => x"0d082210",
			3937 => x"0507ad08",
			3938 => x"00033e04",
			3939 => x"00f23e31",
			3940 => x"00003e31",
			3941 => x"0507ba04",
			3942 => x"fee73e31",
			3943 => x"00003e31",
			3944 => x"06013d04",
			3945 => x"00003e31",
			3946 => x"0b06ee04",
			3947 => x"01443e31",
			3948 => x"00003e31",
			3949 => x"0b06e004",
			3950 => x"ff363e31",
			3951 => x"00003e31",
			3952 => x"0c060f0c",
			3953 => x"01011508",
			3954 => x"0e090704",
			3955 => x"00003e31",
			3956 => x"fecb3e31",
			3957 => x"00003e31",
			3958 => x"0c06120c",
			3959 => x"05082108",
			3960 => x"05080104",
			3961 => x"00003e31",
			3962 => x"00b43e31",
			3963 => x"00003e31",
			3964 => x"ff8f3e31",
			3965 => x"0209000c",
			3966 => x"0100ef08",
			3967 => x"04090804",
			3968 => x"00003e31",
			3969 => x"ffc33e31",
			3970 => x"00003e31",
			3971 => x"01014b10",
			3972 => x"0100e704",
			3973 => x"00003e31",
			3974 => x"040af708",
			3975 => x"0507c704",
			3976 => x"00003e31",
			3977 => x"01083e31",
			3978 => x"00003e31",
			3979 => x"00003e31",
			3980 => x"0507c71c",
			3981 => x"0002e60c",
			3982 => x"0c05f204",
			3983 => x"00003f35",
			3984 => x"0b06bd04",
			3985 => x"00c63f35",
			3986 => x"00003f35",
			3987 => x"0e098708",
			3988 => x"04090804",
			3989 => x"00003f35",
			3990 => x"fe6e3f35",
			3991 => x"06018804",
			3992 => x"00813f35",
			3993 => x"00003f35",
			3994 => x"02093a30",
			3995 => x"0002e624",
			3996 => x"0100e910",
			3997 => x"07065804",
			3998 => x"00003f35",
			3999 => x"03094f08",
			4000 => x"0e08d604",
			4001 => x"00003f35",
			4002 => x"01863f35",
			4003 => x"00003f35",
			4004 => x"02090c10",
			4005 => x"0208e208",
			4006 => x"09018004",
			4007 => x"00003f35",
			4008 => x"00223f35",
			4009 => x"07065904",
			4010 => x"00003f35",
			4011 => x"feea3f35",
			4012 => x"00003f35",
			4013 => x"0100eb04",
			4014 => x"00003f35",
			4015 => x"03098704",
			4016 => x"014d3f35",
			4017 => x"00003f35",
			4018 => x"0901c31c",
			4019 => x"0b07100c",
			4020 => x"0507ea04",
			4021 => x"00513f35",
			4022 => x"0c063004",
			4023 => x"feb13f35",
			4024 => x"00003f35",
			4025 => x"0a020804",
			4026 => x"00dc3f35",
			4027 => x"0a021004",
			4028 => x"ffb63f35",
			4029 => x"0209ce04",
			4030 => x"00403f35",
			4031 => x"00003f35",
			4032 => x"040a3a08",
			4033 => x"0507cc04",
			4034 => x"00003f35",
			4035 => x"01433f35",
			4036 => x"0309ef04",
			4037 => x"fed43f35",
			4038 => x"0c062e08",
			4039 => x"01014504",
			4040 => x"01233f35",
			4041 => x"00003f35",
			4042 => x"07072504",
			4043 => x"ff593f35",
			4044 => x"00003f35",
			4045 => x"00039650",
			4046 => x"0e0a1b44",
			4047 => x"00033524",
			4048 => x"0a021d18",
			4049 => x"00032410",
			4050 => x"08025a08",
			4051 => x"04091d04",
			4052 => x"009e3fd9",
			4053 => x"ff5b3fd9",
			4054 => x"0d087f04",
			4055 => x"00f23fd9",
			4056 => x"ffcf3fd9",
			4057 => x"07062b04",
			4058 => x"00003fd9",
			4059 => x"fe7d3fd9",
			4060 => x"06016204",
			4061 => x"00003fd9",
			4062 => x"0b06bb04",
			4063 => x"00003fd9",
			4064 => x"017d3fd9",
			4065 => x"0e09a210",
			4066 => x"040a0108",
			4067 => x"0d081704",
			4068 => x"00003fd9",
			4069 => x"01073fd9",
			4070 => x"07065c04",
			4071 => x"fe343fd9",
			4072 => x"00003fd9",
			4073 => x"0003700c",
			4074 => x"00034608",
			4075 => x"0b06ef04",
			4076 => x"00003fd9",
			4077 => x"fed03fd9",
			4078 => x"01523fd9",
			4079 => x"fe983fd9",
			4080 => x"0d08b304",
			4081 => x"01573fd9",
			4082 => x"0802ed04",
			4083 => x"ffeb3fd9",
			4084 => x"00003fd9",
			4085 => x"fe7c3fd9",
			4086 => x"0b06dd44",
			4087 => x"0e094024",
			4088 => x"00030c1c",
			4089 => x"08025a14",
			4090 => x"04091d0c",
			4091 => x"0307f404",
			4092 => x"000040fd",
			4093 => x"03091a04",
			4094 => x"003b40fd",
			4095 => x"000040fd",
			4096 => x"0b06cd04",
			4097 => x"fef340fd",
			4098 => x"000040fd",
			4099 => x"0100ed04",
			4100 => x"000040fd",
			4101 => x"00c240fd",
			4102 => x"04097204",
			4103 => x"000040fd",
			4104 => x"fe7540fd",
			4105 => x"0b06cc08",
			4106 => x"00035b04",
			4107 => x"011540fd",
			4108 => x"000040fd",
			4109 => x"0409db04",
			4110 => x"000040fd",
			4111 => x"0901d904",
			4112 => x"fef040fd",
			4113 => x"0901f408",
			4114 => x"0802c304",
			4115 => x"007040fd",
			4116 => x"000040fd",
			4117 => x"0d084a04",
			4118 => x"ff3c40fd",
			4119 => x"000040fd",
			4120 => x"0507f418",
			4121 => x"01013d10",
			4122 => x"0b06fc0c",
			4123 => x"06013d04",
			4124 => x"000040fd",
			4125 => x"00038504",
			4126 => x"014840fd",
			4127 => x"000040fd",
			4128 => x"000040fd",
			4129 => x"0507e604",
			4130 => x"ffbd40fd",
			4131 => x"000040fd",
			4132 => x"0c060f10",
			4133 => x"0e092404",
			4134 => x"000040fd",
			4135 => x"030a2808",
			4136 => x"0c05fa04",
			4137 => x"feb340fd",
			4138 => x"000040fd",
			4139 => x"000040fd",
			4140 => x"0002e610",
			4141 => x"03094f08",
			4142 => x"0f090d04",
			4143 => x"000040fd",
			4144 => x"00a040fd",
			4145 => x"05081f04",
			4146 => x"ff0e40fd",
			4147 => x"000040fd",
			4148 => x"0d08b310",
			4149 => x"0c064d08",
			4150 => x"00039d04",
			4151 => x"00ee40fd",
			4152 => x"000040fd",
			4153 => x"06015204",
			4154 => x"000040fd",
			4155 => x"ffc440fd",
			4156 => x"0901c804",
			4157 => x"000040fd",
			4158 => x"ff3040fd",
			4159 => x"0c05d818",
			4160 => x"00034614",
			4161 => x"07062c08",
			4162 => x"02096004",
			4163 => x"ff544201",
			4164 => x"00004201",
			4165 => x"0a01df04",
			4166 => x"00004201",
			4167 => x"07064004",
			4168 => x"00004201",
			4169 => x"00604201",
			4170 => x"fe844201",
			4171 => x"0507e72c",
			4172 => x"01013d20",
			4173 => x"0d080e0c",
			4174 => x"0002e604",
			4175 => x"00004201",
			4176 => x"07065a04",
			4177 => x"ff0d4201",
			4178 => x"00004201",
			4179 => x"00035b08",
			4180 => x"06013d04",
			4181 => x"00004201",
			4182 => x"01364201",
			4183 => x"0901fa04",
			4184 => x"fff64201",
			4185 => x"030a2804",
			4186 => x"00174201",
			4187 => x"00004201",
			4188 => x"0c05f404",
			4189 => x"00004201",
			4190 => x"0c061504",
			4191 => x"ff204201",
			4192 => x"00004201",
			4193 => x"0507f610",
			4194 => x"0d08660c",
			4195 => x"0309d808",
			4196 => x"0f095604",
			4197 => x"00004201",
			4198 => x"feee4201",
			4199 => x"00004201",
			4200 => x"008a4201",
			4201 => x"0100f118",
			4202 => x"03094f08",
			4203 => x"08025304",
			4204 => x"00004201",
			4205 => x"00f74201",
			4206 => x"07066c08",
			4207 => x"07065a04",
			4208 => x"00004201",
			4209 => x"00c04201",
			4210 => x"0002e604",
			4211 => x"fef54201",
			4212 => x"00004201",
			4213 => x"0d08b30c",
			4214 => x"01015708",
			4215 => x"040b2204",
			4216 => x"01484201",
			4217 => x"00004201",
			4218 => x"00004201",
			4219 => x"0706b704",
			4220 => x"ff274201",
			4221 => x"020a2d04",
			4222 => x"00dd4201",
			4223 => x"ffeb4201",
			4224 => x"00039654",
			4225 => x"0e0a1b48",
			4226 => x"00033524",
			4227 => x"08025a10",
			4228 => x"0601420c",
			4229 => x"07068308",
			4230 => x"06013b04",
			4231 => x"ffcb42ad",
			4232 => x"00c142ad",
			4233 => x"feb942ad",
			4234 => x"fe9142ad",
			4235 => x"02092808",
			4236 => x"0d07fd04",
			4237 => x"000042ad",
			4238 => x"016042ad",
			4239 => x"06016b08",
			4240 => x"00032404",
			4241 => x"003042ad",
			4242 => x"ff1242ad",
			4243 => x"016542ad",
			4244 => x"0e09a214",
			4245 => x"0507ab08",
			4246 => x"0b06bd04",
			4247 => x"ffad42ad",
			4248 => x"009f42ad",
			4249 => x"05080108",
			4250 => x"07062e04",
			4251 => x"000042ad",
			4252 => x"fe5942ad",
			4253 => x"000042ad",
			4254 => x"0003700c",
			4255 => x"00034608",
			4256 => x"0b06ef04",
			4257 => x"000042ad",
			4258 => x"feb942ad",
			4259 => x"015c42ad",
			4260 => x"fe8c42ad",
			4261 => x"0d088204",
			4262 => x"017942ad",
			4263 => x"0802e904",
			4264 => x"ffca42ad",
			4265 => x"000042ad",
			4266 => x"fe7942ad",
			4267 => x"0c05d810",
			4268 => x"0003460c",
			4269 => x"0e093308",
			4270 => x"07064304",
			4271 => x"ff2f43b1",
			4272 => x"000043b1",
			4273 => x"006a43b1",
			4274 => x"fe7943b1",
			4275 => x"0507e730",
			4276 => x"01013d24",
			4277 => x"0507ca18",
			4278 => x"03097810",
			4279 => x"0002e608",
			4280 => x"0c05f204",
			4281 => x"000043b1",
			4282 => x"007c43b1",
			4283 => x"0c05de04",
			4284 => x"000043b1",
			4285 => x"ff4f43b1",
			4286 => x"01013004",
			4287 => x"010443b1",
			4288 => x"000043b1",
			4289 => x"06013d04",
			4290 => x"000043b1",
			4291 => x"00037d04",
			4292 => x"015343b1",
			4293 => x"000043b1",
			4294 => x"0c05f404",
			4295 => x"000043b1",
			4296 => x"0c061504",
			4297 => x"ff1043b1",
			4298 => x"000043b1",
			4299 => x"0507f61c",
			4300 => x"0f095610",
			4301 => x"06014108",
			4302 => x"03092204",
			4303 => x"000043b1",
			4304 => x"fff443b1",
			4305 => x"0e08e104",
			4306 => x"000043b1",
			4307 => x"00fe43b1",
			4308 => x"0309d808",
			4309 => x"0b06e004",
			4310 => x"febb43b1",
			4311 => x"000043b1",
			4312 => x"000043b1",
			4313 => x"0100f118",
			4314 => x"03094f08",
			4315 => x"08025304",
			4316 => x"000043b1",
			4317 => x"012a43b1",
			4318 => x"07066c08",
			4319 => x"07065a04",
			4320 => x"000043b1",
			4321 => x"00d843b1",
			4322 => x"0c063204",
			4323 => x"ff1243b1",
			4324 => x"000043b1",
			4325 => x"0101560c",
			4326 => x"040b2208",
			4327 => x"05088604",
			4328 => x"00fa43b1",
			4329 => x"000043b1",
			4330 => x"000043b1",
			4331 => x"ffcd43b1",
			4332 => x"0c05d508",
			4333 => x"07064304",
			4334 => x"fe7f448d",
			4335 => x"0000448d",
			4336 => x"00032438",
			4337 => x"08025a18",
			4338 => x"04091d0c",
			4339 => x"03092208",
			4340 => x"09017a04",
			4341 => x"0000448d",
			4342 => x"0138448d",
			4343 => x"0000448d",
			4344 => x"02090004",
			4345 => x"fe92448d",
			4346 => x"0c061404",
			4347 => x"ff64448d",
			4348 => x"00c3448d",
			4349 => x"0d087f10",
			4350 => x"0d081808",
			4351 => x"01011304",
			4352 => x"0000448d",
			4353 => x"ff3c448d",
			4354 => x"0309b004",
			4355 => x"015e448d",
			4356 => x"0000448d",
			4357 => x"07068508",
			4358 => x"0100f304",
			4359 => x"fec6448d",
			4360 => x"0042448d",
			4361 => x"06014f04",
			4362 => x"011c448d",
			4363 => x"0000448d",
			4364 => x"0a021d04",
			4365 => x"fe81448d",
			4366 => x"0003350c",
			4367 => x"06016304",
			4368 => x"0000448d",
			4369 => x"02094904",
			4370 => x"0000448d",
			4371 => x"0165448d",
			4372 => x"0e09a210",
			4373 => x"040a0108",
			4374 => x"0d081704",
			4375 => x"0000448d",
			4376 => x"00fc448d",
			4377 => x"07065c04",
			4378 => x"fe42448d",
			4379 => x"0000448d",
			4380 => x"00038508",
			4381 => x"030a1204",
			4382 => x"0000448d",
			4383 => x"014a448d",
			4384 => x"030a4904",
			4385 => x"fec9448d",
			4386 => x"0000448d",
			4387 => x"09017614",
			4388 => x"0600ef10",
			4389 => x"0600ee04",
			4390 => x"000045a1",
			4391 => x"00022e04",
			4392 => x"000045a1",
			4393 => x"00045404",
			4394 => x"002d45a1",
			4395 => x"000045a1",
			4396 => x"fe6d45a1",
			4397 => x"0c05f640",
			4398 => x"00034b20",
			4399 => x"07063f10",
			4400 => x"07062b08",
			4401 => x"0d07fd04",
			4402 => x"000045a1",
			4403 => x"009545a1",
			4404 => x"0b06bc04",
			4405 => x"000045a1",
			4406 => x"fe0845a1",
			4407 => x"0d085b0c",
			4408 => x"09018004",
			4409 => x"000045a1",
			4410 => x"0c05f504",
			4411 => x"018945a1",
			4412 => x"000845a1",
			4413 => x"ff0445a1",
			4414 => x"0b06e010",
			4415 => x"07066d0c",
			4416 => x"0901f804",
			4417 => x"fdc945a1",
			4418 => x"0901fa04",
			4419 => x"000045a1",
			4420 => x"ff4545a1",
			4421 => x"000045a1",
			4422 => x"0c05f304",
			4423 => x"000045a1",
			4424 => x"0c05f508",
			4425 => x"020ad104",
			4426 => x"005345a1",
			4427 => x"000045a1",
			4428 => x"000045a1",
			4429 => x"0d08b328",
			4430 => x"030a011c",
			4431 => x"00035b10",
			4432 => x"06016808",
			4433 => x"02099504",
			4434 => x"003845a1",
			4435 => x"fe7945a1",
			4436 => x"03096804",
			4437 => x"000045a1",
			4438 => x"016645a1",
			4439 => x"0c061508",
			4440 => x"0c05f704",
			4441 => x"000045a1",
			4442 => x"fe6d45a1",
			4443 => x"000045a1",
			4444 => x"01015508",
			4445 => x"00039d04",
			4446 => x"01b945a1",
			4447 => x"fff545a1",
			4448 => x"ffbd45a1",
			4449 => x"0901c30c",
			4450 => x"01010b04",
			4451 => x"ff5e45a1",
			4452 => x"0d090104",
			4453 => x"00bf45a1",
			4454 => x"000045a1",
			4455 => x"fe9445a1",
			4456 => x"0d080e14",
			4457 => x"0002dd0c",
			4458 => x"07061304",
			4459 => x"000046b5",
			4460 => x"0507c704",
			4461 => x"002746b5",
			4462 => x"000046b5",
			4463 => x"07064604",
			4464 => x"fe7646b5",
			4465 => x"000046b5",
			4466 => x"0901dd50",
			4467 => x"0409b330",
			4468 => x"0d083e14",
			4469 => x"0d08180c",
			4470 => x"0c05f608",
			4471 => x"07064404",
			4472 => x"ff5946b5",
			4473 => x"000046b5",
			4474 => x"000046b5",
			4475 => x"0a01e404",
			4476 => x"000046b5",
			4477 => x"016b46b5",
			4478 => x"0002e60c",
			4479 => x"05081f08",
			4480 => x"0208dd04",
			4481 => x"000046b5",
			4482 => x"fe9b46b5",
			4483 => x"ffd646b5",
			4484 => x"00030c08",
			4485 => x"0c05f304",
			4486 => x"000046b5",
			4487 => x"010546b5",
			4488 => x"01010b04",
			4489 => x"febd46b5",
			4490 => x"001a46b5",
			4491 => x"0c066a14",
			4492 => x"040a2810",
			4493 => x"0a021d08",
			4494 => x"07068304",
			4495 => x"fe7446b5",
			4496 => x"000046b5",
			4497 => x"0507d804",
			4498 => x"ffb146b5",
			4499 => x"011546b5",
			4500 => x"fe7c46b5",
			4501 => x"01010604",
			4502 => x"000046b5",
			4503 => x"06019904",
			4504 => x"00e146b5",
			4505 => x"000046b5",
			4506 => x"0003780c",
			4507 => x"0a023304",
			4508 => x"fff346b5",
			4509 => x"05086a04",
			4510 => x"015746b5",
			4511 => x"000046b5",
			4512 => x"0e0a1b04",
			4513 => x"feb146b5",
			4514 => x"06018d08",
			4515 => x"0a025704",
			4516 => x"000046b5",
			4517 => x"ff7e46b5",
			4518 => x"0f0aad08",
			4519 => x"01015504",
			4520 => x"011546b5",
			4521 => x"000046b5",
			4522 => x"0f0ac304",
			4523 => x"000046b5",
			4524 => x"ffc346b5",
			4525 => x"00039a78",
			4526 => x"0100f138",
			4527 => x"07066c20",
			4528 => x"07065a14",
			4529 => x"04091d0c",
			4530 => x"06013d08",
			4531 => x"0600ef04",
			4532 => x"009247a9",
			4533 => x"ff2847a9",
			4534 => x"023c47a9",
			4535 => x"09018304",
			4536 => x"fe6e47a9",
			4537 => x"003547a9",
			4538 => x"0002dd08",
			4539 => x"03092e04",
			4540 => x"000047a9",
			4541 => x"ffd347a9",
			4542 => x"023847a9",
			4543 => x"03094f08",
			4544 => x"08025304",
			4545 => x"000047a9",
			4546 => x"02a247a9",
			4547 => x"0002e604",
			4548 => x"fdeb47a9",
			4549 => x"07066e04",
			4550 => x"fe0a47a9",
			4551 => x"08026904",
			4552 => x"014547a9",
			4553 => x"ff0847a9",
			4554 => x"07065b24",
			4555 => x"040a3a14",
			4556 => x"07065a10",
			4557 => x"0507ba08",
			4558 => x"01012604",
			4559 => x"000e47a9",
			4560 => x"fe5847a9",
			4561 => x"0d084b04",
			4562 => x"014847a9",
			4563 => x"002947a9",
			4564 => x"feae47a9",
			4565 => x"0309d804",
			4566 => x"fdf147a9",
			4567 => x"020a2d04",
			4568 => x"016147a9",
			4569 => x"0802de04",
			4570 => x"fe6647a9",
			4571 => x"000947a9",
			4572 => x"05086a10",
			4573 => x"0100f304",
			4574 => x"000047a9",
			4575 => x"0507ca04",
			4576 => x"000047a9",
			4577 => x"0f0a9204",
			4578 => x"015c47a9",
			4579 => x"027a47a9",
			4580 => x"07072508",
			4581 => x"05088604",
			4582 => x"000047a9",
			4583 => x"feae47a9",
			4584 => x"004147a9",
			4585 => x"fe6a47a9",
			4586 => x"07063f14",
			4587 => x"0409870c",
			4588 => x"01011108",
			4589 => x"0100aa04",
			4590 => x"000048d5",
			4591 => x"004248d5",
			4592 => x"000048d5",
			4593 => x"03097804",
			4594 => x"fe7148d5",
			4595 => x"000048d5",
			4596 => x"0706582c",
			4597 => x"06016c20",
			4598 => x"040a011c",
			4599 => x"0a01f210",
			4600 => x"06013e08",
			4601 => x"0c061004",
			4602 => x"000048d5",
			4603 => x"001d48d5",
			4604 => x"0f08f004",
			4605 => x"000048d5",
			4606 => x"ff9348d5",
			4607 => x"09018b04",
			4608 => x"000048d5",
			4609 => x"03094f04",
			4610 => x"000048d5",
			4611 => x"00ed48d5",
			4612 => x"ff5f48d5",
			4613 => x"00037d08",
			4614 => x"03099604",
			4615 => x"000048d5",
			4616 => x"014b48d5",
			4617 => x"fff548d5",
			4618 => x"06014a24",
			4619 => x"03097818",
			4620 => x"02090010",
			4621 => x"04093108",
			4622 => x"0208c204",
			4623 => x"000048d5",
			4624 => x"005948d5",
			4625 => x"0c061004",
			4626 => x"000048d5",
			4627 => x"ffb248d5",
			4628 => x"05080104",
			4629 => x"000048d5",
			4630 => x"010648d5",
			4631 => x"0002ee04",
			4632 => x"ff4648d5",
			4633 => x"0c061304",
			4634 => x"000048d5",
			4635 => x"007048d5",
			4636 => x"0507f61c",
			4637 => x"07065b0c",
			4638 => x"0d082204",
			4639 => x"000048d5",
			4640 => x"0d085b04",
			4641 => x"fee648d5",
			4642 => x"000048d5",
			4643 => x"07066f08",
			4644 => x"06018904",
			4645 => x"005448d5",
			4646 => x"000048d5",
			4647 => x"0d084b04",
			4648 => x"000048d5",
			4649 => x"ff4248d5",
			4650 => x"0d088208",
			4651 => x"00038c04",
			4652 => x"00c448d5",
			4653 => x"000048d5",
			4654 => x"0c063008",
			4655 => x"05083004",
			4656 => x"000048d5",
			4657 => x"ff1e48d5",
			4658 => x"0100f304",
			4659 => x"000048d5",
			4660 => x"005648d5",
			4661 => x"00039670",
			4662 => x"0901dd4c",
			4663 => x"00030c2c",
			4664 => x"0002e618",
			4665 => x"0d084b0c",
			4666 => x"06013b04",
			4667 => x"000049b9",
			4668 => x"03093704",
			4669 => x"012d49b9",
			4670 => x"000049b9",
			4671 => x"05081f08",
			4672 => x"0c05f604",
			4673 => x"000049b9",
			4674 => x"fe9749b9",
			4675 => x"ffe149b9",
			4676 => x"0507b804",
			4677 => x"ff4b49b9",
			4678 => x"0309a308",
			4679 => x"09017d04",
			4680 => x"000049b9",
			4681 => x"017149b9",
			4682 => x"09018704",
			4683 => x"ff8349b9",
			4684 => x"005349b9",
			4685 => x"0706a11c",
			4686 => x"0a02170c",
			4687 => x"07062b04",
			4688 => x"000049b9",
			4689 => x"0d088d04",
			4690 => x"fe8949b9",
			4691 => x"000049b9",
			4692 => x"040a0108",
			4693 => x"07062e04",
			4694 => x"ff8349b9",
			4695 => x"00e249b9",
			4696 => x"06017404",
			4697 => x"fe9f49b9",
			4698 => x"000049b9",
			4699 => x"008849b9",
			4700 => x"00037810",
			4701 => x"06016b04",
			4702 => x"ff4149b9",
			4703 => x"03098704",
			4704 => x"000049b9",
			4705 => x"05086a04",
			4706 => x"015349b9",
			4707 => x"000049b9",
			4708 => x"0e0a1b04",
			4709 => x"fec249b9",
			4710 => x"06018d08",
			4711 => x"040abb04",
			4712 => x"000049b9",
			4713 => x"ffa349b9",
			4714 => x"0706b404",
			4715 => x"011d49b9",
			4716 => x"000049b9",
			4717 => x"fe8349b9",
			4718 => x"00039a64",
			4719 => x"06018c58",
			4720 => x"00032438",
			4721 => x"07066c1c",
			4722 => x"0507b80c",
			4723 => x"01010f08",
			4724 => x"07061304",
			4725 => x"ff334a85",
			4726 => x"00b14a85",
			4727 => x"fe494a85",
			4728 => x"0a01e908",
			4729 => x"0d082504",
			4730 => x"00e94a85",
			4731 => x"fee54a85",
			4732 => x"0f097104",
			4733 => x"01624a85",
			4734 => x"002e4a85",
			4735 => x"07067010",
			4736 => x"09018308",
			4737 => x"03094f04",
			4738 => x"00004a85",
			4739 => x"fde34a85",
			4740 => x"03099604",
			4741 => x"01494a85",
			4742 => x"fda34a85",
			4743 => x"0b071008",
			4744 => x"0b06ff04",
			4745 => x"01534a85",
			4746 => x"ff1c4a85",
			4747 => x"01d94a85",
			4748 => x"0e09400c",
			4749 => x"00032c08",
			4750 => x"0308f704",
			4751 => x"00004a85",
			4752 => x"fc944a85",
			4753 => x"fe7d4a85",
			4754 => x"0409ed04",
			4755 => x"019a4a85",
			4756 => x"0e098708",
			4757 => x"07064104",
			4758 => x"00914a85",
			4759 => x"fd714a85",
			4760 => x"00037004",
			4761 => x"00b44a85",
			4762 => x"fe9e4a85",
			4763 => x"0b074408",
			4764 => x"05080f04",
			4765 => x"00024a85",
			4766 => x"02754a85",
			4767 => x"ff524a85",
			4768 => x"fe6b4a85",
			4769 => x"0c05d504",
			4770 => x"fe9a4b9b",
			4771 => x"0507f63c",
			4772 => x"0507ea28",
			4773 => x"0507e418",
			4774 => x"01013610",
			4775 => x"07064208",
			4776 => x"00035304",
			4777 => x"00b64b9b",
			4778 => x"00004b9b",
			4779 => x"0507b804",
			4780 => x"fece4b9b",
			4781 => x"00034b9b",
			4782 => x"0d084a04",
			4783 => x"fe714b9b",
			4784 => x"00004b9b",
			4785 => x"0b06ed0c",
			4786 => x"00037d08",
			4787 => x"06013d04",
			4788 => x"00004b9b",
			4789 => x"01664b9b",
			4790 => x"00004b9b",
			4791 => x"00004b9b",
			4792 => x"0d083e04",
			4793 => x"00004b9b",
			4794 => x"01012e0c",
			4795 => x"0b06fe08",
			4796 => x"03094004",
			4797 => x"00004b9b",
			4798 => x"fe924b9b",
			4799 => x"00004b9b",
			4800 => x"00004b9b",
			4801 => x"05082120",
			4802 => x"0002dd0c",
			4803 => x"0d084b04",
			4804 => x"00004b9b",
			4805 => x"07065804",
			4806 => x"00004b9b",
			4807 => x"ffab4b9b",
			4808 => x"0101470c",
			4809 => x"04094504",
			4810 => x"00004b9b",
			4811 => x"0d087f04",
			4812 => x"013c4b9b",
			4813 => x"00004b9b",
			4814 => x"0d087f04",
			4815 => x"ffff4b9b",
			4816 => x"00004b9b",
			4817 => x"0100f310",
			4818 => x"02093508",
			4819 => x"04095904",
			4820 => x"ff9f4b9b",
			4821 => x"00cb4b9b",
			4822 => x"07068504",
			4823 => x"fedd4b9b",
			4824 => x"00004b9b",
			4825 => x"0d08b30c",
			4826 => x"00039608",
			4827 => x"0b070e04",
			4828 => x"00004b9b",
			4829 => x"012c4b9b",
			4830 => x"00004b9b",
			4831 => x"0c066608",
			4832 => x"05089404",
			4833 => x"ff1d4b9b",
			4834 => x"00004b9b",
			4835 => x"01012304",
			4836 => x"00464b9b",
			4837 => x"00004b9b",
			4838 => x"00004b9d",
			4839 => x"00004ba1",
			4840 => x"0c060f04",
			4841 => x"ffff4bb5",
			4842 => x"0c064d04",
			4843 => x"00064bb5",
			4844 => x"00004bb5",
			4845 => x"0b071008",
			4846 => x"0b06bc04",
			4847 => x"00004bc9",
			4848 => x"fff04bc9",
			4849 => x"00004bc9",
			4850 => x"00030208",
			4851 => x"0406ea04",
			4852 => x"00004bdd",
			4853 => x"00064bdd",
			4854 => x"00004bdd",
			4855 => x"00030c08",
			4856 => x"00022e04",
			4857 => x"00004bf1",
			4858 => x"00034bf1",
			4859 => x"00004bf1",
			4860 => x"0507e708",
			4861 => x"0506f104",
			4862 => x"00004c0d",
			4863 => x"00144c0d",
			4864 => x"05081f04",
			4865 => x"fff34c0d",
			4866 => x"00004c0d",
			4867 => x"0b06dd04",
			4868 => x"00004c29",
			4869 => x"02092808",
			4870 => x"0208ce04",
			4871 => x"00004c29",
			4872 => x"00334c29",
			4873 => x"00004c29",
			4874 => x"0209200c",
			4875 => x"04098708",
			4876 => x"0207c504",
			4877 => x"00004c4d",
			4878 => x"001d4c4d",
			4879 => x"00004c4d",
			4880 => x"02097b04",
			4881 => x"ffea4c4d",
			4882 => x"00004c4d",
			4883 => x"0003240c",
			4884 => x"0207c504",
			4885 => x"00004c71",
			4886 => x"02097804",
			4887 => x"00114c71",
			4888 => x"00004c71",
			4889 => x"020a5004",
			4890 => x"fff44c71",
			4891 => x"00004c71",
			4892 => x"0003020c",
			4893 => x"02092808",
			4894 => x"02090004",
			4895 => x"00004c9d",
			4896 => x"00324c9d",
			4897 => x"00004c9d",
			4898 => x"06019108",
			4899 => x"06014704",
			4900 => x"00004c9d",
			4901 => x"fffd4c9d",
			4902 => x"00004c9d",
			4903 => x"00037d10",
			4904 => x"0507e70c",
			4905 => x"07065a08",
			4906 => x"07061304",
			4907 => x"00004cc1",
			4908 => x"003b4cc1",
			4909 => x"00004cc1",
			4910 => x"00004cc1",
			4911 => x"00004cc1",
			4912 => x"0c063010",
			4913 => x"04091d04",
			4914 => x"00004ce5",
			4915 => x"06016f08",
			4916 => x"0c05de04",
			4917 => x"00004ce5",
			4918 => x"ffb54ce5",
			4919 => x"00004ce5",
			4920 => x"00004ce5",
			4921 => x"09017d08",
			4922 => x"0a017904",
			4923 => x"00004d11",
			4924 => x"ffda4d11",
			4925 => x"0a02740c",
			4926 => x"0a01e904",
			4927 => x"00004d11",
			4928 => x"09021d04",
			4929 => x"00174d11",
			4930 => x"00004d11",
			4931 => x"00004d11",
			4932 => x"0b06e004",
			4933 => x"00004d3d",
			4934 => x"05082108",
			4935 => x"0507e404",
			4936 => x"00004d3d",
			4937 => x"00464d3d",
			4938 => x"0b073308",
			4939 => x"0b06fe04",
			4940 => x"00004d3d",
			4941 => x"ffe24d3d",
			4942 => x"00004d3d",
			4943 => x"0901dd0c",
			4944 => x"09018008",
			4945 => x"09017a04",
			4946 => x"00004d71",
			4947 => x"00114d71",
			4948 => x"fffa4d71",
			4949 => x"05086a0c",
			4950 => x"09022408",
			4951 => x"0507a004",
			4952 => x"00004d71",
			4953 => x"001c4d71",
			4954 => x"00004d71",
			4955 => x"00004d71",
			4956 => x"0c05f608",
			4957 => x"0901e304",
			4958 => x"fffd4da5",
			4959 => x"00004da5",
			4960 => x"0b06dd04",
			4961 => x"00004da5",
			4962 => x"040a280c",
			4963 => x"0f08f904",
			4964 => x"00004da5",
			4965 => x"0100e704",
			4966 => x"00004da5",
			4967 => x"00504da5",
			4968 => x"00004da5",
			4969 => x"00037d14",
			4970 => x"0507e710",
			4971 => x"0901f40c",
			4972 => x"0506f104",
			4973 => x"00004dd1",
			4974 => x"00035b04",
			4975 => x"00374dd1",
			4976 => x"00004dd1",
			4977 => x"00004dd1",
			4978 => x"00004dd1",
			4979 => x"00004dd1",
			4980 => x"0c063014",
			4981 => x"04091d04",
			4982 => x"00004dfd",
			4983 => x"06016f0c",
			4984 => x"0c05de04",
			4985 => x"00004dfd",
			4986 => x"07062c04",
			4987 => x"00004dfd",
			4988 => x"ffbd4dfd",
			4989 => x"00004dfd",
			4990 => x"00004dfd",
			4991 => x"00032414",
			4992 => x"0f093d04",
			4993 => x"00004e41",
			4994 => x"0002ee04",
			4995 => x"00004e41",
			4996 => x"0c064d08",
			4997 => x"0b06cd04",
			4998 => x"00004e41",
			4999 => x"00b44e41",
			5000 => x"00004e41",
			5001 => x"0e098704",
			5002 => x"ffd94e41",
			5003 => x"0802e008",
			5004 => x"08029e04",
			5005 => x"00004e41",
			5006 => x"001d4e41",
			5007 => x"00004e41",
			5008 => x"0c063210",
			5009 => x"04091d04",
			5010 => x"00004e85",
			5011 => x"0e0a1b08",
			5012 => x"0b06cc04",
			5013 => x"00004e85",
			5014 => x"ffa34e85",
			5015 => x"00004e85",
			5016 => x"020a9310",
			5017 => x"0002e604",
			5018 => x"00004e85",
			5019 => x"0b06fe04",
			5020 => x"00004e85",
			5021 => x"0d090f04",
			5022 => x"00334e85",
			5023 => x"00004e85",
			5024 => x"00004e85",
			5025 => x"00037018",
			5026 => x"09017d04",
			5027 => x"00004ec1",
			5028 => x"0d080b04",
			5029 => x"00004ec1",
			5030 => x"0d087f0c",
			5031 => x"0a01e904",
			5032 => x"00004ec1",
			5033 => x"07063f04",
			5034 => x"00004ec1",
			5035 => x"00804ec1",
			5036 => x"00004ec1",
			5037 => x"06018d04",
			5038 => x"ffee4ec1",
			5039 => x"00004ec1",
			5040 => x"040a3a18",
			5041 => x"0a01ec04",
			5042 => x"00004efd",
			5043 => x"01013610",
			5044 => x"0100e704",
			5045 => x"00004efd",
			5046 => x"0b06be04",
			5047 => x"00004efd",
			5048 => x"0802bb04",
			5049 => x"005a4efd",
			5050 => x"00004efd",
			5051 => x"00004efd",
			5052 => x"06018804",
			5053 => x"fff74efd",
			5054 => x"00004efd",
			5055 => x"0e093308",
			5056 => x"0d075504",
			5057 => x"00004f39",
			5058 => x"fffe4f39",
			5059 => x"0d089a14",
			5060 => x"09018304",
			5061 => x"00004f39",
			5062 => x"0e0a860c",
			5063 => x"0d080e04",
			5064 => x"00004f39",
			5065 => x"09021b04",
			5066 => x"002c4f39",
			5067 => x"00004f39",
			5068 => x"00004f39",
			5069 => x"00004f39",
			5070 => x"06013e08",
			5071 => x"0c05f204",
			5072 => x"00004f75",
			5073 => x"005b4f75",
			5074 => x"07067014",
			5075 => x"0507e704",
			5076 => x"00004f75",
			5077 => x"0c06320c",
			5078 => x"09021208",
			5079 => x"0d083e04",
			5080 => x"00004f75",
			5081 => x"ffac4f75",
			5082 => x"00004f75",
			5083 => x"00004f75",
			5084 => x"00004f75",
			5085 => x"00037d18",
			5086 => x"0507e714",
			5087 => x"0901f410",
			5088 => x"0507ba04",
			5089 => x"00004fa9",
			5090 => x"09017a04",
			5091 => x"00004fa9",
			5092 => x"00035b04",
			5093 => x"005a4fa9",
			5094 => x"00004fa9",
			5095 => x"00004fa9",
			5096 => x"00004fa9",
			5097 => x"00004fa9",
			5098 => x"05082118",
			5099 => x"0c05f204",
			5100 => x"00004fdd",
			5101 => x"00038510",
			5102 => x"0c062e0c",
			5103 => x"07064604",
			5104 => x"00004fdd",
			5105 => x"07068304",
			5106 => x"00694fdd",
			5107 => x"00004fdd",
			5108 => x"00004fdd",
			5109 => x"00004fdd",
			5110 => x"00004fdd",
			5111 => x"0100f310",
			5112 => x"0e08fd04",
			5113 => x"00005029",
			5114 => x"05084d08",
			5115 => x"0d084c04",
			5116 => x"00005029",
			5117 => x"ffd95029",
			5118 => x"00005029",
			5119 => x"0c05f304",
			5120 => x"00005029",
			5121 => x"00037d10",
			5122 => x"0e093304",
			5123 => x"00005029",
			5124 => x"01014508",
			5125 => x"0507bb04",
			5126 => x"00005029",
			5127 => x"006e5029",
			5128 => x"00005029",
			5129 => x"00005029",
			5130 => x"04098714",
			5131 => x"08025a04",
			5132 => x"0000508d",
			5133 => x"0f09600c",
			5134 => x"0c05d504",
			5135 => x"0000508d",
			5136 => x"0f08dd04",
			5137 => x"0000508d",
			5138 => x"003a508d",
			5139 => x"0000508d",
			5140 => x"06018810",
			5141 => x"0706b70c",
			5142 => x"08026f04",
			5143 => x"0000508d",
			5144 => x"06018004",
			5145 => x"ff83508d",
			5146 => x"0000508d",
			5147 => x"0000508d",
			5148 => x"00039a0c",
			5149 => x"01015408",
			5150 => x"0901fc04",
			5151 => x"0000508d",
			5152 => x"0038508d",
			5153 => x"0000508d",
			5154 => x"0000508d",
			5155 => x"00030c18",
			5156 => x"0a01ec10",
			5157 => x"08024e04",
			5158 => x"000050f9",
			5159 => x"06014008",
			5160 => x"0f08e604",
			5161 => x"000050f9",
			5162 => x"ffb650f9",
			5163 => x"000050f9",
			5164 => x"0f08dd04",
			5165 => x"000050f9",
			5166 => x"001d50f9",
			5167 => x"0a021d0c",
			5168 => x"0b072008",
			5169 => x"06013e04",
			5170 => x"000050f9",
			5171 => x"ffa150f9",
			5172 => x"000050f9",
			5173 => x"0a025710",
			5174 => x"020a2d0c",
			5175 => x"0802db08",
			5176 => x"02093004",
			5177 => x"000050f9",
			5178 => x"002d50f9",
			5179 => x"000050f9",
			5180 => x"000050f9",
			5181 => x"000050f9",
			5182 => x"040a3a20",
			5183 => x"08025a08",
			5184 => x"0100e904",
			5185 => x"0000514d",
			5186 => x"ffff514d",
			5187 => x"07064004",
			5188 => x"0000514d",
			5189 => x"0100e704",
			5190 => x"0000514d",
			5191 => x"07066c0c",
			5192 => x"01012608",
			5193 => x"0d080104",
			5194 => x"0000514d",
			5195 => x"005f514d",
			5196 => x"0000514d",
			5197 => x"0000514d",
			5198 => x"01014908",
			5199 => x"0706c904",
			5200 => x"ffc2514d",
			5201 => x"0000514d",
			5202 => x"0000514d",
			5203 => x"0b06dc0c",
			5204 => x"0e094008",
			5205 => x"03097804",
			5206 => x"ffcd5199",
			5207 => x"00005199",
			5208 => x"00005199",
			5209 => x"040a2818",
			5210 => x"07064604",
			5211 => x"00005199",
			5212 => x"0100e504",
			5213 => x"00005199",
			5214 => x"0002dd04",
			5215 => x"00005199",
			5216 => x"04094504",
			5217 => x"00005199",
			5218 => x"02090004",
			5219 => x"00005199",
			5220 => x"007f5199",
			5221 => x"00005199",
			5222 => x"040a281c",
			5223 => x"0100e704",
			5224 => x"000051dd",
			5225 => x"0d080b04",
			5226 => x"000051dd",
			5227 => x"0309ef10",
			5228 => x"09017d04",
			5229 => x"000051dd",
			5230 => x"0f092a04",
			5231 => x"000051dd",
			5232 => x"01013504",
			5233 => x"006051dd",
			5234 => x"000051dd",
			5235 => x"000051dd",
			5236 => x"0901fc04",
			5237 => x"ffe051dd",
			5238 => x"000051dd",
			5239 => x"0f092a0c",
			5240 => x"0a01f208",
			5241 => x"07064104",
			5242 => x"00005249",
			5243 => x"ff925249",
			5244 => x"00005249",
			5245 => x"0c061418",
			5246 => x"0a021d0c",
			5247 => x"07067008",
			5248 => x"0c05de04",
			5249 => x"00005249",
			5250 => x"ffa25249",
			5251 => x"00005249",
			5252 => x"0a025708",
			5253 => x"07062804",
			5254 => x"00005249",
			5255 => x"00235249",
			5256 => x"00005249",
			5257 => x"0c064d10",
			5258 => x"0d08b30c",
			5259 => x"0100ed04",
			5260 => x"00005249",
			5261 => x"00039d04",
			5262 => x"00b65249",
			5263 => x"00005249",
			5264 => x"00005249",
			5265 => x"00005249",
			5266 => x"0507ba08",
			5267 => x"0e098704",
			5268 => x"ffc752ad",
			5269 => x"000052ad",
			5270 => x"0901b218",
			5271 => x"02091b0c",
			5272 => x"0e08d604",
			5273 => x"000052ad",
			5274 => x"0208db04",
			5275 => x"000052ad",
			5276 => x"001a52ad",
			5277 => x"0e097708",
			5278 => x"02092804",
			5279 => x"000052ad",
			5280 => x"ffcb52ad",
			5281 => x"000052ad",
			5282 => x"020a9310",
			5283 => x"09021d0c",
			5284 => x"0e092404",
			5285 => x"000052ad",
			5286 => x"07062604",
			5287 => x"000052ad",
			5288 => x"004f52ad",
			5289 => x"000052ad",
			5290 => x"000052ad",
			5291 => x"09017d0c",
			5292 => x"06013e04",
			5293 => x"00005301",
			5294 => x"0a01ec04",
			5295 => x"00005301",
			5296 => x"ffdf5301",
			5297 => x"00037d1c",
			5298 => x"07063f04",
			5299 => x"00005301",
			5300 => x"0c062e10",
			5301 => x"0d087f0c",
			5302 => x"05082e08",
			5303 => x"08025304",
			5304 => x"00005301",
			5305 => x"00755301",
			5306 => x"00005301",
			5307 => x"00005301",
			5308 => x"0c063204",
			5309 => x"fffe5301",
			5310 => x"00005301",
			5311 => x"00005301",
			5312 => x"0e09871c",
			5313 => x"0b072018",
			5314 => x"0408db04",
			5315 => x"0000533d",
			5316 => x"0a021d10",
			5317 => x"07062b04",
			5318 => x"0000533d",
			5319 => x"05081f08",
			5320 => x"07068504",
			5321 => x"ffac533d",
			5322 => x"0000533d",
			5323 => x"0000533d",
			5324 => x"0000533d",
			5325 => x"0000533d",
			5326 => x"0000533d",
			5327 => x"09017d04",
			5328 => x"00005379",
			5329 => x"040b2218",
			5330 => x"0c05f604",
			5331 => x"00005379",
			5332 => x"05088610",
			5333 => x"0a01e404",
			5334 => x"00005379",
			5335 => x"09021d08",
			5336 => x"0b06a504",
			5337 => x"00005379",
			5338 => x"00415379",
			5339 => x"00005379",
			5340 => x"00005379",
			5341 => x"00005379",
			5342 => x"0003891c",
			5343 => x"09017a04",
			5344 => x"000053b5",
			5345 => x"07064604",
			5346 => x"000053b5",
			5347 => x"0002e604",
			5348 => x"000053b5",
			5349 => x"0101540c",
			5350 => x"0c05dc04",
			5351 => x"000053b5",
			5352 => x"0100f304",
			5353 => x"000053b5",
			5354 => x"008653b5",
			5355 => x"000053b5",
			5356 => x"000053b5",
			5357 => x"09017a04",
			5358 => x"00005401",
			5359 => x"0409db18",
			5360 => x"05082114",
			5361 => x"0d087f10",
			5362 => x"0c062e0c",
			5363 => x"07064404",
			5364 => x"00005401",
			5365 => x"0a01e404",
			5366 => x"00005401",
			5367 => x"00835401",
			5368 => x"00005401",
			5369 => x"00005401",
			5370 => x"00005401",
			5371 => x"0901dd08",
			5372 => x"06015c04",
			5373 => x"00005401",
			5374 => x"ffd45401",
			5375 => x"00005401",
			5376 => x"0409db18",
			5377 => x"0f08f904",
			5378 => x"00005475",
			5379 => x"0309b010",
			5380 => x"06014104",
			5381 => x"00005475",
			5382 => x"07064404",
			5383 => x"00005475",
			5384 => x"0a022804",
			5385 => x"00ae5475",
			5386 => x"00005475",
			5387 => x"00005475",
			5388 => x"0309d810",
			5389 => x"0c05da04",
			5390 => x"00005475",
			5391 => x"0507ab04",
			5392 => x"00005475",
			5393 => x"0507f604",
			5394 => x"ff7d5475",
			5395 => x"00005475",
			5396 => x"01010204",
			5397 => x"00005475",
			5398 => x"0f0ac30c",
			5399 => x"01015408",
			5400 => x"0a027b04",
			5401 => x"00285475",
			5402 => x"00005475",
			5403 => x"00005475",
			5404 => x"00005475",
			5405 => x"040a0130",
			5406 => x"0d084b18",
			5407 => x"07063f04",
			5408 => x"00005501",
			5409 => x"09017a04",
			5410 => x"00005501",
			5411 => x"0b06f00c",
			5412 => x"0a01e404",
			5413 => x"00005501",
			5414 => x"0d080b04",
			5415 => x"00005501",
			5416 => x"00a45501",
			5417 => x"00005501",
			5418 => x"0b06f00c",
			5419 => x"0309b008",
			5420 => x"0f08f004",
			5421 => x"00005501",
			5422 => x"ffd05501",
			5423 => x"00005501",
			5424 => x"03098708",
			5425 => x"0f092a04",
			5426 => x"00005501",
			5427 => x"006f5501",
			5428 => x"00005501",
			5429 => x"0309d80c",
			5430 => x"0e09a208",
			5431 => x"00033504",
			5432 => x"00005501",
			5433 => x"ff6a5501",
			5434 => x"00005501",
			5435 => x"00037008",
			5436 => x"00033e04",
			5437 => x"00005501",
			5438 => x"00525501",
			5439 => x"00005501",
			5440 => x"00037d28",
			5441 => x"09017a08",
			5442 => x"07067204",
			5443 => x"fe6a5585",
			5444 => x"013e5585",
			5445 => x"0d080108",
			5446 => x"0208e204",
			5447 => x"030e5585",
			5448 => x"fe625585",
			5449 => x"0d08da14",
			5450 => x"0802d20c",
			5451 => x"06013804",
			5452 => x"fe9e5585",
			5453 => x"040a3a04",
			5454 => x"044d5585",
			5455 => x"03145585",
			5456 => x"040a9504",
			5457 => x"04b55585",
			5458 => x"09ba5585",
			5459 => x"fe605585",
			5460 => x"00039514",
			5461 => x"0802e90c",
			5462 => x"0802e504",
			5463 => x"fe5b5585",
			5464 => x"040ae204",
			5465 => x"01ee5585",
			5466 => x"fe7a5585",
			5467 => x"06019104",
			5468 => x"fec25585",
			5469 => x"07865585",
			5470 => x"00039a04",
			5471 => x"feb05585",
			5472 => x"fe5a5585",
			5473 => x"09018314",
			5474 => x"0a01f70c",
			5475 => x"03098708",
			5476 => x"0307f404",
			5477 => x"00005611",
			5478 => x"000a5611",
			5479 => x"00005611",
			5480 => x"0100ef04",
			5481 => x"ffa05611",
			5482 => x"00005611",
			5483 => x"0f096010",
			5484 => x"00031a0c",
			5485 => x"0d088208",
			5486 => x"0d07f104",
			5487 => x"00005611",
			5488 => x"00a75611",
			5489 => x"00005611",
			5490 => x"00005611",
			5491 => x"0309780c",
			5492 => x"0f097d08",
			5493 => x"0507d804",
			5494 => x"00005611",
			5495 => x"ff7b5611",
			5496 => x"00005611",
			5497 => x"00037810",
			5498 => x"00031a04",
			5499 => x"00005611",
			5500 => x"0507c904",
			5501 => x"00005611",
			5502 => x"0901a904",
			5503 => x"00005611",
			5504 => x"00a05611",
			5505 => x"030a4904",
			5506 => x"fff65611",
			5507 => x"00005611",
			5508 => x"040a2828",
			5509 => x"0f097d24",
			5510 => x"07065b14",
			5511 => x"04091d04",
			5512 => x"0000567d",
			5513 => x"0d08650c",
			5514 => x"07062b04",
			5515 => x"0000567d",
			5516 => x"0b06bc04",
			5517 => x"0000567d",
			5518 => x"ffa6567d",
			5519 => x"0000567d",
			5520 => x"0002dd04",
			5521 => x"0000567d",
			5522 => x"09017d04",
			5523 => x"0000567d",
			5524 => x"07068604",
			5525 => x"0068567d",
			5526 => x"0000567d",
			5527 => x"00b6567d",
			5528 => x"0901fc0c",
			5529 => x"0c06e508",
			5530 => x"08029904",
			5531 => x"0000567d",
			5532 => x"ffa1567d",
			5533 => x"0000567d",
			5534 => x"0000567d",
			5535 => x"040a012c",
			5536 => x"0b06cd14",
			5537 => x"02096010",
			5538 => x"0901a904",
			5539 => x"00005711",
			5540 => x"0c05bd04",
			5541 => x"00005711",
			5542 => x"0d080a04",
			5543 => x"00005711",
			5544 => x"ff7a5711",
			5545 => x"00005711",
			5546 => x"0d081704",
			5547 => x"00005711",
			5548 => x"0100e704",
			5549 => x"00005711",
			5550 => x"0209950c",
			5551 => x"0d087f08",
			5552 => x"08025304",
			5553 => x"00005711",
			5554 => x"00915711",
			5555 => x"00005711",
			5556 => x"00005711",
			5557 => x"0601770c",
			5558 => x"0c063408",
			5559 => x"00033504",
			5560 => x"00005711",
			5561 => x"ff495711",
			5562 => x"00005711",
			5563 => x"00037d0c",
			5564 => x"020a2d08",
			5565 => x"0f09c604",
			5566 => x"00005711",
			5567 => x"00735711",
			5568 => x"00005711",
			5569 => x"0802f304",
			5570 => x"00005711",
			5571 => x"00005711",
			5572 => x"040a0130",
			5573 => x"07066c18",
			5574 => x"0c05d704",
			5575 => x"00005785",
			5576 => x"0901db10",
			5577 => x"0100eb04",
			5578 => x"00005785",
			5579 => x"0c062e08",
			5580 => x"0b069c04",
			5581 => x"00005785",
			5582 => x"00815785",
			5583 => x"00005785",
			5584 => x"00005785",
			5585 => x"0b071014",
			5586 => x"05082e10",
			5587 => x"0507ea04",
			5588 => x"00005785",
			5589 => x"0c05f804",
			5590 => x"00005785",
			5591 => x"0c063204",
			5592 => x"ff8f5785",
			5593 => x"00005785",
			5594 => x"00005785",
			5595 => x"00005785",
			5596 => x"0c063308",
			5597 => x"06018804",
			5598 => x"ff755785",
			5599 => x"00005785",
			5600 => x"00005785",
			5601 => x"0d084b18",
			5602 => x"00035310",
			5603 => x"09017a04",
			5604 => x"00005819",
			5605 => x"0b06f008",
			5606 => x"0d080104",
			5607 => x"00005819",
			5608 => x"00c75819",
			5609 => x"00005819",
			5610 => x"0309ef04",
			5611 => x"ffd85819",
			5612 => x"00005819",
			5613 => x"0507f50c",
			5614 => x"08029108",
			5615 => x"0c05f404",
			5616 => x"00005819",
			5617 => x"ff4c5819",
			5618 => x"00005819",
			5619 => x"0d088214",
			5620 => x"0c05f704",
			5621 => x"00005819",
			5622 => x"02090004",
			5623 => x"00005819",
			5624 => x"0b071e08",
			5625 => x"00039604",
			5626 => x"00cf5819",
			5627 => x"00005819",
			5628 => x"00005819",
			5629 => x"0309c004",
			5630 => x"00005819",
			5631 => x"0c06660c",
			5632 => x"05082104",
			5633 => x"00005819",
			5634 => x"05089404",
			5635 => x"ff765819",
			5636 => x"00005819",
			5637 => x"00005819",
			5638 => x"06013e10",
			5639 => x"0c05f204",
			5640 => x"000058a5",
			5641 => x"0c063008",
			5642 => x"0100ef04",
			5643 => x"006158a5",
			5644 => x"000058a5",
			5645 => x"000058a5",
			5646 => x"07067020",
			5647 => x"0901c314",
			5648 => x"0507e704",
			5649 => x"000058a5",
			5650 => x"0d08720c",
			5651 => x"0c05f404",
			5652 => x"000058a5",
			5653 => x"0d083e04",
			5654 => x"000058a5",
			5655 => x"ff6558a5",
			5656 => x"000058a5",
			5657 => x"01013d08",
			5658 => x"07061704",
			5659 => x"000058a5",
			5660 => x"001e58a5",
			5661 => x"000058a5",
			5662 => x"0c060f04",
			5663 => x"000058a5",
			5664 => x"0d08da10",
			5665 => x"0c06500c",
			5666 => x"0d08b308",
			5667 => x"0601a304",
			5668 => x"009958a5",
			5669 => x"000058a5",
			5670 => x"000058a5",
			5671 => x"000058a5",
			5672 => x"000058a5",
			5673 => x"0003853c",
			5674 => x"0100e710",
			5675 => x"0600ef08",
			5676 => x"0f067a04",
			5677 => x"fea35939",
			5678 => x"02e45939",
			5679 => x"09017a04",
			5680 => x"fe565939",
			5681 => x"00005939",
			5682 => x"0d08da24",
			5683 => x"0d080e0c",
			5684 => x"0002e604",
			5685 => x"01d95939",
			5686 => x"0507c704",
			5687 => x"fe475939",
			5688 => x"004a5939",
			5689 => x"0a01e40c",
			5690 => x"03090708",
			5691 => x"08023c04",
			5692 => x"00005939",
			5693 => x"00e75939",
			5694 => x"fe6e5939",
			5695 => x"06018c08",
			5696 => x"00034b04",
			5697 => x"017e5939",
			5698 => x"00a25939",
			5699 => x"03145939",
			5700 => x"07071204",
			5701 => x"fe6a5939",
			5702 => x"00f15939",
			5703 => x"0003960c",
			5704 => x"0802eb04",
			5705 => x"fe6b5939",
			5706 => x"06019404",
			5707 => x"00005939",
			5708 => x"02825939",
			5709 => x"fe645939",
			5710 => x"0f092a0c",
			5711 => x"09018308",
			5712 => x"0100ef04",
			5713 => x"ff9759c5",
			5714 => x"000059c5",
			5715 => x"000059c5",
			5716 => x"0c061424",
			5717 => x"06016b14",
			5718 => x"07067010",
			5719 => x"0507d804",
			5720 => x"000059c5",
			5721 => x"06013e04",
			5722 => x"000059c5",
			5723 => x"0c05f404",
			5724 => x"000059c5",
			5725 => x"ff6f59c5",
			5726 => x"000059c5",
			5727 => x"0706580c",
			5728 => x"00037d08",
			5729 => x"07062804",
			5730 => x"000059c5",
			5731 => x"002b59c5",
			5732 => x"000059c5",
			5733 => x"000059c5",
			5734 => x"0d08da14",
			5735 => x"0100e904",
			5736 => x"000059c5",
			5737 => x"0c064d0c",
			5738 => x"0d08b308",
			5739 => x"0e08fd04",
			5740 => x"000059c5",
			5741 => x"00ab59c5",
			5742 => x"000059c5",
			5743 => x"000059c5",
			5744 => x"000059c5",
			5745 => x"0901b82c",
			5746 => x"00030c24",
			5747 => x"0a01f21c",
			5748 => x"0d084b10",
			5749 => x"0507f50c",
			5750 => x"0100aa04",
			5751 => x"00005a79",
			5752 => x"03093704",
			5753 => x"005b5a79",
			5754 => x"00005a79",
			5755 => x"00005a79",
			5756 => x"0d086d08",
			5757 => x"0208db04",
			5758 => x"00005a79",
			5759 => x"ff505a79",
			5760 => x"00005a79",
			5761 => x"0100ed04",
			5762 => x"00005a79",
			5763 => x"00b15a79",
			5764 => x"0c066604",
			5765 => x"ff455a79",
			5766 => x"00005a79",
			5767 => x"0003530c",
			5768 => x"03094f04",
			5769 => x"00005a79",
			5770 => x"0507bc04",
			5771 => x"00005a79",
			5772 => x"011d5a79",
			5773 => x"0e0a1b10",
			5774 => x"07066d0c",
			5775 => x"0c05d904",
			5776 => x"00005a79",
			5777 => x"06019404",
			5778 => x"ff7f5a79",
			5779 => x"00005a79",
			5780 => x"00005a79",
			5781 => x"040af710",
			5782 => x"0c05f604",
			5783 => x"00005a79",
			5784 => x"0d084a04",
			5785 => x"00005a79",
			5786 => x"09021d04",
			5787 => x"00dc5a79",
			5788 => x"00005a79",
			5789 => x"00005a79",
			5790 => x"0d084b20",
			5791 => x"00035318",
			5792 => x"09017a04",
			5793 => x"00005b1d",
			5794 => x"07063f04",
			5795 => x"00005b1d",
			5796 => x"0b06f00c",
			5797 => x"0d080104",
			5798 => x"00005b1d",
			5799 => x"05080104",
			5800 => x"00e25b1d",
			5801 => x"00005b1d",
			5802 => x"00005b1d",
			5803 => x"0309ef04",
			5804 => x"ffd95b1d",
			5805 => x"00005b1d",
			5806 => x"0507f50c",
			5807 => x"08029108",
			5808 => x"0c05f404",
			5809 => x"00005b1d",
			5810 => x"ff5e5b1d",
			5811 => x"00005b1d",
			5812 => x"0d088214",
			5813 => x"0c05f704",
			5814 => x"00005b1d",
			5815 => x"0002e604",
			5816 => x"00005b1d",
			5817 => x"00039608",
			5818 => x"0c064d04",
			5819 => x"00bb5b1d",
			5820 => x"00005b1d",
			5821 => x"00005b1d",
			5822 => x"0309ef04",
			5823 => x"00005b1d",
			5824 => x"0c06660c",
			5825 => x"05082104",
			5826 => x"00005b1d",
			5827 => x"05089404",
			5828 => x"ff715b1d",
			5829 => x"00005b1d",
			5830 => x"00005b1d",
			5831 => x"0003893c",
			5832 => x"0901760c",
			5833 => x"0600ef08",
			5834 => x"0100a604",
			5835 => x"fe945ba9",
			5836 => x"01e95ba9",
			5837 => x"fe665ba9",
			5838 => x"0507b808",
			5839 => x"01010b04",
			5840 => x"01195ba9",
			5841 => x"fe415ba9",
			5842 => x"05084d18",
			5843 => x"06018c10",
			5844 => x"0c05d908",
			5845 => x"00034604",
			5846 => x"01095ba9",
			5847 => x"fdff5ba9",
			5848 => x"0a01e404",
			5849 => x"ff875ba9",
			5850 => x"018f5ba9",
			5851 => x"05082e04",
			5852 => x"03c65ba9",
			5853 => x"02685ba9",
			5854 => x"040a2804",
			5855 => x"01f15ba9",
			5856 => x"07072408",
			5857 => x"0706b404",
			5858 => x"fd505ba9",
			5859 => x"feb85ba9",
			5860 => x"01115ba9",
			5861 => x"00039508",
			5862 => x"06019404",
			5863 => x"fe6c5ba9",
			5864 => x"01875ba9",
			5865 => x"fe635ba9",
			5866 => x"0409a024",
			5867 => x"0c05d704",
			5868 => x"00005c5d",
			5869 => x"07066c10",
			5870 => x"0101110c",
			5871 => x"0100eb04",
			5872 => x"00005c5d",
			5873 => x"09017a04",
			5874 => x"00005c5d",
			5875 => x"00fd5c5d",
			5876 => x"00005c5d",
			5877 => x"0002e608",
			5878 => x"0002dd04",
			5879 => x"00005c5d",
			5880 => x"ffb15c5d",
			5881 => x"0002ee04",
			5882 => x"00005c5d",
			5883 => x"004d5c5d",
			5884 => x"03097810",
			5885 => x"0c06130c",
			5886 => x"07065908",
			5887 => x"0e096204",
			5888 => x"feda5c5d",
			5889 => x"00005c5d",
			5890 => x"00005c5d",
			5891 => x"00005c5d",
			5892 => x"02099508",
			5893 => x"0100f304",
			5894 => x"00005c5d",
			5895 => x"00ed5c5d",
			5896 => x"0e09870c",
			5897 => x"0c061208",
			5898 => x"07064104",
			5899 => x"00005c5d",
			5900 => x"ff045c5d",
			5901 => x"00005c5d",
			5902 => x"0209c104",
			5903 => x"00a35c5d",
			5904 => x"0b071e08",
			5905 => x"07066d04",
			5906 => x"ffcb5c5d",
			5907 => x"00795c5d",
			5908 => x"0c066a04",
			5909 => x"ff425c5d",
			5910 => x"00005c5d",
			5911 => x"0901c338",
			5912 => x"00030228",
			5913 => x"0309781c",
			5914 => x"0a01ec14",
			5915 => x"04091d0c",
			5916 => x"0507e608",
			5917 => x"0c05f204",
			5918 => x"00005d29",
			5919 => x"004f5d29",
			5920 => x"00005d29",
			5921 => x"04094504",
			5922 => x"ff995d29",
			5923 => x"00005d29",
			5924 => x"09017a04",
			5925 => x"00005d29",
			5926 => x"00cf5d29",
			5927 => x"0c062e08",
			5928 => x"08026404",
			5929 => x"ff625d29",
			5930 => x"00005d29",
			5931 => x"00005d29",
			5932 => x"0c06660c",
			5933 => x"08026f04",
			5934 => x"00005d29",
			5935 => x"0a01fa04",
			5936 => x"00005d29",
			5937 => x"ff375d29",
			5938 => x"00005d29",
			5939 => x"0a021d08",
			5940 => x"0901cc04",
			5941 => x"00005d29",
			5942 => x"ff605d29",
			5943 => x"00037d1c",
			5944 => x"0507ca10",
			5945 => x"07064108",
			5946 => x"07062e04",
			5947 => x"00005d29",
			5948 => x"00465d29",
			5949 => x"040a0104",
			5950 => x"00005d29",
			5951 => x"ff9d5d29",
			5952 => x"030a7808",
			5953 => x"09021504",
			5954 => x"00cf5d29",
			5955 => x"00005d29",
			5956 => x"00005d29",
			5957 => x"030a4908",
			5958 => x"0802eb04",
			5959 => x"ff905d29",
			5960 => x"00005d29",
			5961 => x"00005d29",
			5962 => x"00038944",
			5963 => x"0100e814",
			5964 => x"0a01790c",
			5965 => x"02066104",
			5966 => x"ff235ddd",
			5967 => x"09011b04",
			5968 => x"01045ddd",
			5969 => x"00005ddd",
			5970 => x"09017d04",
			5971 => x"fe735ddd",
			5972 => x"00005ddd",
			5973 => x"00035318",
			5974 => x"0802b310",
			5975 => x"0101360c",
			5976 => x"0309ef08",
			5977 => x"0d084b04",
			5978 => x"01405ddd",
			5979 => x"009b5ddd",
			5980 => x"ff455ddd",
			5981 => x"fc2a5ddd",
			5982 => x"0309a304",
			5983 => x"00005ddd",
			5984 => x"01fd5ddd",
			5985 => x"0309d804",
			5986 => x"fdd95ddd",
			5987 => x"0d088208",
			5988 => x"0b06dd04",
			5989 => x"00005ddd",
			5990 => x"01895ddd",
			5991 => x"0a026408",
			5992 => x"040a8804",
			5993 => x"003d5ddd",
			5994 => x"fead5ddd",
			5995 => x"01105ddd",
			5996 => x"00039514",
			5997 => x"00039104",
			5998 => x"feff5ddd",
			5999 => x"0101570c",
			6000 => x"09021504",
			6001 => x"ffbf5ddd",
			6002 => x"01015104",
			6003 => x"00dc5ddd",
			6004 => x"00005ddd",
			6005 => x"ff885ddd",
			6006 => x"fe675ddd",
			6007 => x"00037840",
			6008 => x"09017a14",
			6009 => x"0100eb10",
			6010 => x"0600ef08",
			6011 => x"0100a304",
			6012 => x"fe765ea1",
			6013 => x"097e5ea1",
			6014 => x"0b070104",
			6015 => x"fe625ea1",
			6016 => x"ffb85ea1",
			6017 => x"01cc5ea1",
			6018 => x"0507b80c",
			6019 => x"03098708",
			6020 => x"01010b04",
			6021 => x"01f65ea1",
			6022 => x"fe585ea1",
			6023 => x"04d35ea1",
			6024 => x"030a781c",
			6025 => x"0100eb0c",
			6026 => x"0a01ec08",
			6027 => x"0507e604",
			6028 => x"04f05ea1",
			6029 => x"fe4c5ea1",
			6030 => x"024e5ea1",
			6031 => x"00035308",
			6032 => x"09017d04",
			6033 => x"05125ea1",
			6034 => x"029d5ea1",
			6035 => x"0309d804",
			6036 => x"fdc35ea1",
			6037 => x"02bf5ea1",
			6038 => x"fe885ea1",
			6039 => x"00038910",
			6040 => x"0802e80c",
			6041 => x"040abb08",
			6042 => x"0802db04",
			6043 => x"fe7b5ea1",
			6044 => x"01395ea1",
			6045 => x"fe645ea1",
			6046 => x"06dc5ea1",
			6047 => x"00039a10",
			6048 => x"0802f10c",
			6049 => x"06019604",
			6050 => x"fe615ea1",
			6051 => x"0802eb04",
			6052 => x"fee65ea1",
			6053 => x"00555ea1",
			6054 => x"04725ea1",
			6055 => x"fe5e5ea1",
			6056 => x"0901b834",
			6057 => x"00030c2c",
			6058 => x"0a01f21c",
			6059 => x"0d084b10",
			6060 => x"0b06ef0c",
			6061 => x"0100aa04",
			6062 => x"00005f65",
			6063 => x"03093704",
			6064 => x"00485f65",
			6065 => x"00005f65",
			6066 => x"00005f65",
			6067 => x"0d086d08",
			6068 => x"09017a04",
			6069 => x"00005f65",
			6070 => x"ff4d5f65",
			6071 => x"00005f65",
			6072 => x"0309a30c",
			6073 => x"07063d04",
			6074 => x"00005f65",
			6075 => x"0f08f004",
			6076 => x"00005f65",
			6077 => x"00c95f65",
			6078 => x"00005f65",
			6079 => x"0c066604",
			6080 => x"ff585f65",
			6081 => x"00005f65",
			6082 => x"00036818",
			6083 => x"03094f04",
			6084 => x"00005f65",
			6085 => x"0c05f30c",
			6086 => x"0c05da08",
			6087 => x"0c05d404",
			6088 => x"00005f65",
			6089 => x"00185f65",
			6090 => x"00005f65",
			6091 => x"0d080e04",
			6092 => x"00005f65",
			6093 => x"01115f65",
			6094 => x"030a1204",
			6095 => x"ffab5f65",
			6096 => x"040af710",
			6097 => x"06018804",
			6098 => x"00005f65",
			6099 => x"040aa904",
			6100 => x"00005f65",
			6101 => x"030a9904",
			6102 => x"00a75f65",
			6103 => x"00005f65",
			6104 => x"00005f65",
			6105 => x"00038940",
			6106 => x"030a1230",
			6107 => x"00036328",
			6108 => x"0901dd20",
			6109 => x"0f096010",
			6110 => x"0100eb08",
			6111 => x"06014104",
			6112 => x"ff645ff1",
			6113 => x"00005ff1",
			6114 => x"0b070e04",
			6115 => x"009a5ff1",
			6116 => x"ffe75ff1",
			6117 => x"0c061308",
			6118 => x"0901c304",
			6119 => x"fecf5ff1",
			6120 => x"ffe45ff1",
			6121 => x"01010204",
			6122 => x"ffaa5ff1",
			6123 => x"00fd5ff1",
			6124 => x"03097804",
			6125 => x"00005ff1",
			6126 => x"01505ff1",
			6127 => x"0c05f404",
			6128 => x"00005ff1",
			6129 => x"feab5ff1",
			6130 => x"020a2d04",
			6131 => x"01465ff1",
			6132 => x"0d088d04",
			6133 => x"00525ff1",
			6134 => x"020a5b04",
			6135 => x"ffb15ff1",
			6136 => x"00005ff1",
			6137 => x"09021504",
			6138 => x"fe895ff1",
			6139 => x"00005ff1",
			6140 => x"00037d40",
			6141 => x"09017a10",
			6142 => x"0b07010c",
			6143 => x"0600ef08",
			6144 => x"0100a604",
			6145 => x"fe8760a5",
			6146 => x"024d60a5",
			6147 => x"fe6560a5",
			6148 => x"000060a5",
			6149 => x"0b06a508",
			6150 => x"0208e904",
			6151 => x"002860a5",
			6152 => x"fe7460a5",
			6153 => x"0d08b320",
			6154 => x"0100ed10",
			6155 => x"07066f08",
			6156 => x"0507f504",
			6157 => x"012360a5",
			6158 => x"febb60a5",
			6159 => x"0b071004",
			6160 => x"014160a5",
			6161 => x"031e60a5",
			6162 => x"00035308",
			6163 => x"0d07f104",
			6164 => x"ff3260a5",
			6165 => x"01d960a5",
			6166 => x"0309d804",
			6167 => x"fdc260a5",
			6168 => x"022460a5",
			6169 => x"00035b04",
			6170 => x"002b60a5",
			6171 => x"fe7460a5",
			6172 => x"00039618",
			6173 => x"0802eb10",
			6174 => x"0003810c",
			6175 => x"01014708",
			6176 => x"0308d604",
			6177 => x"000060a5",
			6178 => x"03a960a5",
			6179 => x"fea660a5",
			6180 => x"fe6760a5",
			6181 => x"06019404",
			6182 => x"001460a5",
			6183 => x"02fd60a5",
			6184 => x"fe6260a5",
			6185 => x"0409db40",
			6186 => x"0a01f220",
			6187 => x"0d084b08",
			6188 => x"09017d04",
			6189 => x"00006199",
			6190 => x"007f6199",
			6191 => x"02090c0c",
			6192 => x"08025a08",
			6193 => x"0c05f304",
			6194 => x"00006199",
			6195 => x"feda6199",
			6196 => x"00006199",
			6197 => x"03098708",
			6198 => x"0c061a04",
			6199 => x"00006199",
			6200 => x"00c66199",
			6201 => x"ffa46199",
			6202 => x"0309c018",
			6203 => x"0d080e08",
			6204 => x"00030c04",
			6205 => x"00006199",
			6206 => x"ffb86199",
			6207 => x"0100ed04",
			6208 => x"00006199",
			6209 => x"01012608",
			6210 => x"03093704",
			6211 => x"00006199",
			6212 => x"01596199",
			6213 => x"00006199",
			6214 => x"0b072f04",
			6215 => x"ffa56199",
			6216 => x"00006199",
			6217 => x"01011f14",
			6218 => x"0c06340c",
			6219 => x"08028704",
			6220 => x"00006199",
			6221 => x"0901ce04",
			6222 => x"fe856199",
			6223 => x"00006199",
			6224 => x"0802b704",
			6225 => x"009b6199",
			6226 => x"00006199",
			6227 => x"00034b08",
			6228 => x"03099604",
			6229 => x"ffaa6199",
			6230 => x"01226199",
			6231 => x"0309d808",
			6232 => x"0b06bd04",
			6233 => x"00006199",
			6234 => x"fecf6199",
			6235 => x"00037008",
			6236 => x"01014904",
			6237 => x"00dd6199",
			6238 => x"00006199",
			6239 => x"0e0a1b08",
			6240 => x"00037804",
			6241 => x"00006199",
			6242 => x"fef86199",
			6243 => x"06019104",
			6244 => x"00006199",
			6245 => x"009b6199",
			6246 => x"040a0140",
			6247 => x"0a021d38",
			6248 => x"01011b30",
			6249 => x"07065b1c",
			6250 => x"04091d0c",
			6251 => x"03091a08",
			6252 => x"0c05ba04",
			6253 => x"0000625d",
			6254 => x"0033625d",
			6255 => x"0000625d",
			6256 => x"06015208",
			6257 => x"0b06cc04",
			6258 => x"0000625d",
			6259 => x"ff4a625d",
			6260 => x"02091304",
			6261 => x"0000625d",
			6262 => x"000b625d",
			6263 => x"07066c08",
			6264 => x"0100eb04",
			6265 => x"0000625d",
			6266 => x"00a1625d",
			6267 => x"0100f308",
			6268 => x"0100eb04",
			6269 => x"0000625d",
			6270 => x"ffd9625d",
			6271 => x"0028625d",
			6272 => x"0c05f304",
			6273 => x"0000625d",
			6274 => x"ff4f625d",
			6275 => x"03094f04",
			6276 => x"0000625d",
			6277 => x"00da625d",
			6278 => x"06017c0c",
			6279 => x"00033504",
			6280 => x"0000625d",
			6281 => x"0c066d04",
			6282 => x"ff09625d",
			6283 => x"0000625d",
			6284 => x"00037d10",
			6285 => x"07063d04",
			6286 => x"0000625d",
			6287 => x"0b073308",
			6288 => x"0309c004",
			6289 => x"0000625d",
			6290 => x"00d3625d",
			6291 => x"0000625d",
			6292 => x"06019104",
			6293 => x"ffab625d",
			6294 => x"0000625d",
			6295 => x"0409db44",
			6296 => x"0a01f224",
			6297 => x"0d084b08",
			6298 => x"09017d04",
			6299 => x"00006341",
			6300 => x"00826341",
			6301 => x"02090c0c",
			6302 => x"08025a08",
			6303 => x"0c05f304",
			6304 => x"00006341",
			6305 => x"febe6341",
			6306 => x"00006341",
			6307 => x"03097808",
			6308 => x"0c061a04",
			6309 => x"00006341",
			6310 => x"00c76341",
			6311 => x"0b071004",
			6312 => x"ff776341",
			6313 => x"00006341",
			6314 => x"0309c018",
			6315 => x"0d082210",
			6316 => x"0c05f608",
			6317 => x"0a020004",
			6318 => x"00006341",
			6319 => x"ff966341",
			6320 => x"0c05f704",
			6321 => x"00506341",
			6322 => x"00006341",
			6323 => x"0100ed04",
			6324 => x"00006341",
			6325 => x"01656341",
			6326 => x"0b072f04",
			6327 => x"ff826341",
			6328 => x"00006341",
			6329 => x"0e098708",
			6330 => x"0b06ee04",
			6331 => x"feb96341",
			6332 => x"00006341",
			6333 => x"040a2804",
			6334 => x"011e6341",
			6335 => x"01011b08",
			6336 => x"0c066a04",
			6337 => x"fe956341",
			6338 => x"00006341",
			6339 => x"030a4910",
			6340 => x"00037008",
			6341 => x"0209dd04",
			6342 => x"00006341",
			6343 => x"00d26341",
			6344 => x"0e0a1b04",
			6345 => x"fede6341",
			6346 => x"00006341",
			6347 => x"0f0ac308",
			6348 => x"00039a04",
			6349 => x"010c6341",
			6350 => x"00006341",
			6351 => x"00006341",
			6352 => x"0901dd50",
			6353 => x"0003243c",
			6354 => x"0d083e10",
			6355 => x"0d081808",
			6356 => x"0901a904",
			6357 => x"0000643d",
			6358 => x"fff5643d",
			6359 => x"09017d04",
			6360 => x"0000643d",
			6361 => x"010e643d",
			6362 => x"0b06ec10",
			6363 => x"0b06cc04",
			6364 => x"0000643d",
			6365 => x"0a021708",
			6366 => x"0208dd04",
			6367 => x"0000643d",
			6368 => x"feef643d",
			6369 => x"0000643d",
			6370 => x"06014110",
			6371 => x"0100e808",
			6372 => x"0b06fe04",
			6373 => x"0000643d",
			6374 => x"005f643d",
			6375 => x"0c063204",
			6376 => x"ff3e643d",
			6377 => x"0000643d",
			6378 => x"0309c008",
			6379 => x"09017d04",
			6380 => x"0000643d",
			6381 => x"00e8643d",
			6382 => x"0000643d",
			6383 => x"0c065008",
			6384 => x"01012a04",
			6385 => x"ff08643d",
			6386 => x"0000643d",
			6387 => x"01010204",
			6388 => x"0000643d",
			6389 => x"01012304",
			6390 => x"001b643d",
			6391 => x"0000643d",
			6392 => x"00036810",
			6393 => x"06016f04",
			6394 => x"0000643d",
			6395 => x"03098704",
			6396 => x"0000643d",
			6397 => x"0b071e04",
			6398 => x"0114643d",
			6399 => x"0000643d",
			6400 => x"0e0a1b0c",
			6401 => x"0c05f404",
			6402 => x"0000643d",
			6403 => x"030a5c04",
			6404 => x"ff6a643d",
			6405 => x"0000643d",
			6406 => x"0f0ac310",
			6407 => x"06018d04",
			6408 => x"0000643d",
			6409 => x"0c05f804",
			6410 => x"0000643d",
			6411 => x"030a2804",
			6412 => x"0000643d",
			6413 => x"00e0643d",
			6414 => x"0000643d",
			6415 => x"07063f14",
			6416 => x"0409870c",
			6417 => x"01011108",
			6418 => x"0100aa04",
			6419 => x"00006521",
			6420 => x"003d6521",
			6421 => x"00006521",
			6422 => x"06016b04",
			6423 => x"fe8c6521",
			6424 => x"00006521",
			6425 => x"07065828",
			6426 => x"06016c1c",
			6427 => x"040a0118",
			6428 => x"0a01f20c",
			6429 => x"06013e04",
			6430 => x"00006521",
			6431 => x"0f08f004",
			6432 => x"00006521",
			6433 => x"ffa56521",
			6434 => x"09018b04",
			6435 => x"00006521",
			6436 => x"03094f04",
			6437 => x"00006521",
			6438 => x"00e16521",
			6439 => x"ff756521",
			6440 => x"00037d08",
			6441 => x"03099604",
			6442 => x"00006521",
			6443 => x"01406521",
			6444 => x"fffb6521",
			6445 => x"0b06dd10",
			6446 => x"0b06cc04",
			6447 => x"00006521",
			6448 => x"0309b008",
			6449 => x"0f08f004",
			6450 => x"00006521",
			6451 => x"fec16521",
			6452 => x"00006521",
			6453 => x"040a2814",
			6454 => x"0100f310",
			6455 => x"03097808",
			6456 => x"0c063004",
			6457 => x"009a6521",
			6458 => x"00006521",
			6459 => x"07068504",
			6460 => x"ff886521",
			6461 => x"00006521",
			6462 => x"01146521",
			6463 => x"030a2808",
			6464 => x"0507f404",
			6465 => x"00006521",
			6466 => x"ff186521",
			6467 => x"05086a08",
			6468 => x"00039e04",
			6469 => x"00a66521",
			6470 => x"00006521",
			6471 => x"00006521",
			6472 => x"00039a40",
			6473 => x"0c05d50c",
			6474 => x"07064104",
			6475 => x"fe5065a5",
			6476 => x"06013904",
			6477 => x"000065a5",
			6478 => x"003865a5",
			6479 => x"0a026d30",
			6480 => x"0d089a1c",
			6481 => x"0003530c",
			6482 => x"0e098708",
			6483 => x"040a0104",
			6484 => x"00ce65a5",
			6485 => x"fea865a5",
			6486 => x"01e665a5",
			6487 => x"0d084a08",
			6488 => x"0f0a0304",
			6489 => x"fdc165a5",
			6490 => x"ff7065a5",
			6491 => x"0e0a1b04",
			6492 => x"00a165a5",
			6493 => x"01fa65a5",
			6494 => x"040a2808",
			6495 => x"07068604",
			6496 => x"000065a5",
			6497 => x"018265a5",
			6498 => x"07072508",
			6499 => x"0802eb04",
			6500 => x"fe2865a5",
			6501 => x"000065a5",
			6502 => x"009c65a5",
			6503 => x"043b65a5",
			6504 => x"fe6865a5",
			6505 => x"0c05f32c",
			6506 => x"0003351c",
			6507 => x"0f094d18",
			6508 => x"0c05d708",
			6509 => x"07064304",
			6510 => x"ff6766b9",
			6511 => x"000066b9",
			6512 => x"0409870c",
			6513 => x"03094f08",
			6514 => x"07061304",
			6515 => x"000066b9",
			6516 => x"004466b9",
			6517 => x"000066b9",
			6518 => x"000066b9",
			6519 => x"00dd66b9",
			6520 => x"07066d0c",
			6521 => x"040a0104",
			6522 => x"000066b9",
			6523 => x"0b06ef04",
			6524 => x"fe7666b9",
			6525 => x"000066b9",
			6526 => x"000066b9",
			6527 => x"0c06133c",
			6528 => x"0d08592c",
			6529 => x"040a491c",
			6530 => x"06014510",
			6531 => x"04091d08",
			6532 => x"06013504",
			6533 => x"000066b9",
			6534 => x"008766b9",
			6535 => x"0f090504",
			6536 => x"000066b9",
			6537 => x"ff4e66b9",
			6538 => x"00035308",
			6539 => x"03093704",
			6540 => x"000066b9",
			6541 => x"014166b9",
			6542 => x"000066b9",
			6543 => x"0309ef08",
			6544 => x"0b06bf04",
			6545 => x"000066b9",
			6546 => x"ff0f66b9",
			6547 => x"020a2d04",
			6548 => x"00ed66b9",
			6549 => x"000066b9",
			6550 => x"02092008",
			6551 => x"0b070104",
			6552 => x"ffcf66b9",
			6553 => x"009d66b9",
			6554 => x"06016704",
			6555 => x"fef266b9",
			6556 => x"000066b9",
			6557 => x"02090008",
			6558 => x"0d085704",
			6559 => x"000066b9",
			6560 => x"ffcc66b9",
			6561 => x"0c064d10",
			6562 => x"00039a0c",
			6563 => x"0507c704",
			6564 => x"000066b9",
			6565 => x"0d08b304",
			6566 => x"012b66b9",
			6567 => x"000066b9",
			6568 => x"000066b9",
			6569 => x"0802b708",
			6570 => x"0b072004",
			6571 => x"000066b9",
			6572 => x"00b166b9",
			6573 => x"ffbf66b9",
			6574 => x"09017a10",
			6575 => x"0a01790c",
			6576 => x"02066104",
			6577 => x"febc678d",
			6578 => x"0600f704",
			6579 => x"01f5678d",
			6580 => x"0000678d",
			6581 => x"fe63678d",
			6582 => x"0d08b344",
			6583 => x"07064024",
			6584 => x"02092e0c",
			6585 => x"0507ab04",
			6586 => x"ff15678d",
			6587 => x"0507e704",
			6588 => x"0196678d",
			6589 => x"0049678d",
			6590 => x"0c05f60c",
			6591 => x"0a021d04",
			6592 => x"fc61678d",
			6593 => x"0a023004",
			6594 => x"00c3678d",
			6595 => x"fe10678d",
			6596 => x"0d082504",
			6597 => x"fe61678d",
			6598 => x"040a9504",
			6599 => x"0177678d",
			6600 => x"0000678d",
			6601 => x"0a02751c",
			6602 => x"0e0a1b10",
			6603 => x"08025a08",
			6604 => x"04091d04",
			6605 => x"01a5678d",
			6606 => x"febb678d",
			6607 => x"01013904",
			6608 => x"0138678d",
			6609 => x"ffdd678d",
			6610 => x"0e0a6308",
			6611 => x"040aed04",
			6612 => x"026b678d",
			6613 => x"0000678d",
			6614 => x"05d6678d",
			6615 => x"fe8b678d",
			6616 => x"0901c314",
			6617 => x"0c063a04",
			6618 => x"ff4a678d",
			6619 => x"0706cb08",
			6620 => x"0b076304",
			6621 => x"01d1678d",
			6622 => x"0000678d",
			6623 => x"0c06a704",
			6624 => x"ff8b678d",
			6625 => x"0000678d",
			6626 => x"fe72678d",
			6627 => x"0c05d810",
			6628 => x"0003460c",
			6629 => x"0e093308",
			6630 => x"07064304",
			6631 => x"ff406881",
			6632 => x"00006881",
			6633 => x"00616881",
			6634 => x"fe7d6881",
			6635 => x"0901c344",
			6636 => x"02092024",
			6637 => x"0d081708",
			6638 => x"0002e604",
			6639 => x"00006881",
			6640 => x"ff406881",
			6641 => x"0002dd10",
			6642 => x"03092e08",
			6643 => x"0a01df04",
			6644 => x"00006881",
			6645 => x"00d06881",
			6646 => x"0100ed04",
			6647 => x"ff1f6881",
			6648 => x"00006881",
			6649 => x"0a01e904",
			6650 => x"00006881",
			6651 => x"03097804",
			6652 => x"01526881",
			6653 => x"00006881",
			6654 => x"0c063010",
			6655 => x"0c05f404",
			6656 => x"00006881",
			6657 => x"0b06cc04",
			6658 => x"00006881",
			6659 => x"0d083e04",
			6660 => x"00006881",
			6661 => x"ff226881",
			6662 => x"0a020804",
			6663 => x"01056881",
			6664 => x"0100f304",
			6665 => x"ff336881",
			6666 => x"020a2d04",
			6667 => x"00ce6881",
			6668 => x"00006881",
			6669 => x"040a3a0c",
			6670 => x"03094f04",
			6671 => x"ffbe6881",
			6672 => x"01013504",
			6673 => x"01586881",
			6674 => x"00006881",
			6675 => x"0209e808",
			6676 => x"0b06cf04",
			6677 => x"00006881",
			6678 => x"febc6881",
			6679 => x"00037808",
			6680 => x"01014b04",
			6681 => x"012f6881",
			6682 => x"00006881",
			6683 => x"0e0a1b04",
			6684 => x"ff0d6881",
			6685 => x"0f0ab204",
			6686 => x"00f26881",
			6687 => x"00006881",
			6688 => x"0901760c",
			6689 => x"0a017908",
			6690 => x"0406a304",
			6691 => x"0000694d",
			6692 => x"0021694d",
			6693 => x"fe6c694d",
			6694 => x"04091d0c",
			6695 => x"03092e08",
			6696 => x"09017a04",
			6697 => x"0000694d",
			6698 => x"01c1694d",
			6699 => x"ffa0694d",
			6700 => x"07063f28",
			6701 => x"0309781c",
			6702 => x"04098710",
			6703 => x"01011108",
			6704 => x"09019604",
			6705 => x"0000694d",
			6706 => x"009d694d",
			6707 => x"07062904",
			6708 => x"0000694d",
			6709 => x"ff66694d",
			6710 => x"07062b08",
			6711 => x"07062604",
			6712 => x"ffbe694d",
			6713 => x"0000694d",
			6714 => x"fda1694d",
			6715 => x"040a5b04",
			6716 => x"0118694d",
			6717 => x"0b06e004",
			6718 => x"feab694d",
			6719 => x"0000694d",
			6720 => x"08025a0c",
			6721 => x"0f092a08",
			6722 => x"0a01ec04",
			6723 => x"fe39694d",
			6724 => x"0000694d",
			6725 => x"007e694d",
			6726 => x"0209280c",
			6727 => x"0b071e08",
			6728 => x"03090704",
			6729 => x"0000694d",
			6730 => x"0172694d",
			6731 => x"0000694d",
			6732 => x"0e093308",
			6733 => x"0b071004",
			6734 => x"fea7694d",
			6735 => x"000c694d",
			6736 => x"02099504",
			6737 => x"00ff694d",
			6738 => x"fff5694d",
			6739 => x"0c05d808",
			6740 => x"00034604",
			6741 => x"00006a21",
			6742 => x"ff0c6a21",
			6743 => x"0c061a34",
			6744 => x"0b071e2c",
			6745 => x"07063f18",
			6746 => x"07062c0c",
			6747 => x"00035308",
			6748 => x"07061304",
			6749 => x"00006a21",
			6750 => x"00a36a21",
			6751 => x"00006a21",
			6752 => x"0309a308",
			6753 => x"0409a004",
			6754 => x"00006a21",
			6755 => x"ff426a21",
			6756 => x"00006a21",
			6757 => x"00038910",
			6758 => x"0100ef08",
			6759 => x"07066c04",
			6760 => x"002c6a21",
			6761 => x"00006a21",
			6762 => x"0b06be04",
			6763 => x"00006a21",
			6764 => x"011f6a21",
			6765 => x"00006a21",
			6766 => x"09019c04",
			6767 => x"ffa36a21",
			6768 => x"00006a21",
			6769 => x"0b070e0c",
			6770 => x"06018d08",
			6771 => x"0c063204",
			6772 => x"ff3f6a21",
			6773 => x"00006a21",
			6774 => x"00006a21",
			6775 => x"0d08b310",
			6776 => x"07066e04",
			6777 => x"00006a21",
			6778 => x"0c065008",
			6779 => x"0003aa04",
			6780 => x"00d16a21",
			6781 => x"00006a21",
			6782 => x"00006a21",
			6783 => x"0706b708",
			6784 => x"09022104",
			6785 => x"ff886a21",
			6786 => x"00006a21",
			6787 => x"01012308",
			6788 => x"0b079304",
			6789 => x"003c6a21",
			6790 => x"00006a21",
			6791 => x"00006a21",
			6792 => x"00038970",
			6793 => x"0c05f53c",
			6794 => x"00034b28",
			6795 => x"09018310",
			6796 => x"0c05f204",
			6797 => x"fe6e6b2d",
			6798 => x"0c05f304",
			6799 => x"01496b2d",
			6800 => x"0c05f404",
			6801 => x"00006b2d",
			6802 => x"fe076b2d",
			6803 => x"0d084b10",
			6804 => x"0d080b08",
			6805 => x"00030c04",
			6806 => x"00d06b2d",
			6807 => x"fece6b2d",
			6808 => x"01012604",
			6809 => x"01d16b2d",
			6810 => x"00bc6b2d",
			6811 => x"0409a004",
			6812 => x"01266b2d",
			6813 => x"febd6b2d",
			6814 => x"0601770c",
			6815 => x"0802b308",
			6816 => x"0f097d04",
			6817 => x"ff766b2d",
			6818 => x"fbca6b2d",
			6819 => x"fe636b2d",
			6820 => x"0309c004",
			6821 => x"febb6b2d",
			6822 => x"01126b2d",
			6823 => x"05084d24",
			6824 => x"0100e808",
			6825 => x"09017a04",
			6826 => x"fe806b2d",
			6827 => x"fff66b2d",
			6828 => x"0c061610",
			6829 => x"0100f108",
			6830 => x"03097804",
			6831 => x"01056b2d",
			6832 => x"fe096b2d",
			6833 => x"040a4904",
			6834 => x"01626b2d",
			6835 => x"001d6b2d",
			6836 => x"0f08f904",
			6837 => x"fede6b2d",
			6838 => x"05082e04",
			6839 => x"021f6b2d",
			6840 => x"00da6b2d",
			6841 => x"040a2804",
			6842 => x"015a6b2d",
			6843 => x"0c066a04",
			6844 => x"fd716b2d",
			6845 => x"030a7804",
			6846 => x"013c6b2d",
			6847 => x"fece6b2d",
			6848 => x"00039514",
			6849 => x"00039104",
			6850 => x"feec6b2d",
			6851 => x"0101570c",
			6852 => x"09021504",
			6853 => x"ffac6b2d",
			6854 => x"01015104",
			6855 => x"00ea6b2d",
			6856 => x"00006b2d",
			6857 => x"ff6d6b2d",
			6858 => x"fe676b2d",
			6859 => x"0003897c",
			6860 => x"0c05f534",
			6861 => x"00034b24",
			6862 => x"0901830c",
			6863 => x"0600ef08",
			6864 => x"0c054604",
			6865 => x"ff026c49",
			6866 => x"00f36c49",
			6867 => x"fe7d6c49",
			6868 => x"0d084b10",
			6869 => x"0d080b08",
			6870 => x"0208d004",
			6871 => x"00de6c49",
			6872 => x"fec16c49",
			6873 => x"0802aa04",
			6874 => x"014d6c49",
			6875 => x"025a6c49",
			6876 => x"07065a04",
			6877 => x"fe896c49",
			6878 => x"01316c49",
			6879 => x"0802b308",
			6880 => x"0f098b04",
			6881 => x"ff5e6c49",
			6882 => x"fad76c49",
			6883 => x"0b06dc04",
			6884 => x"fe4f6c49",
			6885 => x"00a76c49",
			6886 => x"05082124",
			6887 => x"05081f1c",
			6888 => x"09017d0c",
			6889 => x"0002e608",
			6890 => x"0b06ff04",
			6891 => x"feab6c49",
			6892 => x"fc596c49",
			6893 => x"00586c49",
			6894 => x"0c061008",
			6895 => x"00035304",
			6896 => x"01076c49",
			6897 => x"feea6c49",
			6898 => x"06013d04",
			6899 => x"ffa66c49",
			6900 => x"01966c49",
			6901 => x"0100ef04",
			6902 => x"03826c49",
			6903 => x"01996c49",
			6904 => x"07067010",
			6905 => x"0100f108",
			6906 => x"08025f04",
			6907 => x"00566c49",
			6908 => x"fd136c49",
			6909 => x"030a0104",
			6910 => x"01656c49",
			6911 => x"00006c49",
			6912 => x"0209c908",
			6913 => x"0b071004",
			6914 => x"00496c49",
			6915 => x"01a96c49",
			6916 => x"01011904",
			6917 => x"fe496c49",
			6918 => x"01014304",
			6919 => x"019b6c49",
			6920 => x"feeb6c49",
			6921 => x"00039510",
			6922 => x"00039204",
			6923 => x"ff106c49",
			6924 => x"01015708",
			6925 => x"01014d04",
			6926 => x"00006c49",
			6927 => x"00776c49",
			6928 => x"00006c49",
			6929 => x"fe676c49",
			6930 => x"0c05d508",
			6931 => x"07064104",
			6932 => x"fe6b6cf5",
			6933 => x"00006cf5",
			6934 => x"040af74c",
			6935 => x"0b06ef2c",
			6936 => x"0101391c",
			6937 => x"0d084b10",
			6938 => x"03098708",
			6939 => x"01012404",
			6940 => x"00a16cf5",
			6941 => x"fdcf6cf5",
			6942 => x"00035304",
			6943 => x"01ab6cf5",
			6944 => x"00006cf5",
			6945 => x"08029108",
			6946 => x"0c05f404",
			6947 => x"00006cf5",
			6948 => x"fe5e6cf5",
			6949 => x"01586cf5",
			6950 => x"0309d804",
			6951 => x"fd5b6cf5",
			6952 => x"00037004",
			6953 => x"01386cf5",
			6954 => x"0c05f404",
			6955 => x"00006cf5",
			6956 => x"fece6cf5",
			6957 => x"02090008",
			6958 => x"0c061204",
			6959 => x"00006cf5",
			6960 => x"fe946cf5",
			6961 => x"03097808",
			6962 => x"0c060f04",
			6963 => x"00006cf5",
			6964 => x"01ce6cf5",
			6965 => x"0100ff08",
			6966 => x"0c061304",
			6967 => x"fe886cf5",
			6968 => x"005f6cf5",
			6969 => x"0d08b304",
			6970 => x"018e6cf5",
			6971 => x"ffac6cf5",
			6972 => x"fea96cf5",
			6973 => x"00039a6c",
			6974 => x"07067048",
			6975 => x"07066e38",
			6976 => x"07064018",
			6977 => x"07062c0c",
			6978 => x"07061304",
			6979 => x"ff046dd1",
			6980 => x"0d083204",
			6981 => x"00b76dd1",
			6982 => x"00006dd1",
			6983 => x"0208e404",
			6984 => x"00006dd1",
			6985 => x"0b06bc04",
			6986 => x"00006dd1",
			6987 => x"fe8f6dd1",
			6988 => x"0507c710",
			6989 => x"0b06bc08",
			6990 => x"0b06af04",
			6991 => x"00006dd1",
			6992 => x"01846dd1",
			6993 => x"01010f04",
			6994 => x"00206dd1",
			6995 => x"fdf36dd1",
			6996 => x"01013d08",
			6997 => x"08026404",
			6998 => x"00006dd1",
			6999 => x"00fd6dd1",
			7000 => x"0b06de04",
			7001 => x"fe8b6dd1",
			7002 => x"003d6dd1",
			7003 => x"06014104",
			7004 => x"00006dd1",
			7005 => x"0d084b04",
			7006 => x"00006dd1",
			7007 => x"06016704",
			7008 => x"fe796dd1",
			7009 => x"00006dd1",
			7010 => x"0d088208",
			7011 => x"08025304",
			7012 => x"00006dd1",
			7013 => x"01686dd1",
			7014 => x"0b072008",
			7015 => x"05083004",
			7016 => x"00096dd1",
			7017 => x"fe386dd1",
			7018 => x"0d08b308",
			7019 => x"0d088d04",
			7020 => x"00006dd1",
			7021 => x"01576dd1",
			7022 => x"07072508",
			7023 => x"06019704",
			7024 => x"ff466dd1",
			7025 => x"00006dd1",
			7026 => x"00006dd1",
			7027 => x"fe766dd1",
			7028 => x"0c05d508",
			7029 => x"07064104",
			7030 => x"fec56ed5",
			7031 => x"00006ed5",
			7032 => x"02099548",
			7033 => x"0a01f220",
			7034 => x"0507d708",
			7035 => x"0c05d904",
			7036 => x"00006ed5",
			7037 => x"00736ed5",
			7038 => x"0209110c",
			7039 => x"08025f08",
			7040 => x"0208e204",
			7041 => x"00006ed5",
			7042 => x"fee96ed5",
			7043 => x"00006ed5",
			7044 => x"02092808",
			7045 => x"0100eb04",
			7046 => x"00006ed5",
			7047 => x"00e86ed5",
			7048 => x"ff3f6ed5",
			7049 => x"0507ca18",
			7050 => x"0507ac0c",
			7051 => x"07063f04",
			7052 => x"00006ed5",
			7053 => x"00034604",
			7054 => x"00b56ed5",
			7055 => x"00006ed5",
			7056 => x"0901cc08",
			7057 => x"0b06ce04",
			7058 => x"00456ed5",
			7059 => x"00006ed5",
			7060 => x"ff0b6ed5",
			7061 => x"0309c008",
			7062 => x"0100ed04",
			7063 => x"00006ed5",
			7064 => x"015b6ed5",
			7065 => x"02097b04",
			7066 => x"ffa56ed5",
			7067 => x"00006ed5",
			7068 => x"0e098710",
			7069 => x"06015e04",
			7070 => x"00006ed5",
			7071 => x"07062c04",
			7072 => x"00006ed5",
			7073 => x"0f09a304",
			7074 => x"00006ed5",
			7075 => x"feb06ed5",
			7076 => x"0209c104",
			7077 => x"00f16ed5",
			7078 => x"0e0a1b10",
			7079 => x"0b074408",
			7080 => x"07065804",
			7081 => x"00006ed5",
			7082 => x"ff076ed5",
			7083 => x"020a3a04",
			7084 => x"00636ed5",
			7085 => x"00006ed5",
			7086 => x"06019108",
			7087 => x"00037804",
			7088 => x"00006ed5",
			7089 => x"ffe36ed5",
			7090 => x"00039a04",
			7091 => x"01036ed5",
			7092 => x"00006ed5",
			7093 => x"00039a7c",
			7094 => x"0b06ef40",
			7095 => x"04091d14",
			7096 => x"09017a0c",
			7097 => x"0801cb08",
			7098 => x"0b05e504",
			7099 => x"fff56fd1",
			7100 => x"01026fd1",
			7101 => x"fee76fd1",
			7102 => x"0507e604",
			7103 => x"01906fd1",
			7104 => x"00006fd1",
			7105 => x"0e09871c",
			7106 => x"02099510",
			7107 => x"0e094008",
			7108 => x"00032404",
			7109 => x"ffdf6fd1",
			7110 => x"fdb76fd1",
			7111 => x"0c05f304",
			7112 => x"ffe66fd1",
			7113 => x"01a26fd1",
			7114 => x"07065908",
			7115 => x"0c05da04",
			7116 => x"00006fd1",
			7117 => x"fe356fd1",
			7118 => x"fbe46fd1",
			7119 => x"00037008",
			7120 => x"0901d904",
			7121 => x"ff856fd1",
			7122 => x"01a86fd1",
			7123 => x"020a4604",
			7124 => x"fe8a6fd1",
			7125 => x"00006fd1",
			7126 => x"0508211c",
			7127 => x"08025304",
			7128 => x"feea6fd1",
			7129 => x"0b071e10",
			7130 => x"0c060f08",
			7131 => x"0c05f504",
			7132 => x"00836fd1",
			7133 => x"ffb26fd1",
			7134 => x"0c063a04",
			7135 => x"01e56fd1",
			7136 => x"00006fd1",
			7137 => x"0f095604",
			7138 => x"ff436fd1",
			7139 => x"00996fd1",
			7140 => x"0802e818",
			7141 => x"0c06300c",
			7142 => x"05083e08",
			7143 => x"09018704",
			7144 => x"ff1b6fd1",
			7145 => x"01096fd1",
			7146 => x"fe526fd1",
			7147 => x"00037008",
			7148 => x"0f094d04",
			7149 => x"ff5c6fd1",
			7150 => x"013d6fd1",
			7151 => x"fef86fd1",
			7152 => x"0b074404",
			7153 => x"02226fd1",
			7154 => x"00006fd1",
			7155 => x"fe6c6fd1",
			7156 => x"00039a78",
			7157 => x"07064024",
			7158 => x"0409720c",
			7159 => x"0100ef08",
			7160 => x"0600ef04",
			7161 => x"000070c5",
			7162 => x"ff9e70c5",
			7163 => x"00c770c5",
			7164 => x"06016b08",
			7165 => x"0a020004",
			7166 => x"000070c5",
			7167 => x"fea670c5",
			7168 => x"0a02530c",
			7169 => x"0b06bc04",
			7170 => x"000070c5",
			7171 => x"0e094004",
			7172 => x"000070c5",
			7173 => x"00fe70c5",
			7174 => x"feee70c5",
			7175 => x"0706581c",
			7176 => x"0e098714",
			7177 => x"0f09b110",
			7178 => x"08024e08",
			7179 => x"0507ad04",
			7180 => x"000070c5",
			7181 => x"ff8f70c5",
			7182 => x"0b06be04",
			7183 => x"000070c5",
			7184 => x"013670c5",
			7185 => x"ff4470c5",
			7186 => x"0a025c04",
			7187 => x"01b470c5",
			7188 => x"000070c5",
			7189 => x"0f096820",
			7190 => x"07066c10",
			7191 => x"06013d08",
			7192 => x"0507d804",
			7193 => x"000070c5",
			7194 => x"ffc570c5",
			7195 => x"0d081804",
			7196 => x"000070c5",
			7197 => x"017170c5",
			7198 => x"0002ee08",
			7199 => x"03094f04",
			7200 => x"017970c5",
			7201 => x"fed170c5",
			7202 => x"0e090704",
			7203 => x"000070c5",
			7204 => x"015e70c5",
			7205 => x"0e09c10c",
			7206 => x"00034b08",
			7207 => x"06016204",
			7208 => x"feda70c5",
			7209 => x"015570c5",
			7210 => x"fe0a70c5",
			7211 => x"0802ee08",
			7212 => x"01014704",
			7213 => x"008b70c5",
			7214 => x"feb770c5",
			7215 => x"018370c5",
			7216 => x"fe7370c5",
			7217 => x"00039a80",
			7218 => x"0100f13c",
			7219 => x"0309782c",
			7220 => x"0209001c",
			7221 => x"04091d0c",
			7222 => x"06013d08",
			7223 => x"0600ef04",
			7224 => x"007e71cb",
			7225 => x"ff2d71cb",
			7226 => x"01e271cb",
			7227 => x"06014108",
			7228 => x"08025a04",
			7229 => x"fe1571cb",
			7230 => x"ffca71cb",
			7231 => x"03091a04",
			7232 => x"ffad71cb",
			7233 => x"007671cb",
			7234 => x"0b07010c",
			7235 => x"06014104",
			7236 => x"fe9371cb",
			7237 => x"0100e904",
			7238 => x"ff6d71cb",
			7239 => x"01d871cb",
			7240 => x"024c71cb",
			7241 => x"09017d04",
			7242 => x"fdfc71cb",
			7243 => x"03098704",
			7244 => x"010071cb",
			7245 => x"0b071004",
			7246 => x"fe7f71cb",
			7247 => x"00f071cb",
			7248 => x"07065b20",
			7249 => x"0100ff04",
			7250 => x"016871cb",
			7251 => x"0901b80c",
			7252 => x"02093a08",
			7253 => x"0a01fa04",
			7254 => x"feb071cb",
			7255 => x"012c71cb",
			7256 => x"fdeb71cb",
			7257 => x"0e092408",
			7258 => x"04098704",
			7259 => x"006571cb",
			7260 => x"fe8d71cb",
			7261 => x"040a3a04",
			7262 => x"014771cb",
			7263 => x"ffaf71cb",
			7264 => x"05086a18",
			7265 => x"09018708",
			7266 => x"04098704",
			7267 => x"008471cb",
			7268 => x"ffcc71cb",
			7269 => x"0b06dc08",
			7270 => x"040a3a04",
			7271 => x"00f571cb",
			7272 => x"ff9f71cb",
			7273 => x"0706a104",
			7274 => x"01a671cb",
			7275 => x"003771cb",
			7276 => x"07072508",
			7277 => x"05088604",
			7278 => x"000071cb",
			7279 => x"febd71cb",
			7280 => x"003471cb",
			7281 => x"fe6a71cb",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(2358, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(4838, initial_addr_3'length));
	end generate gen_rom_2;

	gen_rom_3: if SELECT_ROM = 3 generate
		bank <= (
			0 => x"00000005",
			1 => x"00000009",
			2 => x"0000000d",
			3 => x"00000011",
			4 => x"00000015",
			5 => x"00000019",
			6 => x"0000001d",
			7 => x"00000021",
			8 => x"00000025",
			9 => x"00000029",
			10 => x"0000002d",
			11 => x"00000031",
			12 => x"00000035",
			13 => x"00000039",
			14 => x"0000003d",
			15 => x"00000041",
			16 => x"00000045",
			17 => x"00000049",
			18 => x"0000004d",
			19 => x"00000051",
			20 => x"00000055",
			21 => x"00000059",
			22 => x"00021b04",
			23 => x"00000065",
			24 => x"ffeb0065",
			25 => x"0c052504",
			26 => x"fff20071",
			27 => x"00000071",
			28 => x"02061a04",
			29 => x"0025007d",
			30 => x"0000007d",
			31 => x"0405d204",
			32 => x"00000089",
			33 => x"fffd0089",
			34 => x"0f060a04",
			35 => x"00000095",
			36 => x"ffea0095",
			37 => x"0406ea04",
			38 => x"000b00a1",
			39 => x"000000a1",
			40 => x"02061a04",
			41 => x"002e00ad",
			42 => x"000000ad",
			43 => x"0406a304",
			44 => x"00bd00c1",
			45 => x"09011304",
			46 => x"ffc600c1",
			47 => x"000000c1",
			48 => x"0900f304",
			49 => x"ffe700d5",
			50 => x"09017404",
			51 => x"001a00d5",
			52 => x"000000d5",
			53 => x"00021b04",
			54 => x"003400e9",
			55 => x"0f08b104",
			56 => x"fff600e9",
			57 => x"000000e9",
			58 => x"0f062f08",
			59 => x"0002d504",
			60 => x"002200fd",
			61 => x"000000fd",
			62 => x"000000fd",
			63 => x"00028d08",
			64 => x"0e070104",
			65 => x"01c40111",
			66 => x"d5d10111",
			67 => x"c3d10111",
			68 => x"0a016608",
			69 => x"0c054304",
			70 => x"0136012d",
			71 => x"0000012d",
			72 => x"0900f704",
			73 => x"fff3012d",
			74 => x"0000012d",
			75 => x"02061a08",
			76 => x"0600d704",
			77 => x"00000149",
			78 => x"00aa0149",
			79 => x"01009d04",
			80 => x"ffc50149",
			81 => x"00000149",
			82 => x"02061a08",
			83 => x"0c04d004",
			84 => x"00000165",
			85 => x"00550165",
			86 => x"07069b04",
			87 => x"ffaa0165",
			88 => x"00000165",
			89 => x"0900f70c",
			90 => x"02059a04",
			91 => x"00000181",
			92 => x"01009704",
			93 => x"ff850181",
			94 => x"00000181",
			95 => x"00000181",
			96 => x"01009204",
			97 => x"0000019d",
			98 => x"0e073b08",
			99 => x"08024704",
			100 => x"0064019d",
			101 => x"0000019d",
			102 => x"0000019d",
			103 => x"0900f30c",
			104 => x"0e059d04",
			105 => x"000001b9",
			106 => x"01009704",
			107 => x"ffdd01b9",
			108 => x"000001b9",
			109 => x"000001b9",
			110 => x"0406a304",
			111 => x"000001d5",
			112 => x"00021b04",
			113 => x"000001d5",
			114 => x"0f067a04",
			115 => x"000001d5",
			116 => x"fffa01d5",
			117 => x"00021b08",
			118 => x"0c054304",
			119 => x"00bb01f9",
			120 => x"000001f9",
			121 => x"0100a108",
			122 => x"0c056204",
			123 => x"ff8001f9",
			124 => x"000001f9",
			125 => x"000001f9",
			126 => x"02077710",
			127 => x"0900f308",
			128 => x"0e059d04",
			129 => x"0000021d",
			130 => x"ffae021d",
			131 => x"0f06de04",
			132 => x"00e6021d",
			133 => x"0000021d",
			134 => x"ff0e021d",
			135 => x"0c04d40c",
			136 => x"0405d204",
			137 => x"00000249",
			138 => x"07051f04",
			139 => x"ff4e0249",
			140 => x"00000249",
			141 => x"0b059708",
			142 => x"0002d504",
			143 => x"006e0249",
			144 => x"00000249",
			145 => x"00000249",
			146 => x"0900ef04",
			147 => x"0000026d",
			148 => x"0901740c",
			149 => x"07053104",
			150 => x"0000026d",
			151 => x"0308e704",
			152 => x"0028026d",
			153 => x"0000026d",
			154 => x"0000026d",
			155 => x"0900f304",
			156 => x"00000291",
			157 => x"0901740c",
			158 => x"0d083808",
			159 => x"0d064704",
			160 => x"00000291",
			161 => x"00220291",
			162 => x"00000291",
			163 => x"00000291",
			164 => x"0406ea10",
			165 => x"0900f70c",
			166 => x"0305b904",
			167 => x"000002bd",
			168 => x"07051a04",
			169 => x"000002bd",
			170 => x"ffd202bd",
			171 => x"006202bd",
			172 => x"09012004",
			173 => x"ff1e02bd",
			174 => x"000002bd",
			175 => x"01009210",
			176 => x"0f05ad04",
			177 => x"000002e9",
			178 => x"0b058508",
			179 => x"07054904",
			180 => x"ff7202e9",
			181 => x"000002e9",
			182 => x"000002e9",
			183 => x"0f06de04",
			184 => x"012f02e9",
			185 => x"000002e9",
			186 => x"02061a08",
			187 => x"01009204",
			188 => x"00000315",
			189 => x"00b10315",
			190 => x"0901200c",
			191 => x"0100ad08",
			192 => x"04065904",
			193 => x"00000315",
			194 => x"ffae0315",
			195 => x"00000315",
			196 => x"00000315",
			197 => x"0c052808",
			198 => x"0900fb04",
			199 => x"ffd00341",
			200 => x"00000341",
			201 => x"0901740c",
			202 => x"0c061508",
			203 => x"0900e004",
			204 => x"00000341",
			205 => x"00340341",
			206 => x"00000341",
			207 => x"00000341",
			208 => x"02077714",
			209 => x"0900f30c",
			210 => x"0e059d04",
			211 => x"0000036d",
			212 => x"07051a04",
			213 => x"0000036d",
			214 => x"ff95036d",
			215 => x"0f06de04",
			216 => x"00f7036d",
			217 => x"0000036d",
			218 => x"ff04036d",
			219 => x"0900fb0c",
			220 => x"0e059d04",
			221 => x"000003a1",
			222 => x"01009b04",
			223 => x"ffca03a1",
			224 => x"000003a1",
			225 => x"0100e50c",
			226 => x"0e087f08",
			227 => x"07051f04",
			228 => x"000003a1",
			229 => x"002f03a1",
			230 => x"000003a1",
			231 => x"000003a1",
			232 => x"0406ea14",
			233 => x"0100920c",
			234 => x"0305b904",
			235 => x"000003dd",
			236 => x"07051a04",
			237 => x"000003dd",
			238 => x"ffd503dd",
			239 => x"0600ea04",
			240 => x"000003dd",
			241 => x"005903dd",
			242 => x"07058c08",
			243 => x"0c056404",
			244 => x"ff2d03dd",
			245 => x"000003dd",
			246 => x"000003dd",
			247 => x"0900f310",
			248 => x"0405d204",
			249 => x"00000419",
			250 => x"01009708",
			251 => x"07055d04",
			252 => x"ff9e0419",
			253 => x"00000419",
			254 => x"00000419",
			255 => x"0a01df0c",
			256 => x"0e087f08",
			257 => x"0100a104",
			258 => x"00000419",
			259 => x"00660419",
			260 => x"00000419",
			261 => x"00000419",
			262 => x"08024718",
			263 => x"0900f30c",
			264 => x"0f060a08",
			265 => x"07050104",
			266 => x"0000044d",
			267 => x"0080044d",
			268 => x"ffb5044d",
			269 => x"07054904",
			270 => x"0000044d",
			271 => x"0308e704",
			272 => x"00e1044d",
			273 => x"0000044d",
			274 => x"ff42044d",
			275 => x"0b053508",
			276 => x"0405d204",
			277 => x"00000481",
			278 => x"ff980481",
			279 => x"0408ea10",
			280 => x"0900f304",
			281 => x"00000481",
			282 => x"0e087f08",
			283 => x"0100e504",
			284 => x"004c0481",
			285 => x"00000481",
			286 => x"00000481",
			287 => x"00000481",
			288 => x"0900f308",
			289 => x"0c054604",
			290 => x"ffea04b5",
			291 => x"000004b5",
			292 => x"09017410",
			293 => x"0507d70c",
			294 => x"07051f04",
			295 => x"000004b5",
			296 => x"0c061504",
			297 => x"002704b5",
			298 => x"000004b5",
			299 => x"000004b5",
			300 => x"000004b5",
			301 => x"00021b04",
			302 => x"007804e1",
			303 => x"0100a104",
			304 => x"ff5d04e1",
			305 => x"02088b0c",
			306 => x"06013808",
			307 => x"0507c904",
			308 => x"003604e1",
			309 => x"000004e1",
			310 => x"000004e1",
			311 => x"000004e1",
			312 => x"00028d14",
			313 => x"0c04d004",
			314 => x"ffc2051d",
			315 => x"0f076d0c",
			316 => x"01009b08",
			317 => x"03064804",
			318 => x"01b2051d",
			319 => x"fdee051d",
			320 => x"01c1051d",
			321 => x"ff8c051d",
			322 => x"0408ab08",
			323 => x"0a01cc04",
			324 => x"fea4051d",
			325 => x"0349051d",
			326 => x"fe65051d",
			327 => x"0c05280c",
			328 => x"0a014504",
			329 => x"00000559",
			330 => x"0100a104",
			331 => x"ffaa0559",
			332 => x"00000559",
			333 => x"01009304",
			334 => x"00000559",
			335 => x"02088b0c",
			336 => x"0100e508",
			337 => x"0308e704",
			338 => x"00830559",
			339 => x"00000559",
			340 => x"00000559",
			341 => x"00000559",
			342 => x"00028d18",
			343 => x"0f060a08",
			344 => x"0b053504",
			345 => x"0031058d",
			346 => x"019a058d",
			347 => x"0900fb04",
			348 => x"fd9a058d",
			349 => x"0f070104",
			350 => x"019a058d",
			351 => x"09013804",
			352 => x"fe05058d",
			353 => x"0140058d",
			354 => x"fe67058d",
			355 => x"0a01b618",
			356 => x"03076c14",
			357 => x"0c04d008",
			358 => x"0405d204",
			359 => x"028205d1",
			360 => x"ff5b05d1",
			361 => x"0f070108",
			362 => x"02066104",
			363 => x"028705d1",
			364 => x"024305d1",
			365 => x"009a05d1",
			366 => x"06b005d1",
			367 => x"0408ab08",
			368 => x"04089204",
			369 => x"fe7405d1",
			370 => x"ffd905d1",
			371 => x"fe5f05d1",
			372 => x"0c052810",
			373 => x"02059a04",
			374 => x"00000615",
			375 => x"0900fb08",
			376 => x"0d068504",
			377 => x"ffaf0615",
			378 => x"00000615",
			379 => x"00000615",
			380 => x"0900ef04",
			381 => x"00000615",
			382 => x"02088b0c",
			383 => x"09017608",
			384 => x"0507d704",
			385 => x"00740615",
			386 => x"00000615",
			387 => x"00000615",
			388 => x"00000615",
			389 => x"00028d18",
			390 => x"01007904",
			391 => x"ff320661",
			392 => x"0f07010c",
			393 => x"0c04ed08",
			394 => x"03060904",
			395 => x"01b70661",
			396 => x"ff300661",
			397 => x"01a40661",
			398 => x"0705a104",
			399 => x"fda50661",
			400 => x"01e90661",
			401 => x"0408ea0c",
			402 => x"0a01d704",
			403 => x"fe7e0661",
			404 => x"08024704",
			405 => x"04130661",
			406 => x"ffba0661",
			407 => x"fe650661",
			408 => x"01009b18",
			409 => x"0f060a0c",
			410 => x"0c04cf04",
			411 => x"000006b5",
			412 => x"06011c04",
			413 => x"002906b5",
			414 => x"000006b5",
			415 => x"0c056008",
			416 => x"0600e604",
			417 => x"000006b5",
			418 => x"ff1606b5",
			419 => x"000006b5",
			420 => x"02088b10",
			421 => x"0600f104",
			422 => x"000006b5",
			423 => x"0100e508",
			424 => x"0507d704",
			425 => x"009706b5",
			426 => x"000006b5",
			427 => x"000006b5",
			428 => x"000006b5",
			429 => x"0408ab20",
			430 => x"01009910",
			431 => x"04062708",
			432 => x"0600cd04",
			433 => x"000006f9",
			434 => x"014c06f9",
			435 => x"01009204",
			436 => x"feb906f9",
			437 => x"ffdf06f9",
			438 => x"0f070104",
			439 => x"015d06f9",
			440 => x"0d071604",
			441 => x"ffc106f9",
			442 => x"0f087a04",
			443 => x"009706f9",
			444 => x"000006f9",
			445 => x"fe7206f9",
			446 => x"0b053508",
			447 => x"0405d204",
			448 => x"0000073d",
			449 => x"ff4b073d",
			450 => x"0406a304",
			451 => x"0071073d",
			452 => x"0c06140c",
			453 => x"0c04e904",
			454 => x"0000073d",
			455 => x"0c054804",
			456 => x"ffa6073d",
			457 => x"0000073d",
			458 => x"0c061508",
			459 => x"0b06cf04",
			460 => x"0000073d",
			461 => x"003d073d",
			462 => x"0000073d",
			463 => x"0b053508",
			464 => x"0405d204",
			465 => x"00000789",
			466 => x"ff410789",
			467 => x"0f067a08",
			468 => x"00030204",
			469 => x"00810789",
			470 => x"00000789",
			471 => x"0100a108",
			472 => x"0c056204",
			473 => x"ffa80789",
			474 => x"00000789",
			475 => x"0802470c",
			476 => x"0e087f08",
			477 => x"0801cb04",
			478 => x"00000789",
			479 => x"00560789",
			480 => x"00000789",
			481 => x"00000789",
			482 => x"08024724",
			483 => x"01009b14",
			484 => x"0801a50c",
			485 => x"0e059d04",
			486 => x"007d07d5",
			487 => x"07051b04",
			488 => x"ff9b07d5",
			489 => x"000007d5",
			490 => x"0c050b04",
			491 => x"000007d5",
			492 => x"ff3807d5",
			493 => x"0e087f0c",
			494 => x"0507d708",
			495 => x"02088b04",
			496 => x"009707d5",
			497 => x"000007d5",
			498 => x"000007d5",
			499 => x"000007d5",
			500 => x"fed107d5",
			501 => x"0408ab1c",
			502 => x"01006c04",
			503 => x"fefe0811",
			504 => x"0f060a04",
			505 => x"018d0811",
			506 => x"0705490c",
			507 => x"01009b04",
			508 => x"fe9d0811",
			509 => x"0c051104",
			510 => x"004b0811",
			511 => x"ffbf0811",
			512 => x"0f087a04",
			513 => x"01480811",
			514 => x"00000811",
			515 => x"fe6a0811",
			516 => x"08024724",
			517 => x"01009b10",
			518 => x"00021b0c",
			519 => x"01007904",
			520 => x"0000085d",
			521 => x"01009504",
			522 => x"00f5085d",
			523 => x"0000085d",
			524 => x"ff1a085d",
			525 => x"0f070104",
			526 => x"00f7085d",
			527 => x"0c061404",
			528 => x"ffb9085d",
			529 => x"0002bf04",
			530 => x"0000085d",
			531 => x"0208ab04",
			532 => x"00a4085d",
			533 => x"0000085d",
			534 => x"fe9d085d",
			535 => x"08024728",
			536 => x"0100a614",
			537 => x"0e059d08",
			538 => x"0600e604",
			539 => x"002e08b1",
			540 => x"000008b1",
			541 => x"01009204",
			542 => x"ff4f08b1",
			543 => x"0600f204",
			544 => x"000608b1",
			545 => x"fffe08b1",
			546 => x"0e087f10",
			547 => x"0600f204",
			548 => x"000008b1",
			549 => x"0c052704",
			550 => x"000008b1",
			551 => x"0507c904",
			552 => x"00a808b1",
			553 => x"000008b1",
			554 => x"000008b1",
			555 => x"ff0708b1",
			556 => x"0002cc1c",
			557 => x"0c04d004",
			558 => x"ff8208ed",
			559 => x"0406a304",
			560 => x"010908ed",
			561 => x"0c052a04",
			562 => x"ff8f08ed",
			563 => x"0e087f0c",
			564 => x"09012004",
			565 => x"000008ed",
			566 => x"0308e704",
			567 => x"00e408ed",
			568 => x"000008ed",
			569 => x"000008ed",
			570 => x"fe8908ed",
			571 => x"0002cc24",
			572 => x"0706581c",
			573 => x"02077718",
			574 => x"0900f30c",
			575 => x"04062708",
			576 => x"0c04cf04",
			577 => x"fff70939",
			578 => x"01640939",
			579 => x"fe5a0939",
			580 => x"0f070104",
			581 => x"01850939",
			582 => x"0506e204",
			583 => x"ff630939",
			584 => x"012a0939",
			585 => x"fee50939",
			586 => x"02089004",
			587 => x"03840939",
			588 => x"00000939",
			589 => x"fe6d0939",
			590 => x"0408ab20",
			591 => x"01006f04",
			592 => x"fe00097d",
			593 => x"02076714",
			594 => x"01009210",
			595 => x"0f05d20c",
			596 => x"0e059d04",
			597 => x"01b5097d",
			598 => x"0e05ac04",
			599 => x"0000097d",
			600 => x"013c097d",
			601 => x"fdcb097d",
			602 => x"019c097d",
			603 => x"09016504",
			604 => x"fe8b097d",
			605 => x"0473097d",
			606 => x"fe66097d",
			607 => x"0002cc28",
			608 => x"0c06141c",
			609 => x"02077718",
			610 => x"0900f30c",
			611 => x"04062708",
			612 => x"0c04cf04",
			613 => x"000009d1",
			614 => x"015e09d1",
			615 => x"fe8809d1",
			616 => x"0e06ce04",
			617 => x"018009d1",
			618 => x"0705a204",
			619 => x"feea09d1",
			620 => x"013f09d1",
			621 => x"fef609d1",
			622 => x"0b06cf04",
			623 => x"000009d1",
			624 => x"0507d804",
			625 => x"02f309d1",
			626 => x"000009d1",
			627 => x"fe6e09d1",
			628 => x"0002cc24",
			629 => x"0706581c",
			630 => x"0f077b18",
			631 => x"0c04d008",
			632 => x"0405d204",
			633 => x"00eb0a1d",
			634 => x"feac0a1d",
			635 => x"0c051104",
			636 => x"01700a1d",
			637 => x"0100a108",
			638 => x"03064804",
			639 => x"00c80a1d",
			640 => x"ff110a1d",
			641 => x"015c0a1d",
			642 => x"ff080a1d",
			643 => x"0308e704",
			644 => x"02870a1d",
			645 => x"00000a1d",
			646 => x"fe6f0a1d",
			647 => x"08024724",
			648 => x"01007908",
			649 => x"0f058504",
			650 => x"00000a69",
			651 => x"ff0b0a69",
			652 => x"0b059904",
			653 => x"014b0a69",
			654 => x"0c052a08",
			655 => x"0f067a04",
			656 => x"00000a69",
			657 => x"fef70a69",
			658 => x"0e087f0c",
			659 => x"0100a604",
			660 => x"00000a69",
			661 => x"0600f204",
			662 => x"00000a69",
			663 => x"00ff0a69",
			664 => x"00000a69",
			665 => x"fe860a69",
			666 => x"0002cc2c",
			667 => x"0100a614",
			668 => x"00021b0c",
			669 => x"0c04d004",
			670 => x"ff7d0ac5",
			671 => x"0c054304",
			672 => x"01430ac5",
			673 => x"00000ac5",
			674 => x"0100a104",
			675 => x"fe8b0ac5",
			676 => x"00000ac5",
			677 => x"0600f104",
			678 => x"00000ac5",
			679 => x"02088b10",
			680 => x"0c052704",
			681 => x"00000ac5",
			682 => x"0100e508",
			683 => x"0507c904",
			684 => x"01590ac5",
			685 => x"00000ac5",
			686 => x"00000ac5",
			687 => x"00000ac5",
			688 => x"fe7b0ac5",
			689 => x"0002cc28",
			690 => x"0c04d004",
			691 => x"ffa80b1b",
			692 => x"0f067a0c",
			693 => x"0900f308",
			694 => x"0900ef04",
			695 => x"006e0b1b",
			696 => x"00000b1b",
			697 => x"01320b1b",
			698 => x"0a017908",
			699 => x"0100b404",
			700 => x"ff510b1b",
			701 => x"00000b1b",
			702 => x"0e087f0c",
			703 => x"0c052a04",
			704 => x"00000b1b",
			705 => x"0308e704",
			706 => x"00bc0b1b",
			707 => x"00000b1b",
			708 => x"00000b1b",
			709 => x"fe900b1b",
			710 => x"00000b1d",
			711 => x"00000b21",
			712 => x"00000b25",
			713 => x"00000b29",
			714 => x"00000b2d",
			715 => x"00000b31",
			716 => x"00000b35",
			717 => x"00000b39",
			718 => x"00000b3d",
			719 => x"00000b41",
			720 => x"00000b45",
			721 => x"00000b49",
			722 => x"00000b4d",
			723 => x"00000b51",
			724 => x"00000b55",
			725 => x"00000b59",
			726 => x"00000b5d",
			727 => x"00000b61",
			728 => x"00000b65",
			729 => x"00000b69",
			730 => x"00000b6d",
			731 => x"00000b71",
			732 => x"00021b04",
			733 => x"00000b7d",
			734 => x"fff50b7d",
			735 => x"0c052504",
			736 => x"fff60b89",
			737 => x"00000b89",
			738 => x"02061a04",
			739 => x"00240b95",
			740 => x"00000b95",
			741 => x"0405d204",
			742 => x"00000ba1",
			743 => x"fffe0ba1",
			744 => x"0f060a04",
			745 => x"00000bad",
			746 => x"ffee0bad",
			747 => x"0406ea04",
			748 => x"00080bb9",
			749 => x"00000bb9",
			750 => x"02061a04",
			751 => x"002b0bc5",
			752 => x"00000bc5",
			753 => x"02066104",
			754 => x"00ae0bd9",
			755 => x"09011304",
			756 => x"ffce0bd9",
			757 => x"00000bd9",
			758 => x"0900f304",
			759 => x"ffec0bed",
			760 => x"09017404",
			761 => x"00140bed",
			762 => x"00000bed",
			763 => x"00021b04",
			764 => x"002f0c01",
			765 => x"0f08b104",
			766 => x"fffc0c01",
			767 => x"00000c01",
			768 => x"0c061408",
			769 => x"03054f04",
			770 => x"00000c15",
			771 => x"fff70c15",
			772 => x"00000c15",
			773 => x"0a016608",
			774 => x"0c054304",
			775 => x"016e0c31",
			776 => x"00000c31",
			777 => x"0900f704",
			778 => x"fff00c31",
			779 => x"00000c31",
			780 => x"0900f308",
			781 => x"0405d204",
			782 => x"00000c4d",
			783 => x"ff980c4d",
			784 => x"0f069f04",
			785 => x"00c70c4d",
			786 => x"00000c4d",
			787 => x"02061a08",
			788 => x"0c04d004",
			789 => x"00000c69",
			790 => x"00940c69",
			791 => x"0c052a04",
			792 => x"ffe30c69",
			793 => x"00000c69",
			794 => x"02061a08",
			795 => x"0c04d004",
			796 => x"00000c85",
			797 => x"004e0c85",
			798 => x"09012004",
			799 => x"ffad0c85",
			800 => x"00000c85",
			801 => x"0900f70c",
			802 => x"02059a04",
			803 => x"00000ca1",
			804 => x"01009704",
			805 => x"ff940ca1",
			806 => x"00000ca1",
			807 => x"00000ca1",
			808 => x"01009204",
			809 => x"00000cbd",
			810 => x"0e073b08",
			811 => x"07051b04",
			812 => x"00000cbd",
			813 => x"00530cbd",
			814 => x"00000cbd",
			815 => x"0406a304",
			816 => x"00000cd9",
			817 => x"00021b04",
			818 => x"00000cd9",
			819 => x"0f067a04",
			820 => x"00000cd9",
			821 => x"fff70cd9",
			822 => x"00021b08",
			823 => x"0c054304",
			824 => x"00aa0cfd",
			825 => x"00000cfd",
			826 => x"0100a108",
			827 => x"0c056204",
			828 => x"ff2e0cfd",
			829 => x"00000cfd",
			830 => x"00000cfd",
			831 => x"00021b08",
			832 => x"0c054304",
			833 => x"00b20d21",
			834 => x"00000d21",
			835 => x"0100a108",
			836 => x"0c056204",
			837 => x"ff870d21",
			838 => x"00000d21",
			839 => x"00000d21",
			840 => x"02077710",
			841 => x"01009b08",
			842 => x"0801b004",
			843 => x"00000d45",
			844 => x"ffe40d45",
			845 => x"0e05c304",
			846 => x"00000d45",
			847 => x"005e0d45",
			848 => x"ff8d0d45",
			849 => x"0f062f0c",
			850 => x"0c04d004",
			851 => x"00000d71",
			852 => x"00046404",
			853 => x"00a10d71",
			854 => x"00000d71",
			855 => x"09012008",
			856 => x"0100ad04",
			857 => x"ffd00d71",
			858 => x"00000d71",
			859 => x"00000d71",
			860 => x"0900f304",
			861 => x"00000d95",
			862 => x"0901740c",
			863 => x"0d083808",
			864 => x"0d063804",
			865 => x"00000d95",
			866 => x"002b0d95",
			867 => x"00000d95",
			868 => x"00000d95",
			869 => x"0900f304",
			870 => x"ffe90db9",
			871 => x"0901740c",
			872 => x"0d083808",
			873 => x"0d064704",
			874 => x"00000db9",
			875 => x"00140db9",
			876 => x"00000db9",
			877 => x"00000db9",
			878 => x"0b053508",
			879 => x"0a014504",
			880 => x"00000de5",
			881 => x"ff9f0de5",
			882 => x"0002cc0c",
			883 => x"0900f304",
			884 => x"00000de5",
			885 => x"0e087f04",
			886 => x"00440de5",
			887 => x"00000de5",
			888 => x"00000de5",
			889 => x"01009210",
			890 => x"02059a04",
			891 => x"00000e11",
			892 => x"0b058508",
			893 => x"07054904",
			894 => x"ff7f0e11",
			895 => x"00000e11",
			896 => x"00000e11",
			897 => x"0406ea04",
			898 => x"01180e11",
			899 => x"00000e11",
			900 => x"0c052808",
			901 => x"0100a104",
			902 => x"ffbc0e3d",
			903 => x"00000e3d",
			904 => x"0100e50c",
			905 => x"0c061508",
			906 => x"0900e004",
			907 => x"00000e3d",
			908 => x"004b0e3d",
			909 => x"00000e3d",
			910 => x"00000e3d",
			911 => x"01009208",
			912 => x"0b058504",
			913 => x"ffd80e69",
			914 => x"00000e69",
			915 => x"0100e50c",
			916 => x"0507c908",
			917 => x"05060804",
			918 => x"00000e69",
			919 => x"000e0e69",
			920 => x"00000e69",
			921 => x"00000e69",
			922 => x"00028d14",
			923 => x"0900f30c",
			924 => x"0e059d04",
			925 => x"00000e95",
			926 => x"07051a04",
			927 => x"00000e95",
			928 => x"ffb40e95",
			929 => x"0f06de04",
			930 => x"00d60e95",
			931 => x"00000e95",
			932 => x"ff1d0e95",
			933 => x"0100920c",
			934 => x"0305a004",
			935 => x"00000ec9",
			936 => x"07054904",
			937 => x"ffba0ec9",
			938 => x"00000ec9",
			939 => x"0100e50c",
			940 => x"0308e708",
			941 => x"07050404",
			942 => x"00000ec9",
			943 => x"00170ec9",
			944 => x"00000ec9",
			945 => x"00000ec9",
			946 => x"00028d14",
			947 => x"0e071510",
			948 => x"0c04d008",
			949 => x"0f057204",
			950 => x"02250ef5",
			951 => x"003f0ef5",
			952 => x"0f06de04",
			953 => x"02cb0ef5",
			954 => x"01c90ef5",
			955 => x"06c20ef5",
			956 => x"fe5f0ef5",
			957 => x"02076714",
			958 => x"04062704",
			959 => x"00a20f29",
			960 => x"0100a10c",
			961 => x"07055d08",
			962 => x"0600e804",
			963 => x"00000f29",
			964 => x"ff3e0f29",
			965 => x"00000f29",
			966 => x"00940f29",
			967 => x"07069b04",
			968 => x"fedc0f29",
			969 => x"00000f29",
			970 => x"0406ea14",
			971 => x"0900f710",
			972 => x"0305b904",
			973 => x"00000f5d",
			974 => x"01009708",
			975 => x"07051a04",
			976 => x"00000f5d",
			977 => x"ffb60f5d",
			978 => x"00000f5d",
			979 => x"006c0f5d",
			980 => x"09012004",
			981 => x"ff120f5d",
			982 => x"00000f5d",
			983 => x"01009208",
			984 => x"0b058504",
			985 => x"ffda0f91",
			986 => x"00000f91",
			987 => x"0100e510",
			988 => x"0507d70c",
			989 => x"0c061508",
			990 => x"05060604",
			991 => x"00000f91",
			992 => x"00110f91",
			993 => x"00000f91",
			994 => x"00000f91",
			995 => x"00000f91",
			996 => x"0408ab14",
			997 => x"04062704",
			998 => x"00960fbd",
			999 => x"0900f304",
			1000 => x"ff390fbd",
			1001 => x"0f067a04",
			1002 => x"00b30fbd",
			1003 => x"0100a104",
			1004 => x"ff830fbd",
			1005 => x"000c0fbd",
			1006 => x"feef0fbd",
			1007 => x"00028d18",
			1008 => x"0406ea0c",
			1009 => x"0e060f04",
			1010 => x"01d81001",
			1011 => x"0d068404",
			1012 => x"ff871001",
			1013 => x"01be1001",
			1014 => x"0c054304",
			1015 => x"fcc61001",
			1016 => x"0100ba04",
			1017 => x"00ff1001",
			1018 => x"02501001",
			1019 => x"0408ab08",
			1020 => x"0002b704",
			1021 => x"fe851001",
			1022 => x"05b51001",
			1023 => x"fe641001",
			1024 => x"0100920c",
			1025 => x"0b058508",
			1026 => x"07054904",
			1027 => x"ffd0103d",
			1028 => x"0000103d",
			1029 => x"0000103d",
			1030 => x"0100e510",
			1031 => x"0507d70c",
			1032 => x"0c061508",
			1033 => x"07050404",
			1034 => x"0000103d",
			1035 => x"0014103d",
			1036 => x"0000103d",
			1037 => x"0000103d",
			1038 => x"0000103d",
			1039 => x"0100920c",
			1040 => x"0e059d04",
			1041 => x"00001079",
			1042 => x"0b058504",
			1043 => x"ffbb1079",
			1044 => x"00001079",
			1045 => x"0100e510",
			1046 => x"0e087f0c",
			1047 => x"0507c908",
			1048 => x"05060804",
			1049 => x"00001079",
			1050 => x"001a1079",
			1051 => x"00001079",
			1052 => x"00001079",
			1053 => x"00001079",
			1054 => x"00028d18",
			1055 => x"0f060a08",
			1056 => x"01007904",
			1057 => x"002910ad",
			1058 => x"019410ad",
			1059 => x"0900fb04",
			1060 => x"fe2f10ad",
			1061 => x"0f070104",
			1062 => x"019310ad",
			1063 => x"0100be04",
			1064 => x"fe3c10ad",
			1065 => x"015410ad",
			1066 => x"fe6810ad",
			1067 => x"00028d14",
			1068 => x"0c04d004",
			1069 => x"000010f1",
			1070 => x"0207770c",
			1071 => x"03075408",
			1072 => x"0f06de04",
			1073 => x"020510f1",
			1074 => x"015710f1",
			1075 => x"046510f1",
			1076 => x"fe7110f1",
			1077 => x"0408ea0c",
			1078 => x"0a01d704",
			1079 => x"fe6c10f1",
			1080 => x"08024704",
			1081 => x"05b110f1",
			1082 => x"ff6e10f1",
			1083 => x"fe6210f1",
			1084 => x"0a01b61c",
			1085 => x"0100a114",
			1086 => x"03064808",
			1087 => x"0c04d004",
			1088 => x"fff5112d",
			1089 => x"0197112d",
			1090 => x"07055d08",
			1091 => x"0600eb04",
			1092 => x"fd78112d",
			1093 => x"ff1d112d",
			1094 => x"0074112d",
			1095 => x"02076704",
			1096 => x"0194112d",
			1097 => x"ff36112d",
			1098 => x"fe68112d",
			1099 => x"02066104",
			1100 => x"00ff1161",
			1101 => x"0100a104",
			1102 => x"fe941161",
			1103 => x"0408ea10",
			1104 => x"07065808",
			1105 => x"0f077b04",
			1106 => x"00451161",
			1107 => x"ff921161",
			1108 => x"0a01d404",
			1109 => x"00001161",
			1110 => x"008c1161",
			1111 => x"ffc51161",
			1112 => x"0a01b618",
			1113 => x"0f077b14",
			1114 => x"0c04ce04",
			1115 => x"000f11a5",
			1116 => x"0f07250c",
			1117 => x"0f06f308",
			1118 => x"0f06d904",
			1119 => x"01d211a5",
			1120 => x"00ee11a5",
			1121 => x"fff411a5",
			1122 => x"034a11a5",
			1123 => x"fe9211a5",
			1124 => x"0408ab08",
			1125 => x"04089204",
			1126 => x"fe8e11a5",
			1127 => x"001e11a5",
			1128 => x"fe6311a5",
			1129 => x"0002cc20",
			1130 => x"0100a110",
			1131 => x"0f062f08",
			1132 => x"0c054304",
			1133 => x"014c11e9",
			1134 => x"000011e9",
			1135 => x"01009d04",
			1136 => x"fe5311e9",
			1137 => x"000011e9",
			1138 => x"0e087f0c",
			1139 => x"09016f08",
			1140 => x"0f077b04",
			1141 => x"012a11e9",
			1142 => x"000011e9",
			1143 => x"026811e9",
			1144 => x"000011e9",
			1145 => x"fe7511e9",
			1146 => x"0b053508",
			1147 => x"0405d204",
			1148 => x"0000122d",
			1149 => x"ff54122d",
			1150 => x"02066104",
			1151 => x"0065122d",
			1152 => x"0c06140c",
			1153 => x"0c04e904",
			1154 => x"0000122d",
			1155 => x"0c054804",
			1156 => x"ffb1122d",
			1157 => x"0000122d",
			1158 => x"0c061508",
			1159 => x"0b06cf04",
			1160 => x"0000122d",
			1161 => x"002a122d",
			1162 => x"0000122d",
			1163 => x"0002c420",
			1164 => x"00021b0c",
			1165 => x"0c054304",
			1166 => x"016a1271",
			1167 => x"0c054504",
			1168 => x"fef81271",
			1169 => x"00bf1271",
			1170 => x"09010f04",
			1171 => x"fedf1271",
			1172 => x"0f087a0c",
			1173 => x"0c052a04",
			1174 => x"00001271",
			1175 => x"07057504",
			1176 => x"00001271",
			1177 => x"017b1271",
			1178 => x"ffa01271",
			1179 => x"fe6c1271",
			1180 => x"0a01b624",
			1181 => x"0406ea14",
			1182 => x"07050104",
			1183 => x"005f12d5",
			1184 => x"0d066b04",
			1185 => x"01a812d5",
			1186 => x"0d067704",
			1187 => x"ff6212d5",
			1188 => x"0d067b04",
			1189 => x"00d912d5",
			1190 => x"01a412d5",
			1191 => x"09012008",
			1192 => x"05068904",
			1193 => x"fd6412d5",
			1194 => x"ff3c12d5",
			1195 => x"0e073b04",
			1196 => x"01b112d5",
			1197 => x"000012d5",
			1198 => x"0408ea0c",
			1199 => x"0a01db04",
			1200 => x"fe9212d5",
			1201 => x"0408db04",
			1202 => x"000012d5",
			1203 => x"0d5e12d5",
			1204 => x"fe6612d5",
			1205 => x"00028d20",
			1206 => x"02069d14",
			1207 => x"07050104",
			1208 => x"001e1339",
			1209 => x"03064804",
			1210 => x"01a01339",
			1211 => x"0d067704",
			1212 => x"fe8d1339",
			1213 => x"0d067b04",
			1214 => x"00761339",
			1215 => x"01981339",
			1216 => x"0100a804",
			1217 => x"fddb1339",
			1218 => x"0e072504",
			1219 => x"01931339",
			1220 => x"00491339",
			1221 => x"08024710",
			1222 => x"0a01db04",
			1223 => x"fe9e1339",
			1224 => x"0002c404",
			1225 => x"00001339",
			1226 => x"0a01df04",
			1227 => x"06381339",
			1228 => x"00001339",
			1229 => x"fe671339",
			1230 => x"08024728",
			1231 => x"01009b18",
			1232 => x"0e059d08",
			1233 => x"01006f04",
			1234 => x"0000138d",
			1235 => x"0085138d",
			1236 => x"01009204",
			1237 => x"ff14138d",
			1238 => x"01009504",
			1239 => x"0047138d",
			1240 => x"07054b04",
			1241 => x"0000138d",
			1242 => x"ff4d138d",
			1243 => x"0e087f0c",
			1244 => x"0507d708",
			1245 => x"02088b04",
			1246 => x"00a7138d",
			1247 => x"0000138d",
			1248 => x"0000138d",
			1249 => x"0000138d",
			1250 => x"fec9138d",
			1251 => x"0002cc20",
			1252 => x"0b06cf18",
			1253 => x"0f060a04",
			1254 => x"016313d1",
			1255 => x"0900fb04",
			1256 => x"feb313d1",
			1257 => x"0f070104",
			1258 => x"014b13d1",
			1259 => x"06010c04",
			1260 => x"ff6a13d1",
			1261 => x"06011904",
			1262 => x"005e13d1",
			1263 => x"000013d1",
			1264 => x"0e087f04",
			1265 => x"02cf13d1",
			1266 => x"000013d1",
			1267 => x"fe7313d1",
			1268 => x"0408ea24",
			1269 => x"0c06141c",
			1270 => x"02077718",
			1271 => x"01009910",
			1272 => x"04062708",
			1273 => x"0c04cf04",
			1274 => x"0000141d",
			1275 => x"0188141d",
			1276 => x"0900f304",
			1277 => x"fdce141d",
			1278 => x"ffde141d",
			1279 => x"0f070104",
			1280 => x"0190141d",
			1281 => x"008b141d",
			1282 => x"fec8141d",
			1283 => x"0b06cc04",
			1284 => x"0000141d",
			1285 => x"057d141d",
			1286 => x"fe69141d",
			1287 => x"0408ea24",
			1288 => x"0406a308",
			1289 => x"0c04d004",
			1290 => x"00001469",
			1291 => x"01071469",
			1292 => x"0100ad08",
			1293 => x"0c04e904",
			1294 => x"00001469",
			1295 => x"ff251469",
			1296 => x"0e087f10",
			1297 => x"0c054604",
			1298 => x"00001469",
			1299 => x"0100e508",
			1300 => x"0308e704",
			1301 => x"00711469",
			1302 => x"00001469",
			1303 => x"00001469",
			1304 => x"00001469",
			1305 => x"feae1469",
			1306 => x"0408ab20",
			1307 => x"01006f04",
			1308 => x"fe2214ad",
			1309 => x"02076714",
			1310 => x"01009210",
			1311 => x"0f05d20c",
			1312 => x"0e059d04",
			1313 => x"01ad14ad",
			1314 => x"0e05ac04",
			1315 => x"000014ad",
			1316 => x"012914ad",
			1317 => x"fe1114ad",
			1318 => x"019114ad",
			1319 => x"07064404",
			1320 => x"fe9514ad",
			1321 => x"037314ad",
			1322 => x"fe6614ad",
			1323 => x"0a01df28",
			1324 => x"0100a610",
			1325 => x"0e059d08",
			1326 => x"01006c04",
			1327 => x"00001501",
			1328 => x"00291501",
			1329 => x"01009204",
			1330 => x"ff631501",
			1331 => x"00001501",
			1332 => x"0308e714",
			1333 => x"09010f04",
			1334 => x"00001501",
			1335 => x"0c052704",
			1336 => x"00001501",
			1337 => x"0507c908",
			1338 => x"0100e504",
			1339 => x"009a1501",
			1340 => x"00001501",
			1341 => x"00001501",
			1342 => x"00001501",
			1343 => x"ff111501",
			1344 => x"0408ea24",
			1345 => x"01007908",
			1346 => x"02059a04",
			1347 => x"0000154d",
			1348 => x"fe8a154d",
			1349 => x"0b059904",
			1350 => x"0158154d",
			1351 => x"0c052a08",
			1352 => x"0100a104",
			1353 => x"fef3154d",
			1354 => x"0000154d",
			1355 => x"02088b0c",
			1356 => x"0100a604",
			1357 => x"0000154d",
			1358 => x"0600f204",
			1359 => x"0000154d",
			1360 => x"0124154d",
			1361 => x"0000154d",
			1362 => x"fe80154d",
			1363 => x"08024728",
			1364 => x"0100a110",
			1365 => x"00021b0c",
			1366 => x"0c04d004",
			1367 => x"ff9415a1",
			1368 => x"0c054304",
			1369 => x"013815a1",
			1370 => x"000015a1",
			1371 => x"fe9e15a1",
			1372 => x"0e087f14",
			1373 => x"0600f104",
			1374 => x"000015a1",
			1375 => x"0100a604",
			1376 => x"000015a1",
			1377 => x"0c052704",
			1378 => x"000015a1",
			1379 => x"0507c904",
			1380 => x"013f15a1",
			1381 => x"000015a1",
			1382 => x"000015a1",
			1383 => x"fe7d15a1",
			1384 => x"0002cc24",
			1385 => x"0c04d004",
			1386 => x"ff9615ed",
			1387 => x"0f067a0c",
			1388 => x"0900f308",
			1389 => x"0900ef04",
			1390 => x"007715ed",
			1391 => x"000015ed",
			1392 => x"013c15ed",
			1393 => x"0c052a04",
			1394 => x"ff8e15ed",
			1395 => x"0e087f0c",
			1396 => x"09011b04",
			1397 => x"000015ed",
			1398 => x"0308e704",
			1399 => x"00d215ed",
			1400 => x"000015ed",
			1401 => x"000015ed",
			1402 => x"fe8c15ed",
			1403 => x"0002cc30",
			1404 => x"0100a618",
			1405 => x"00021b10",
			1406 => x"0c04d004",
			1407 => x"ff681653",
			1408 => x"0c054304",
			1409 => x"014b1653",
			1410 => x"0d067704",
			1411 => x"ffff1653",
			1412 => x"00001653",
			1413 => x"0100a104",
			1414 => x"fe771653",
			1415 => x"00001653",
			1416 => x"0e087f14",
			1417 => x"0600f104",
			1418 => x"00001653",
			1419 => x"0c052704",
			1420 => x"00001653",
			1421 => x"0507c908",
			1422 => x"0308e704",
			1423 => x"01721653",
			1424 => x"00001653",
			1425 => x"00001653",
			1426 => x"00001653",
			1427 => x"fe781653",
			1428 => x"00001655",
			1429 => x"00001659",
			1430 => x"0000165d",
			1431 => x"00001661",
			1432 => x"00001665",
			1433 => x"00001669",
			1434 => x"0000166d",
			1435 => x"00001671",
			1436 => x"00001675",
			1437 => x"00001679",
			1438 => x"0000167d",
			1439 => x"00001681",
			1440 => x"00001685",
			1441 => x"00001689",
			1442 => x"0000168d",
			1443 => x"00001691",
			1444 => x"00001695",
			1445 => x"00001699",
			1446 => x"0000169d",
			1447 => x"000016a1",
			1448 => x"000016a5",
			1449 => x"00021b04",
			1450 => x"000016b1",
			1451 => x"ffe716b1",
			1452 => x"00021b04",
			1453 => x"002a16bd",
			1454 => x"000016bd",
			1455 => x"0c052504",
			1456 => x"fff816c9",
			1457 => x"000016c9",
			1458 => x"0405d204",
			1459 => x"000016d5",
			1460 => x"fffc16d5",
			1461 => x"0f060a04",
			1462 => x"000016e1",
			1463 => x"ffe516e1",
			1464 => x"0406ea04",
			1465 => x"000e16ed",
			1466 => x"000016ed",
			1467 => x"02061a04",
			1468 => x"003016f9",
			1469 => x"000016f9",
			1470 => x"0406a304",
			1471 => x"0067170d",
			1472 => x"07058c04",
			1473 => x"ff87170d",
			1474 => x"0000170d",
			1475 => x"0406a304",
			1476 => x"00a31721",
			1477 => x"09011304",
			1478 => x"ffcc1721",
			1479 => x"00001721",
			1480 => x"0d067704",
			1481 => x"fffb1735",
			1482 => x"0d083804",
			1483 => x"00011735",
			1484 => x"00001735",
			1485 => x"02061a08",
			1486 => x"0f05b604",
			1487 => x"00001749",
			1488 => x"00021749",
			1489 => x"ffff1749",
			1490 => x"0900f304",
			1491 => x"fff3175d",
			1492 => x"09017404",
			1493 => x"0006175d",
			1494 => x"0000175d",
			1495 => x"02061a08",
			1496 => x"01009204",
			1497 => x"00001779",
			1498 => x"01411779",
			1499 => x"0900f704",
			1500 => x"fff21779",
			1501 => x"00001779",
			1502 => x"0900f308",
			1503 => x"0405d204",
			1504 => x"00001795",
			1505 => x"ffa41795",
			1506 => x"0f069f04",
			1507 => x"00a61795",
			1508 => x"00001795",
			1509 => x"02061a08",
			1510 => x"0c04d004",
			1511 => x"000017b1",
			1512 => x"005d17b1",
			1513 => x"07069b04",
			1514 => x"ffa017b1",
			1515 => x"000017b1",
			1516 => x"0406a304",
			1517 => x"007017cd",
			1518 => x"0100a108",
			1519 => x"05068904",
			1520 => x"ff3c17cd",
			1521 => x"000017cd",
			1522 => x"000017cd",
			1523 => x"0900f70c",
			1524 => x"02059a04",
			1525 => x"000017e9",
			1526 => x"01009704",
			1527 => x"ffa117e9",
			1528 => x"000017e9",
			1529 => x"000017e9",
			1530 => x"0900f30c",
			1531 => x"0405d204",
			1532 => x"00001805",
			1533 => x"01009704",
			1534 => x"ffb21805",
			1535 => x"00001805",
			1536 => x"00001805",
			1537 => x"0406a304",
			1538 => x"00001821",
			1539 => x"00021b04",
			1540 => x"00001821",
			1541 => x"0f067a04",
			1542 => x"00001821",
			1543 => x"fff91821",
			1544 => x"00021b08",
			1545 => x"0c054304",
			1546 => x"00c61845",
			1547 => x"00001845",
			1548 => x"0100a108",
			1549 => x"0c056204",
			1550 => x"ff791845",
			1551 => x"00001845",
			1552 => x"00001845",
			1553 => x"0100920c",
			1554 => x"0e059d04",
			1555 => x"00001869",
			1556 => x"0b058504",
			1557 => x"ffc31869",
			1558 => x"00001869",
			1559 => x"0e064304",
			1560 => x"00171869",
			1561 => x"00001869",
			1562 => x"02077710",
			1563 => x"01009b08",
			1564 => x"0801b004",
			1565 => x"0000188d",
			1566 => x"ffea188d",
			1567 => x"0e05c304",
			1568 => x"0000188d",
			1569 => x"0057188d",
			1570 => x"ff95188d",
			1571 => x"08024710",
			1572 => x"0900b304",
			1573 => x"000018b1",
			1574 => x"0308e708",
			1575 => x"0900f304",
			1576 => x"000018b1",
			1577 => x"009718b1",
			1578 => x"000018b1",
			1579 => x"ff4c18b1",
			1580 => x"0900f304",
			1581 => x"000018d5",
			1582 => x"0901740c",
			1583 => x"0d083808",
			1584 => x"0d063804",
			1585 => x"000018d5",
			1586 => x"002718d5",
			1587 => x"000018d5",
			1588 => x"000018d5",
			1589 => x"0900f304",
			1590 => x"ffed18f9",
			1591 => x"0901740c",
			1592 => x"0d083808",
			1593 => x"0d064704",
			1594 => x"000018f9",
			1595 => x"000d18f9",
			1596 => x"000018f9",
			1597 => x"000018f9",
			1598 => x"0900fb08",
			1599 => x"01009b04",
			1600 => x"ffdd1925",
			1601 => x"00001925",
			1602 => x"0100e50c",
			1603 => x"0507d708",
			1604 => x"07051f04",
			1605 => x"00001925",
			1606 => x"00261925",
			1607 => x"00001925",
			1608 => x"00001925",
			1609 => x"01009210",
			1610 => x"0f05ad04",
			1611 => x"00001951",
			1612 => x"0b058508",
			1613 => x"07054904",
			1614 => x"ff8a1951",
			1615 => x"00001951",
			1616 => x"00001951",
			1617 => x"0f06de04",
			1618 => x"01021951",
			1619 => x"00001951",
			1620 => x"0c052808",
			1621 => x"0100a104",
			1622 => x"ffc4197d",
			1623 => x"0000197d",
			1624 => x"0100e50c",
			1625 => x"0c061508",
			1626 => x"0900e004",
			1627 => x"0000197d",
			1628 => x"003f197d",
			1629 => x"0000197d",
			1630 => x"0000197d",
			1631 => x"0900f30c",
			1632 => x"02059a08",
			1633 => x"08019004",
			1634 => x"006f19b1",
			1635 => x"000019b1",
			1636 => x"fe9b19b1",
			1637 => x"02076708",
			1638 => x"0900fb04",
			1639 => x"000019b1",
			1640 => x"00d919b1",
			1641 => x"07069b04",
			1642 => x"ff4719b1",
			1643 => x"000019b1",
			1644 => x"0900fb0c",
			1645 => x"0e059d04",
			1646 => x"000019e5",
			1647 => x"01009b04",
			1648 => x"ffbf19e5",
			1649 => x"000019e5",
			1650 => x"0100e50c",
			1651 => x"0e087f08",
			1652 => x"07051f04",
			1653 => x"000019e5",
			1654 => x"003719e5",
			1655 => x"000019e5",
			1656 => x"000019e5",
			1657 => x"0c05280c",
			1658 => x"0f05ad04",
			1659 => x"00001a19",
			1660 => x"0100a104",
			1661 => x"ff9a1a19",
			1662 => x"00001a19",
			1663 => x"01009304",
			1664 => x"00001a19",
			1665 => x"02088b08",
			1666 => x"0100e504",
			1667 => x"00931a19",
			1668 => x"00001a19",
			1669 => x"00001a19",
			1670 => x"00028d10",
			1671 => x"0c04d004",
			1672 => x"00001a55",
			1673 => x"0f077b08",
			1674 => x"02071704",
			1675 => x"02201a55",
			1676 => x"06581a55",
			1677 => x"fe691a55",
			1678 => x"0408ea0c",
			1679 => x"08024104",
			1680 => x"fe6a1a55",
			1681 => x"08024704",
			1682 => x"0b9d1a55",
			1683 => x"ff281a55",
			1684 => x"fe611a55",
			1685 => x"0408ea18",
			1686 => x"0900f30c",
			1687 => x"0f060a08",
			1688 => x"07050104",
			1689 => x"00001a89",
			1690 => x"00891a89",
			1691 => x"ffae1a89",
			1692 => x"07054904",
			1693 => x"00001a89",
			1694 => x"0e087f04",
			1695 => x"00f21a89",
			1696 => x"00001a89",
			1697 => x"ff381a89",
			1698 => x"01009b08",
			1699 => x"0801b004",
			1700 => x"00001abd",
			1701 => x"ff1e1abd",
			1702 => x"02088b10",
			1703 => x"0600f104",
			1704 => x"00001abd",
			1705 => x"0100e508",
			1706 => x"0507d704",
			1707 => x"00871abd",
			1708 => x"00001abd",
			1709 => x"00001abd",
			1710 => x"00001abd",
			1711 => x"0900f308",
			1712 => x"07055d04",
			1713 => x"ffe51af1",
			1714 => x"00001af1",
			1715 => x"09017410",
			1716 => x"0507d70c",
			1717 => x"07051f04",
			1718 => x"00001af1",
			1719 => x"0c061504",
			1720 => x"002c1af1",
			1721 => x"00001af1",
			1722 => x"00001af1",
			1723 => x"00001af1",
			1724 => x"00021b04",
			1725 => x"007f1b1d",
			1726 => x"0100a104",
			1727 => x"ff541b1d",
			1728 => x"02088b0c",
			1729 => x"06013808",
			1730 => x"0507c904",
			1731 => x"00401b1d",
			1732 => x"00001b1d",
			1733 => x"00001b1d",
			1734 => x"00001b1d",
			1735 => x"00028d14",
			1736 => x"0406ea0c",
			1737 => x"04062704",
			1738 => x"01a41b61",
			1739 => x"0900fb04",
			1740 => x"feed1b61",
			1741 => x"01a11b61",
			1742 => x"09012004",
			1743 => x"fe011b61",
			1744 => x"017f1b61",
			1745 => x"0408ea0c",
			1746 => x"0a01db04",
			1747 => x"fe9a1b61",
			1748 => x"0408db04",
			1749 => x"00001b61",
			1750 => x"082a1b61",
			1751 => x"fe671b61",
			1752 => x"0900f30c",
			1753 => x"01009708",
			1754 => x"07055d04",
			1755 => x"ffd81b9d",
			1756 => x"00001b9d",
			1757 => x"00001b9d",
			1758 => x"0100e510",
			1759 => x"0507d70c",
			1760 => x"07051f04",
			1761 => x"00001b9d",
			1762 => x"0c061504",
			1763 => x"00331b9d",
			1764 => x"00001b9d",
			1765 => x"00001b9d",
			1766 => x"00001b9d",
			1767 => x"0900f314",
			1768 => x"0406270c",
			1769 => x"0405d204",
			1770 => x"00591be9",
			1771 => x"0600df04",
			1772 => x"ff921be9",
			1773 => x"00001be9",
			1774 => x"01009704",
			1775 => x"fe921be9",
			1776 => x"00001be9",
			1777 => x"0e073b0c",
			1778 => x"0900fb04",
			1779 => x"00001be9",
			1780 => x"0002cc04",
			1781 => x"00c71be9",
			1782 => x"00001be9",
			1783 => x"07069b04",
			1784 => x"ff6a1be9",
			1785 => x"00001be9",
			1786 => x"02076718",
			1787 => x"04062704",
			1788 => x"00b41c25",
			1789 => x"0900f308",
			1790 => x"0600ea04",
			1791 => x"ff0e1c25",
			1792 => x"00001c25",
			1793 => x"0f067a04",
			1794 => x"00ba1c25",
			1795 => x"0c054304",
			1796 => x"ff9c1c25",
			1797 => x"00121c25",
			1798 => x"07069b04",
			1799 => x"fed31c25",
			1800 => x"00001c25",
			1801 => x"0207671c",
			1802 => x"0900fb14",
			1803 => x"0f05ad08",
			1804 => x"01006f04",
			1805 => x"00001c69",
			1806 => x"00881c69",
			1807 => x"0900f308",
			1808 => x"07051a04",
			1809 => x"00001c69",
			1810 => x"ff071c69",
			1811 => x"00001c69",
			1812 => x"0f070104",
			1813 => x"00db1c69",
			1814 => x"00001c69",
			1815 => x"07069b04",
			1816 => x"feb71c69",
			1817 => x"00001c69",
			1818 => x"0408ab1c",
			1819 => x"0100990c",
			1820 => x"04062708",
			1821 => x"0600cd04",
			1822 => x"00001ca5",
			1823 => x"015c1ca5",
			1824 => x"feed1ca5",
			1825 => x"0f070104",
			1826 => x"016a1ca5",
			1827 => x"03076c04",
			1828 => x"ff8d1ca5",
			1829 => x"0f087a04",
			1830 => x"00961ca5",
			1831 => x"00001ca5",
			1832 => x"fe6f1ca5",
			1833 => x"01009b18",
			1834 => x"0f060a0c",
			1835 => x"0c04cf04",
			1836 => x"00001cf9",
			1837 => x"06011c04",
			1838 => x"002c1cf9",
			1839 => x"00001cf9",
			1840 => x"0c056008",
			1841 => x"0600e604",
			1842 => x"00001cf9",
			1843 => x"ff081cf9",
			1844 => x"00001cf9",
			1845 => x"02088b10",
			1846 => x"0600f104",
			1847 => x"00001cf9",
			1848 => x"0100e508",
			1849 => x"0e087f04",
			1850 => x"00a91cf9",
			1851 => x"00001cf9",
			1852 => x"00001cf9",
			1853 => x"00001cf9",
			1854 => x"0408ab20",
			1855 => x"01009910",
			1856 => x"04062708",
			1857 => x"0600cd04",
			1858 => x"00001d3d",
			1859 => x"01551d3d",
			1860 => x"01009204",
			1861 => x"fea11d3d",
			1862 => x"ffd51d3d",
			1863 => x"0f070104",
			1864 => x"01641d3d",
			1865 => x"0d071604",
			1866 => x"ffbb1d3d",
			1867 => x"0f087a04",
			1868 => x"00a11d3d",
			1869 => x"00001d3d",
			1870 => x"fe711d3d",
			1871 => x"0002cc20",
			1872 => x"0100a110",
			1873 => x"0f062f08",
			1874 => x"0c054304",
			1875 => x"013c1d81",
			1876 => x"00001d81",
			1877 => x"01009d04",
			1878 => x"fe741d81",
			1879 => x"00001d81",
			1880 => x"0308e70c",
			1881 => x"0600f104",
			1882 => x"00001d81",
			1883 => x"02088b04",
			1884 => x"017e1d81",
			1885 => x"00001d81",
			1886 => x"00001d81",
			1887 => x"fe771d81",
			1888 => x"00021b04",
			1889 => x"00861db5",
			1890 => x"0100a104",
			1891 => x"ff4a1db5",
			1892 => x"06013610",
			1893 => x"0e087f0c",
			1894 => x"0507c908",
			1895 => x"0c052704",
			1896 => x"00001db5",
			1897 => x"00511db5",
			1898 => x"00001db5",
			1899 => x"00001db5",
			1900 => x"00001db5",
			1901 => x"00028d1c",
			1902 => x"0f077b18",
			1903 => x"0f072514",
			1904 => x"0406ea0c",
			1905 => x"0f069f04",
			1906 => x"01ed1e01",
			1907 => x"0e068d04",
			1908 => x"00651e01",
			1909 => x"01d21e01",
			1910 => x"06010004",
			1911 => x"fdec1e01",
			1912 => x"01eb1e01",
			1913 => x"03d81e01",
			1914 => x"fe841e01",
			1915 => x"0408ab08",
			1916 => x"04089204",
			1917 => x"fe871e01",
			1918 => x"00011e01",
			1919 => x"fe621e01",
			1920 => x"00028d18",
			1921 => x"09014114",
			1922 => x"0f076d10",
			1923 => x"0c04d004",
			1924 => x"00191e55",
			1925 => x"0f06f308",
			1926 => x"0f06de04",
			1927 => x"024e1e55",
			1928 => x"019b1e55",
			1929 => x"03201e55",
			1930 => x"fe5b1e55",
			1931 => x"05cb1e55",
			1932 => x"0002cc10",
			1933 => x"08024104",
			1934 => x"fe671e55",
			1935 => x"08024708",
			1936 => x"0a01d704",
			1937 => x"ff601e55",
			1938 => x"03641e55",
			1939 => x"ff231e55",
			1940 => x"fe601e55",
			1941 => x"00028d20",
			1942 => x"01007904",
			1943 => x"ff091eb1",
			1944 => x"0f070114",
			1945 => x"01008208",
			1946 => x"0e052604",
			1947 => x"01af1eb1",
			1948 => x"ffc61eb1",
			1949 => x"0e060f04",
			1950 => x"01c01eb1",
			1951 => x"0c052504",
			1952 => x"fff81eb1",
			1953 => x"01c01eb1",
			1954 => x"0705a104",
			1955 => x"fd861eb1",
			1956 => x"021d1eb1",
			1957 => x"0002cc0c",
			1958 => x"08024104",
			1959 => x"fe771eb1",
			1960 => x"08024704",
			1961 => x"02c11eb1",
			1962 => x"ffb71eb1",
			1963 => x"fe651eb1",
			1964 => x"08024728",
			1965 => x"01009b14",
			1966 => x"0801a50c",
			1967 => x"0e059d04",
			1968 => x"00741f05",
			1969 => x"0f05c304",
			1970 => x"ffb11f05",
			1971 => x"00001f05",
			1972 => x"0900f304",
			1973 => x"ff301f05",
			1974 => x"00001f05",
			1975 => x"0e087f10",
			1976 => x"0507d70c",
			1977 => x"0308e708",
			1978 => x"02088b04",
			1979 => x"008f1f05",
			1980 => x"00001f05",
			1981 => x"00001f05",
			1982 => x"00001f05",
			1983 => x"00001f05",
			1984 => x"fed91f05",
			1985 => x"08024720",
			1986 => x"01007908",
			1987 => x"02059a04",
			1988 => x"00001f49",
			1989 => x"ff061f49",
			1990 => x"0f067a04",
			1991 => x"00e91f49",
			1992 => x"0100a604",
			1993 => x"ff541f49",
			1994 => x"0e087f0c",
			1995 => x"0600f704",
			1996 => x"00001f49",
			1997 => x"0507d704",
			1998 => x"00b01f49",
			1999 => x"00001f49",
			2000 => x"00001f49",
			2001 => x"fe941f49",
			2002 => x"0408ea24",
			2003 => x"0c06141c",
			2004 => x"02077718",
			2005 => x"01009910",
			2006 => x"04062708",
			2007 => x"0c04cf04",
			2008 => x"00001f95",
			2009 => x"01841f95",
			2010 => x"0900f304",
			2011 => x"fdfb1f95",
			2012 => x"fff51f95",
			2013 => x"0f070104",
			2014 => x"018c1f95",
			2015 => x"007d1f95",
			2016 => x"fed81f95",
			2017 => x"0b06cc04",
			2018 => x"00001f95",
			2019 => x"03ae1f95",
			2020 => x"fe6a1f95",
			2021 => x"0a01b61c",
			2022 => x"01007904",
			2023 => x"feea1ff1",
			2024 => x"02077714",
			2025 => x"0f061204",
			2026 => x"01cc1ff1",
			2027 => x"01009b04",
			2028 => x"fd661ff1",
			2029 => x"07054908",
			2030 => x"0600f604",
			2031 => x"01b41ff1",
			2032 => x"ff721ff1",
			2033 => x"01d71ff1",
			2034 => x"feb81ff1",
			2035 => x"0408ea10",
			2036 => x"0a01d704",
			2037 => x"fe761ff1",
			2038 => x"0a01df08",
			2039 => x"08024104",
			2040 => x"00001ff1",
			2041 => x"08131ff1",
			2042 => x"ffa91ff1",
			2043 => x"fe641ff1",
			2044 => x"08024720",
			2045 => x"02066104",
			2046 => x"00f22035",
			2047 => x"0100ad08",
			2048 => x"0c04e904",
			2049 => x"00002035",
			2050 => x"ff142035",
			2051 => x"0e087f10",
			2052 => x"0c054604",
			2053 => x"00002035",
			2054 => x"0507d708",
			2055 => x"02088b04",
			2056 => x"007d2035",
			2057 => x"00002035",
			2058 => x"00002035",
			2059 => x"00002035",
			2060 => x"fea82035",
			2061 => x"01009210",
			2062 => x"02059a04",
			2063 => x"000b2099",
			2064 => x"07054908",
			2065 => x"0b058504",
			2066 => x"fed92099",
			2067 => x"00002099",
			2068 => x"00002099",
			2069 => x"00021b04",
			2070 => x"00842099",
			2071 => x"0100a60c",
			2072 => x"0e064304",
			2073 => x"00002099",
			2074 => x"07052f04",
			2075 => x"00002099",
			2076 => x"ff812099",
			2077 => x"02088b10",
			2078 => x"0c052704",
			2079 => x"00002099",
			2080 => x"09011304",
			2081 => x"00002099",
			2082 => x"0100e504",
			2083 => x"00a72099",
			2084 => x"00002099",
			2085 => x"00002099",
			2086 => x"0408ea24",
			2087 => x"01007908",
			2088 => x"02059a04",
			2089 => x"000020e5",
			2090 => x"fe9f20e5",
			2091 => x"0b059904",
			2092 => x"014f20e5",
			2093 => x"0c052a08",
			2094 => x"0100a104",
			2095 => x"ff0f20e5",
			2096 => x"000020e5",
			2097 => x"0e087f0c",
			2098 => x"0100a604",
			2099 => x"000020e5",
			2100 => x"0600f204",
			2101 => x"000020e5",
			2102 => x"011220e5",
			2103 => x"000020e5",
			2104 => x"fe8320e5",
			2105 => x"08024728",
			2106 => x"01007908",
			2107 => x"0f05ad04",
			2108 => x"00002139",
			2109 => x"ff142139",
			2110 => x"0f067a0c",
			2111 => x"0b059904",
			2112 => x"01172139",
			2113 => x"0b05a604",
			2114 => x"00002139",
			2115 => x"005a2139",
			2116 => x"0100a604",
			2117 => x"ff612139",
			2118 => x"0e087f0c",
			2119 => x"0600f704",
			2120 => x"00002139",
			2121 => x"0507d704",
			2122 => x"009f2139",
			2123 => x"00002139",
			2124 => x"00002139",
			2125 => x"fe992139",
			2126 => x"08024728",
			2127 => x"0c061420",
			2128 => x"0207771c",
			2129 => x"01009910",
			2130 => x"0801a508",
			2131 => x"0c04cf04",
			2132 => x"0000218d",
			2133 => x"018d218d",
			2134 => x"0001fa04",
			2135 => x"007e218d",
			2136 => x"fe0f218d",
			2137 => x"07054908",
			2138 => x"0f064204",
			2139 => x"0150218d",
			2140 => x"0000218d",
			2141 => x"0199218d",
			2142 => x"feb7218d",
			2143 => x"0308e704",
			2144 => x"0b20218d",
			2145 => x"0000218d",
			2146 => x"fe69218d",
			2147 => x"0408ab24",
			2148 => x"0900af04",
			2149 => x"ff0a21db",
			2150 => x"0f060a04",
			2151 => x"018921db",
			2152 => x"0705490c",
			2153 => x"0900fe04",
			2154 => x"febf21db",
			2155 => x"0c052504",
			2156 => x"003721db",
			2157 => x"ffc021db",
			2158 => x"0f078104",
			2159 => x"015421db",
			2160 => x"02086c04",
			2161 => x"ff3f21db",
			2162 => x"02087404",
			2163 => x"019521db",
			2164 => x"000021db",
			2165 => x"fe6b21db",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(710, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(1428, initial_addr_3'length));
	end generate gen_rom_3;

	gen_rom_4: if SELECT_ROM = 4 generate
		bank <= (
			0 => x"00000005",
			1 => x"00000009",
			2 => x"0000000d",
			3 => x"00000011",
			4 => x"00000015",
			5 => x"00000019",
			6 => x"0000001d",
			7 => x"00000021",
			8 => x"00000025",
			9 => x"0b071008",
			10 => x"0b06dc04",
			11 => x"00000041",
			12 => x"00220041",
			13 => x"0b086604",
			14 => x"ffe00041",
			15 => x"00000041",
			16 => x"0a01ec08",
			17 => x"0a016e04",
			18 => x"0000005d",
			19 => x"0022005d",
			20 => x"0a028304",
			21 => x"fff7005d",
			22 => x"0000005d",
			23 => x"01009204",
			24 => x"00000079",
			25 => x"0d087f08",
			26 => x"07068304",
			27 => x"ffd90079",
			28 => x"00000079",
			29 => x"00000079",
			30 => x"0508210c",
			31 => x"07065804",
			32 => x"0000009d",
			33 => x"0507c704",
			34 => x"0000009d",
			35 => x"ffca009d",
			36 => x"07076804",
			37 => x"002c009d",
			38 => x"0000009d",
			39 => x"0900f70c",
			40 => x"0e059d04",
			41 => x"000000c1",
			42 => x"0002b704",
			43 => x"001000c1",
			44 => x"000000c1",
			45 => x"06013e04",
			46 => x"ffaf00c1",
			47 => x"000000c1",
			48 => x"07066c08",
			49 => x"07065804",
			50 => x"000000e5",
			51 => x"ffe000e5",
			52 => x"03097804",
			53 => x"000000e5",
			54 => x"030cb804",
			55 => x"000700e5",
			56 => x"000000e5",
			57 => x"0b06d20c",
			58 => x"0c052804",
			59 => x"00000111",
			60 => x"0c061504",
			61 => x"ffeb0111",
			62 => x"00000111",
			63 => x"0100f308",
			64 => x"07069b04",
			65 => x"00310111",
			66 => x"00000111",
			67 => x"00000111",
			68 => x"0a01ec0c",
			69 => x"00021b04",
			70 => x"0000013d",
			71 => x"0002f604",
			72 => x"002b013d",
			73 => x"0000013d",
			74 => x"0a028308",
			75 => x"0002e604",
			76 => x"0000013d",
			77 => x"fff6013d",
			78 => x"0000013d",
			79 => x"0b071010",
			80 => x"0b066304",
			81 => x"00000161",
			82 => x"0100f108",
			83 => x"0100cd04",
			84 => x"00000161",
			85 => x"00310161",
			86 => x"00000161",
			87 => x"00000161",
			88 => x"0409db10",
			89 => x"02092004",
			90 => x"00000185",
			91 => x"02097b08",
			92 => x"08027904",
			93 => x"00320185",
			94 => x"00000185",
			95 => x"00000185",
			96 => x"00000185",
			97 => x"0c052804",
			98 => x"000001a9",
			99 => x"0508210c",
			100 => x"0d087f08",
			101 => x"07068304",
			102 => x"ffbd01a9",
			103 => x"000001a9",
			104 => x"000001a9",
			105 => x"000001a9",
			106 => x"05088610",
			107 => x"0002bf08",
			108 => x"0a018404",
			109 => x"fff501dd",
			110 => x"000101dd",
			111 => x"0a01d704",
			112 => x"000001dd",
			113 => x"ffbf01dd",
			114 => x"06019608",
			115 => x"01013b04",
			116 => x"001201dd",
			117 => x"000001dd",
			118 => x"000001dd",
			119 => x"07066c10",
			120 => x"0f061204",
			121 => x"00000211",
			122 => x"0f097d08",
			123 => x"0b070e04",
			124 => x"ffd30211",
			125 => x"00000211",
			126 => x"00000211",
			127 => x"0f094d08",
			128 => x"0f090d04",
			129 => x"00000211",
			130 => x"00220211",
			131 => x"00000211",
			132 => x"0a01e910",
			133 => x"0a014504",
			134 => x"00000245",
			135 => x"0002e608",
			136 => x"0a01db04",
			137 => x"00100245",
			138 => x"00000245",
			139 => x"00000245",
			140 => x"0002dd04",
			141 => x"00000245",
			142 => x"0a028a04",
			143 => x"fff40245",
			144 => x"00000245",
			145 => x"0308ff0c",
			146 => x"0900f304",
			147 => x"00000279",
			148 => x"01009304",
			149 => x"00000279",
			150 => x"ffea0279",
			151 => x"0209810c",
			152 => x"0b072008",
			153 => x"0100f304",
			154 => x"003f0279",
			155 => x"00000279",
			156 => x"00000279",
			157 => x"00000279",
			158 => x"0a01e40c",
			159 => x"0e059d04",
			160 => x"000002b5",
			161 => x"07051a04",
			162 => x"000002b5",
			163 => x"001d02b5",
			164 => x"03097808",
			165 => x"05082104",
			166 => x"ffee02b5",
			167 => x"000002b5",
			168 => x"05080f04",
			169 => x"000002b5",
			170 => x"0509f004",
			171 => x"000a02b5",
			172 => x"000002b5",
			173 => x"0409db14",
			174 => x"02092004",
			175 => x"000002e9",
			176 => x"0b07200c",
			177 => x"09019008",
			178 => x"0100f304",
			179 => x"006802e9",
			180 => x"000002e9",
			181 => x"000002e9",
			182 => x"000002e9",
			183 => x"0b086704",
			184 => x"fff802e9",
			185 => x"000002e9",
			186 => x"0c052504",
			187 => x"00000315",
			188 => x"05082110",
			189 => x"0d087f0c",
			190 => x"0c063008",
			191 => x"0209ce04",
			192 => x"ffb60315",
			193 => x"00000315",
			194 => x"00000315",
			195 => x"00000315",
			196 => x"00000315",
			197 => x"08032914",
			198 => x"0e059d04",
			199 => x"00000341",
			200 => x"0100e70c",
			201 => x"0a020808",
			202 => x"07051a04",
			203 => x"00000341",
			204 => x"001f0341",
			205 => x"00000341",
			206 => x"00000341",
			207 => x"00000341",
			208 => x"0e064304",
			209 => x"ff6e0375",
			210 => x"05081208",
			211 => x"0c060f04",
			212 => x"00000375",
			213 => x"ffb60375",
			214 => x"0c06de0c",
			215 => x"05082104",
			216 => x"00000375",
			217 => x"0c060f04",
			218 => x"00000375",
			219 => x"00110375",
			220 => x"00000375",
			221 => x"07054b10",
			222 => x"0c04cf04",
			223 => x"000003b9",
			224 => x"0c054308",
			225 => x"0100ad04",
			226 => x"ffea03b9",
			227 => x"000003b9",
			228 => x"000003b9",
			229 => x"0100f110",
			230 => x"0706850c",
			231 => x"0c050b04",
			232 => x"000003b9",
			233 => x"01009504",
			234 => x"000003b9",
			235 => x"002603b9",
			236 => x"000003b9",
			237 => x"000003b9",
			238 => x"03091a10",
			239 => x"0f061204",
			240 => x"00000405",
			241 => x"0d083e08",
			242 => x"0c061504",
			243 => x"ffbf0405",
			244 => x"00000405",
			245 => x"00000405",
			246 => x"0f093308",
			247 => x"06014504",
			248 => x"004c0405",
			249 => x"00000405",
			250 => x"0e0c2c0c",
			251 => x"0002e604",
			252 => x"00000405",
			253 => x"0e090704",
			254 => x"00000405",
			255 => x"ffa60405",
			256 => x"00000405",
			257 => x"0002ee20",
			258 => x"0f06b50c",
			259 => x"01009208",
			260 => x"0e059d04",
			261 => x"00000451",
			262 => x"00550451",
			263 => x"fef50451",
			264 => x"0706580c",
			265 => x"09018008",
			266 => x"0a018404",
			267 => x"00000451",
			268 => x"00990451",
			269 => x"00000451",
			270 => x"07066c04",
			271 => x"ffbf0451",
			272 => x"00160451",
			273 => x"06013b04",
			274 => x"00000451",
			275 => x"ff760451",
			276 => x"03091a1c",
			277 => x"0900f30c",
			278 => x"0e059d04",
			279 => x"000004a5",
			280 => x"0002d504",
			281 => x"002c04a5",
			282 => x"000004a5",
			283 => x"01009304",
			284 => x"000004a5",
			285 => x"0d083e08",
			286 => x"0c061504",
			287 => x"ffaf04a5",
			288 => x"000004a5",
			289 => x"000004a5",
			290 => x"0a02900c",
			291 => x"0507d704",
			292 => x"000004a5",
			293 => x"01013704",
			294 => x"003004a5",
			295 => x"000004a5",
			296 => x"000004a5",
			297 => x"0d07960c",
			298 => x"0801b004",
			299 => x"000004e9",
			300 => x"0e07dc04",
			301 => x"ffd104e9",
			302 => x"000004e9",
			303 => x"0100f814",
			304 => x"0c066610",
			305 => x"0601670c",
			306 => x"0c056304",
			307 => x"000004e9",
			308 => x"0d07d804",
			309 => x"000004e9",
			310 => x"006404e9",
			311 => x"000004e9",
			312 => x"000004e9",
			313 => x"000004e9",
			314 => x"09014f18",
			315 => x"0c052810",
			316 => x"07051a04",
			317 => x"0000053d",
			318 => x"0e059d04",
			319 => x"0000053d",
			320 => x"0002d504",
			321 => x"0025053d",
			322 => x"0000053d",
			323 => x"09014d04",
			324 => x"ff6a053d",
			325 => x"0000053d",
			326 => x"0100f110",
			327 => x"0706850c",
			328 => x"0705a504",
			329 => x"0000053d",
			330 => x"06016b04",
			331 => x"0070053d",
			332 => x"0000053d",
			333 => x"0000053d",
			334 => x"0000053d",
			335 => x"05081204",
			336 => x"ffaa0571",
			337 => x"07066c04",
			338 => x"00000571",
			339 => x"07068510",
			340 => x"02097b0c",
			341 => x"0b06fc04",
			342 => x"00000571",
			343 => x"09019004",
			344 => x"00a70571",
			345 => x"00000571",
			346 => x"00000571",
			347 => x"00000571",
			348 => x"0706721c",
			349 => x"0f061204",
			350 => x"000005ad",
			351 => x"03091a0c",
			352 => x"07065908",
			353 => x"0d083e04",
			354 => x"ffbc05ad",
			355 => x"000005ad",
			356 => x"000005ad",
			357 => x"0f093304",
			358 => x"000005ad",
			359 => x"0f097d04",
			360 => x"fffa05ad",
			361 => x"000005ad",
			362 => x"000005ad",
			363 => x"0506440c",
			364 => x"0f061a04",
			365 => x"00000601",
			366 => x"0e067104",
			367 => x"ff540601",
			368 => x"00000601",
			369 => x"09017614",
			370 => x"0e060f04",
			371 => x"00000601",
			372 => x"0d086d0c",
			373 => x"0a024108",
			374 => x"0b059904",
			375 => x"00000601",
			376 => x"00780601",
			377 => x"00000601",
			378 => x"00000601",
			379 => x"0d087408",
			380 => x"03097804",
			381 => x"ffe40601",
			382 => x"00000601",
			383 => x"00000601",
			384 => x"0002e624",
			385 => x"0507e718",
			386 => x"07058c0c",
			387 => x"02059a04",
			388 => x"0000065d",
			389 => x"0c056204",
			390 => x"002c065d",
			391 => x"0000065d",
			392 => x"0c061508",
			393 => x"0208e404",
			394 => x"ffd8065d",
			395 => x"0000065d",
			396 => x"0000065d",
			397 => x"06014208",
			398 => x"0c061004",
			399 => x"0000065d",
			400 => x"0051065d",
			401 => x"0000065d",
			402 => x"0f0b5108",
			403 => x"0a01ec04",
			404 => x"0000065d",
			405 => x"ffbd065d",
			406 => x"0000065d",
			407 => x"0506440c",
			408 => x"0c054308",
			409 => x"0600df04",
			410 => x"000006c1",
			411 => x"fe9306c1",
			412 => x"000006c1",
			413 => x"0100e410",
			414 => x"0d07a304",
			415 => x"000006c1",
			416 => x"05083e08",
			417 => x"0100cd04",
			418 => x"000006c1",
			419 => x"007906c1",
			420 => x"000006c1",
			421 => x"0d087f0c",
			422 => x"05082108",
			423 => x"09016f04",
			424 => x"000006c1",
			425 => x"ffbe06c1",
			426 => x"000006c1",
			427 => x"01013608",
			428 => x"09018004",
			429 => x"000006c1",
			430 => x"001206c1",
			431 => x"000006c1",
			432 => x"0a01e918",
			433 => x"0900f710",
			434 => x"0100970c",
			435 => x"02059a04",
			436 => x"0000072d",
			437 => x"00022e04",
			438 => x"0074072d",
			439 => x"0000072d",
			440 => x"0000072d",
			441 => x"0207cf04",
			442 => x"fff5072d",
			443 => x"0005072d",
			444 => x"0309780c",
			445 => x"0f096808",
			446 => x"0100ef04",
			447 => x"ffb7072d",
			448 => x"0000072d",
			449 => x"0000072d",
			450 => x"0c061204",
			451 => x"0000072d",
			452 => x"05083e0c",
			453 => x"0100f108",
			454 => x"07068504",
			455 => x"005a072d",
			456 => x"0000072d",
			457 => x"0000072d",
			458 => x"0000072d",
			459 => x"03091a1c",
			460 => x"0900f310",
			461 => x"00022e0c",
			462 => x"02059a04",
			463 => x"00000791",
			464 => x"0405d204",
			465 => x"00000791",
			466 => x"00320791",
			467 => x"00000791",
			468 => x"0c052804",
			469 => x"00000791",
			470 => x"0308e704",
			471 => x"ffa30791",
			472 => x"00000791",
			473 => x"09014f04",
			474 => x"00000791",
			475 => x"01013710",
			476 => x"0d082204",
			477 => x"00000791",
			478 => x"0a029008",
			479 => x"0c05d204",
			480 => x"00000791",
			481 => x"00470791",
			482 => x"00000791",
			483 => x"00000791",
			484 => x"0d08661c",
			485 => x"03062104",
			486 => x"000007dd",
			487 => x"0a01f214",
			488 => x"09018310",
			489 => x"0c050b04",
			490 => x"000007dd",
			491 => x"0f060a04",
			492 => x"000007dd",
			493 => x"0c061204",
			494 => x"006d07dd",
			495 => x"000007dd",
			496 => x"000007dd",
			497 => x"000007dd",
			498 => x"0a01f708",
			499 => x"02092804",
			500 => x"ffc207dd",
			501 => x"000007dd",
			502 => x"000007dd",
			503 => x"07061414",
			504 => x"0207800c",
			505 => x"01009208",
			506 => x"0e059d04",
			507 => x"00000851",
			508 => x"00530851",
			509 => x"00000851",
			510 => x"0c05f404",
			511 => x"ff990851",
			512 => x"00000851",
			513 => x"0c061310",
			514 => x"0901800c",
			515 => x"07067108",
			516 => x"040b8304",
			517 => x"00ab0851",
			518 => x"00000851",
			519 => x"00000851",
			520 => x"00000851",
			521 => x"03095808",
			522 => x"0507c704",
			523 => x"00000851",
			524 => x"ffdf0851",
			525 => x"0507f604",
			526 => x"00000851",
			527 => x"030cb808",
			528 => x"03096804",
			529 => x"00000851",
			530 => x"001e0851",
			531 => x"00000851",
			532 => x"0600eb0c",
			533 => x"01009708",
			534 => x"0e059d04",
			535 => x"000008b5",
			536 => x"005408b5",
			537 => x"000008b5",
			538 => x"05081218",
			539 => x"0a01d704",
			540 => x"000008b5",
			541 => x"03091a08",
			542 => x"08024104",
			543 => x"000008b5",
			544 => x"ff4f08b5",
			545 => x"08025304",
			546 => x"000008b5",
			547 => x"08029104",
			548 => x"ffea08b5",
			549 => x"000008b5",
			550 => x"0c06340c",
			551 => x"0100f808",
			552 => x"03097804",
			553 => x"000008b5",
			554 => x"006d08b5",
			555 => x"000008b5",
			556 => x"000008b5",
			557 => x"0a021d20",
			558 => x"0f062f08",
			559 => x"0c054304",
			560 => x"fff208f9",
			561 => x"000008f9",
			562 => x"0100f114",
			563 => x"07066f10",
			564 => x"0c06320c",
			565 => x"0c050b04",
			566 => x"000008f9",
			567 => x"09018704",
			568 => x"007c08f9",
			569 => x"000008f9",
			570 => x"000008f9",
			571 => x"000008f9",
			572 => x"000008f9",
			573 => x"000008f9",
			574 => x"0a01ec24",
			575 => x"03077c14",
			576 => x"0900fb10",
			577 => x"0c05250c",
			578 => x"0f05ad04",
			579 => x"0000097d",
			580 => x"0c04cd04",
			581 => x"0000097d",
			582 => x"0036097d",
			583 => x"0000097d",
			584 => x"ffb3097d",
			585 => x"0601400c",
			586 => x"0c061608",
			587 => x"09018304",
			588 => x"0087097d",
			589 => x"0000097d",
			590 => x"0000097d",
			591 => x"0000097d",
			592 => x"03097808",
			593 => x"0f094d04",
			594 => x"ff4c097d",
			595 => x"0000097d",
			596 => x"09017d0c",
			597 => x"09014f04",
			598 => x"0000097d",
			599 => x"06017004",
			600 => x"0080097d",
			601 => x"0000097d",
			602 => x"07076408",
			603 => x"0002ee04",
			604 => x"0000097d",
			605 => x"ffe0097d",
			606 => x"0000097d",
			607 => x"0506440c",
			608 => x"0c054308",
			609 => x"0600df04",
			610 => x"000009f1",
			611 => x"feb209f1",
			612 => x"000009f1",
			613 => x"0309681c",
			614 => x"0100e410",
			615 => x"03077c04",
			616 => x"000009f1",
			617 => x"0c061708",
			618 => x"0c051104",
			619 => x"000009f1",
			620 => x"002a09f1",
			621 => x"000009f1",
			622 => x"0c05f704",
			623 => x"000009f1",
			624 => x"0c063004",
			625 => x"ffad09f1",
			626 => x"000009f1",
			627 => x"0c061504",
			628 => x"000009f1",
			629 => x"0101360c",
			630 => x"0c06de08",
			631 => x"0100d404",
			632 => x"000009f1",
			633 => x"004e09f1",
			634 => x"000009f1",
			635 => x"000009f1",
			636 => x"0e087f1c",
			637 => x"0002bf18",
			638 => x"0a018410",
			639 => x"0506500c",
			640 => x"03064804",
			641 => x"00000a75",
			642 => x"0600ee04",
			643 => x"00360a75",
			644 => x"00000a75",
			645 => x"ff730a75",
			646 => x"0f070104",
			647 => x"00000a75",
			648 => x"005b0a75",
			649 => x"fec10a75",
			650 => x"0100f11c",
			651 => x"03097814",
			652 => x"0601410c",
			653 => x"0d086d08",
			654 => x"0a01ec04",
			655 => x"00d90a75",
			656 => x"00000a75",
			657 => x"00000a75",
			658 => x"0100e904",
			659 => x"00000a75",
			660 => x"ff740a75",
			661 => x"06017004",
			662 => x"00e10a75",
			663 => x"00000a75",
			664 => x"05088604",
			665 => x"ff9f0a75",
			666 => x"0a028504",
			667 => x"002e0a75",
			668 => x"00000a75",
			669 => x"0002e630",
			670 => x"0507e71c",
			671 => x"0c05f210",
			672 => x"07051804",
			673 => x"00000b09",
			674 => x"0e059d04",
			675 => x"00000b09",
			676 => x"0a01d704",
			677 => x"006e0b09",
			678 => x"00000b09",
			679 => x"04093108",
			680 => x"09017a04",
			681 => x"00000b09",
			682 => x"ff980b09",
			683 => x"00000b09",
			684 => x"0100e804",
			685 => x"00000b09",
			686 => x"0901830c",
			687 => x"0d083e04",
			688 => x"00000b09",
			689 => x"0c05f604",
			690 => x"00000b09",
			691 => x"01080b09",
			692 => x"00000b09",
			693 => x"0b06cc08",
			694 => x"0002f604",
			695 => x"00000b09",
			696 => x"feea0b09",
			697 => x"0b06ec08",
			698 => x"09018304",
			699 => x"00400b09",
			700 => x"00000b09",
			701 => x"05088608",
			702 => x"0c05f404",
			703 => x"00000b09",
			704 => x"ff9a0b09",
			705 => x"00000b09",
			706 => x"0002e628",
			707 => x"03094f24",
			708 => x"06013818",
			709 => x"07051804",
			710 => x"00000b7d",
			711 => x"0a01840c",
			712 => x"05065008",
			713 => x"0e059d04",
			714 => x"00000b7d",
			715 => x"00610b7d",
			716 => x"ffd90b7d",
			717 => x"0f077b04",
			718 => x"00000b7d",
			719 => x"00c00b7d",
			720 => x"06013e08",
			721 => x"0a01e404",
			722 => x"00000b7d",
			723 => x"ff860b7d",
			724 => x"00000b7d",
			725 => x"00ec0b7d",
			726 => x"0309a308",
			727 => x"0209ce04",
			728 => x"ff160b7d",
			729 => x"00000b7d",
			730 => x"0100f808",
			731 => x"0b072004",
			732 => x"005f0b7d",
			733 => x"00000b7d",
			734 => x"ffb20b7d",
			735 => x"0309962c",
			736 => x"08025f28",
			737 => x"0c052810",
			738 => x"0100a10c",
			739 => x"02059a04",
			740 => x"00000bf1",
			741 => x"01007804",
			742 => x"00000bf1",
			743 => x"005d0bf1",
			744 => x"00000bf1",
			745 => x"03091a10",
			746 => x"01009504",
			747 => x"00000bf1",
			748 => x"0c061508",
			749 => x"0d083e04",
			750 => x"ff8f0bf1",
			751 => x"00000bf1",
			752 => x"00000bf1",
			753 => x"0100eb04",
			754 => x"00620bf1",
			755 => x"00000bf1",
			756 => x"ffb50bf1",
			757 => x"0601960c",
			758 => x"0c061304",
			759 => x"00000bf1",
			760 => x"01013604",
			761 => x"00720bf1",
			762 => x"00000bf1",
			763 => x"00000bf1",
			764 => x"0a01f230",
			765 => x"0e072514",
			766 => x"0c04d008",
			767 => x"07050804",
			768 => x"fea10c9d",
			769 => x"051e0c9d",
			770 => x"02066104",
			771 => x"fe690c9d",
			772 => x"09010f04",
			773 => x"027d0c9d",
			774 => x"fe580c9d",
			775 => x"09018318",
			776 => x"03098714",
			777 => x"05081f0c",
			778 => x"0e07dc04",
			779 => x"01c70c9d",
			780 => x"02091104",
			781 => x"02cd0c9d",
			782 => x"03d80c9d",
			783 => x"02090c04",
			784 => x"02cb0c9d",
			785 => x"fe050c9d",
			786 => x"05150c9d",
			787 => x"fe7b0c9d",
			788 => x"0a021d14",
			789 => x"0209780c",
			790 => x"03099604",
			791 => x"fe5f0c9d",
			792 => x"07066e04",
			793 => x"02d80c9d",
			794 => x"fe760c9d",
			795 => x"0100f804",
			796 => x"05520c9d",
			797 => x"fe9a0c9d",
			798 => x"0a022308",
			799 => x"0d085804",
			800 => x"fe7b0c9d",
			801 => x"015e0c9d",
			802 => x"0d0a5f04",
			803 => x"fe5c0c9d",
			804 => x"0b086904",
			805 => x"02cf0c9d",
			806 => x"fe620c9d",
			807 => x"0409db38",
			808 => x"03096828",
			809 => x"0a01e91c",
			810 => x"0b05990c",
			811 => x"01009008",
			812 => x"0e059d04",
			813 => x"00000d19",
			814 => x"00240d19",
			815 => x"ffac0d19",
			816 => x"0100ef0c",
			817 => x"0e07dc04",
			818 => x"00000d19",
			819 => x"0f090d04",
			820 => x"008d0d19",
			821 => x"00000d19",
			822 => x"00000d19",
			823 => x"0002dd04",
			824 => x"00000d19",
			825 => x"06013904",
			826 => x"00000d19",
			827 => x"ff560d19",
			828 => x"0b07200c",
			829 => x"09019008",
			830 => x"0100f304",
			831 => x"00530d19",
			832 => x"00000d19",
			833 => x"00000d19",
			834 => x"00000d19",
			835 => x"0d0a6c04",
			836 => x"ff6d0d19",
			837 => x"00000d19",
			838 => x"0409db38",
			839 => x"07058c10",
			840 => x"07051804",
			841 => x"00000d9d",
			842 => x"01009b08",
			843 => x"0f05ad04",
			844 => x"00000d9d",
			845 => x"00820d9d",
			846 => x"00000d9d",
			847 => x"0308e708",
			848 => x"0f08bf04",
			849 => x"ff4d0d9d",
			850 => x"00000d9d",
			851 => x"06013d08",
			852 => x"0d086504",
			853 => x"00950d9d",
			854 => x"00000d9d",
			855 => x"0309580c",
			856 => x"0a01e404",
			857 => x"00000d9d",
			858 => x"07064304",
			859 => x"00000d9d",
			860 => x"ff7d0d9d",
			861 => x"09017d04",
			862 => x"00680d9d",
			863 => x"03099604",
			864 => x"ffc30d9d",
			865 => x"00000d9d",
			866 => x"0f0b5108",
			867 => x"040aa104",
			868 => x"00000d9d",
			869 => x"ff000d9d",
			870 => x"00000d9d",
			871 => x"03092e28",
			872 => x"06013520",
			873 => x"0e064308",
			874 => x"0600cd04",
			875 => x"00000e31",
			876 => x"ffa20e31",
			877 => x"0c056210",
			878 => x"0b059904",
			879 => x"00000e31",
			880 => x"0f067a04",
			881 => x"00000e31",
			882 => x"07058c04",
			883 => x"00880e31",
			884 => x"00000e31",
			885 => x"0b064b04",
			886 => x"ffb10e31",
			887 => x"00290e31",
			888 => x"0a01d704",
			889 => x"00000e31",
			890 => x"fef70e31",
			891 => x"09014f04",
			892 => x"00000e31",
			893 => x"09018318",
			894 => x"07066f0c",
			895 => x"06013e04",
			896 => x"00000e31",
			897 => x"03094004",
			898 => x"00000e31",
			899 => x"00cc0e31",
			900 => x"0b071008",
			901 => x"0b06ff04",
			902 => x"00000e31",
			903 => x"00340e31",
			904 => x"00000e31",
			905 => x"0309ef04",
			906 => x"00000e31",
			907 => x"00040e31",
			908 => x"0c050b08",
			909 => x"0600df04",
			910 => x"00000eb5",
			911 => x"ff060eb5",
			912 => x"0309ef2c",
			913 => x"08025f20",
			914 => x"0b06ff14",
			915 => x"0207cf0c",
			916 => x"0c054508",
			917 => x"0600e804",
			918 => x"00000eb5",
			919 => x"00720eb5",
			920 => x"ff810eb5",
			921 => x"0100eb04",
			922 => x"00d20eb5",
			923 => x"00000eb5",
			924 => x"03097808",
			925 => x"02090004",
			926 => x"00000eb5",
			927 => x"ffa30eb5",
			928 => x"00000eb5",
			929 => x"0309c008",
			930 => x"0209f704",
			931 => x"ff780eb5",
			932 => x"00000eb5",
			933 => x"00000eb5",
			934 => x"0601960c",
			935 => x"0c061a04",
			936 => x"00000eb5",
			937 => x"01013804",
			938 => x"00a10eb5",
			939 => x"00000eb5",
			940 => x"00000eb5",
			941 => x"07051a04",
			942 => x"ff000f39",
			943 => x"03097828",
			944 => x"0802531c",
			945 => x"0207cf10",
			946 => x"0900f308",
			947 => x"0e059d04",
			948 => x"00000f39",
			949 => x"00570f39",
			950 => x"09011304",
			951 => x"ff670f39",
			952 => x"00000f39",
			953 => x"09018008",
			954 => x"06013d04",
			955 => x"00cd0f39",
			956 => x"00000f39",
			957 => x"00000f39",
			958 => x"0c063008",
			959 => x"0c060f04",
			960 => x"00000f39",
			961 => x"ff330f39",
			962 => x"00000f39",
			963 => x"07068508",
			964 => x"09019004",
			965 => x"00cf0f39",
			966 => x"00000f39",
			967 => x"05088604",
			968 => x"ffac0f39",
			969 => x"06019608",
			970 => x"0901fa04",
			971 => x"00530f39",
			972 => x"00000f39",
			973 => x"00000f39",
			974 => x"00033540",
			975 => x"09017d18",
			976 => x"07051804",
			977 => x"00000fcd",
			978 => x"0c061710",
			979 => x"0706720c",
			980 => x"0e07dc08",
			981 => x"0f063b04",
			982 => x"00f10fcd",
			983 => x"ffe10fcd",
			984 => x"00f70fcd",
			985 => x"00000fcd",
			986 => x"00000fcd",
			987 => x"0b06fc0c",
			988 => x"0100eb04",
			989 => x"00000fcd",
			990 => x"08024e04",
			991 => x"00000fcd",
			992 => x"ff120fcd",
			993 => x"0b071010",
			994 => x"0a01f208",
			995 => x"06014104",
			996 => x"00fb0fcd",
			997 => x"00000fcd",
			998 => x"02094304",
			999 => x"ff890fcd",
			1000 => x"00000fcd",
			1001 => x"06015204",
			1002 => x"ff140fcd",
			1003 => x"0a021004",
			1004 => x"00a60fcd",
			1005 => x"00000fcd",
			1006 => x"0f0b5104",
			1007 => x"fea70fcd",
			1008 => x"06018d04",
			1009 => x"008c0fcd",
			1010 => x"00000fcd",
			1011 => x"08025a2c",
			1012 => x"0f076d1c",
			1013 => x"0f070118",
			1014 => x"0c04ea08",
			1015 => x"0e059604",
			1016 => x"ce541089",
			1017 => x"d8831089",
			1018 => x"0f06d90c",
			1019 => x"0e060f04",
			1020 => x"ce3c1089",
			1021 => x"09010604",
			1022 => x"d5e81089",
			1023 => x"ce411089",
			1024 => x"d0e71089",
			1025 => x"d4781089",
			1026 => x"09018008",
			1027 => x"0207fa04",
			1028 => x"e3991089",
			1029 => x"eff71089",
			1030 => x"0d085804",
			1031 => x"ce4f1089",
			1032 => x"e3991089",
			1033 => x"08025f0c",
			1034 => x"09017a04",
			1035 => x"e9c01089",
			1036 => x"0f093304",
			1037 => x"ce591089",
			1038 => x"d6191089",
			1039 => x"08027914",
			1040 => x"02097010",
			1041 => x"09017d08",
			1042 => x"0207f804",
			1043 => x"ce9d1089",
			1044 => x"d74c1089",
			1045 => x"0309b004",
			1046 => x"ce3e1089",
			1047 => x"d21c1089",
			1048 => x"dba91089",
			1049 => x"0a022310",
			1050 => x"040a2808",
			1051 => x"0a020804",
			1052 => x"d03c1089",
			1053 => x"ce3e1089",
			1054 => x"0802a504",
			1055 => x"d3c71089",
			1056 => x"ce651089",
			1057 => x"ce391089",
			1058 => x"00033548",
			1059 => x"06014128",
			1060 => x"0e07dc14",
			1061 => x"06010a10",
			1062 => x"0c05480c",
			1063 => x"0e059d04",
			1064 => x"ffe51135",
			1065 => x"0900f704",
			1066 => x"014c1135",
			1067 => x"00691135",
			1068 => x"ffbd1135",
			1069 => x"fe7a1135",
			1070 => x"09018310",
			1071 => x"0706850c",
			1072 => x"09017a04",
			1073 => x"01821135",
			1074 => x"07066c04",
			1075 => x"fffb1135",
			1076 => x"01af1135",
			1077 => x"00001135",
			1078 => x"ffa71135",
			1079 => x"0309a314",
			1080 => x"0209090c",
			1081 => x"05080408",
			1082 => x"08025304",
			1083 => x"00001135",
			1084 => x"feff1135",
			1085 => x"00d51135",
			1086 => x"0100eb04",
			1087 => x"00001135",
			1088 => x"fe951135",
			1089 => x"0100f808",
			1090 => x"0c063204",
			1091 => x"014a1135",
			1092 => x"00001135",
			1093 => x"00001135",
			1094 => x"0f0b5104",
			1095 => x"fe6d1135",
			1096 => x"06019d08",
			1097 => x"01014304",
			1098 => x"019b1135",
			1099 => x"00001135",
			1100 => x"fef31135",
			1101 => x"0409db44",
			1102 => x"0900fb10",
			1103 => x"00022e0c",
			1104 => x"0f05ad04",
			1105 => x"000011d1",
			1106 => x"01009b04",
			1107 => x"006d11d1",
			1108 => x"000011d1",
			1109 => x"000011d1",
			1110 => x"0308e714",
			1111 => x"0100dc08",
			1112 => x"09011b04",
			1113 => x"fff111d1",
			1114 => x"000011d1",
			1115 => x"09016304",
			1116 => x"000011d1",
			1117 => x"02088b04",
			1118 => x"ff3911d1",
			1119 => x"000011d1",
			1120 => x"06013d08",
			1121 => x"0d086504",
			1122 => x"008f11d1",
			1123 => x"000011d1",
			1124 => x"0309580c",
			1125 => x"0a01e404",
			1126 => x"000011d1",
			1127 => x"0c05d604",
			1128 => x"000011d1",
			1129 => x"ff9b11d1",
			1130 => x"0b072008",
			1131 => x"0507f504",
			1132 => x"000011d1",
			1133 => x"003a11d1",
			1134 => x"000011d1",
			1135 => x"0f0b5108",
			1136 => x"040aa104",
			1137 => x"000011d1",
			1138 => x"ff0c11d1",
			1139 => x"000011d1",
			1140 => x"0003dd40",
			1141 => x"0c05a41c",
			1142 => x"06010a14",
			1143 => x"01009b10",
			1144 => x"0e059d04",
			1145 => x"00001255",
			1146 => x"0c052a08",
			1147 => x"07051804",
			1148 => x"00001255",
			1149 => x"00441255",
			1150 => x"00001255",
			1151 => x"00001255",
			1152 => x"07061404",
			1153 => x"ff7f1255",
			1154 => x"00001255",
			1155 => x"0100e708",
			1156 => x"09014f04",
			1157 => x"00001255",
			1158 => x"00b01255",
			1159 => x"0309680c",
			1160 => x"0100e908",
			1161 => x"0507cc04",
			1162 => x"00001255",
			1163 => x"ffcf1255",
			1164 => x"00001255",
			1165 => x"0100f308",
			1166 => x"05081f04",
			1167 => x"00461255",
			1168 => x"00001255",
			1169 => x"05091b04",
			1170 => x"fff21255",
			1171 => x"00001255",
			1172 => x"ff9d1255",
			1173 => x"07051a04",
			1174 => x"feee12e9",
			1175 => x"03097828",
			1176 => x"0002dd18",
			1177 => x"0207cf10",
			1178 => x"0900f308",
			1179 => x"0e059d04",
			1180 => x"000012e9",
			1181 => x"009412e9",
			1182 => x"09011304",
			1183 => x"ff4112e9",
			1184 => x"000012e9",
			1185 => x"06013b04",
			1186 => x"00c112e9",
			1187 => x"000012e9",
			1188 => x"08025304",
			1189 => x"000012e9",
			1190 => x"0b06f004",
			1191 => x"000012e9",
			1192 => x"02094904",
			1193 => x"ff0912e9",
			1194 => x"000012e9",
			1195 => x"07068510",
			1196 => x"0901900c",
			1197 => x"0100f308",
			1198 => x"06014104",
			1199 => x"000012e9",
			1200 => x"010812e9",
			1201 => x"000012e9",
			1202 => x"000012e9",
			1203 => x"0d08da04",
			1204 => x"ff9512e9",
			1205 => x"06019608",
			1206 => x"01013b04",
			1207 => x"005112e9",
			1208 => x"000012e9",
			1209 => x"000012e9",
			1210 => x"00033554",
			1211 => x"09017d24",
			1212 => x"00020a10",
			1213 => x"0900f30c",
			1214 => x"0f05ad04",
			1215 => x"000013a5",
			1216 => x"07051a04",
			1217 => x"000013a5",
			1218 => x"017613a5",
			1219 => x"000013a5",
			1220 => x"03077c08",
			1221 => x"0900fb04",
			1222 => x"000013a5",
			1223 => x"ff3613a5",
			1224 => x"0c061708",
			1225 => x"07067204",
			1226 => x"010013a5",
			1227 => x"000013a5",
			1228 => x"000013a5",
			1229 => x"03098718",
			1230 => x"0002dd0c",
			1231 => x"0d084c08",
			1232 => x"0c05f404",
			1233 => x"000013a5",
			1234 => x"ffb413a5",
			1235 => x"00cb13a5",
			1236 => x"07068308",
			1237 => x"0c060f04",
			1238 => x"000013a5",
			1239 => x"fe8f13a5",
			1240 => x"000013a5",
			1241 => x"0c06320c",
			1242 => x"0b070104",
			1243 => x"000013a5",
			1244 => x"0100f804",
			1245 => x"00ff13a5",
			1246 => x"000013a5",
			1247 => x"06015204",
			1248 => x"ff2a13a5",
			1249 => x"0d088d04",
			1250 => x"004513a5",
			1251 => x"000013a5",
			1252 => x"0f0b5104",
			1253 => x"fe9313a5",
			1254 => x"06018d04",
			1255 => x"00af13a5",
			1256 => x"000013a5",
			1257 => x"08025f34",
			1258 => x"0e07251c",
			1259 => x"0600d908",
			1260 => x"0305b604",
			1261 => x"feb51471",
			1262 => x"063e1471",
			1263 => x"0c04ce04",
			1264 => x"00cf1471",
			1265 => x"0b059904",
			1266 => x"fe471471",
			1267 => x"09010608",
			1268 => x"0c052a04",
			1269 => x"04261471",
			1270 => x"ff191471",
			1271 => x"fe6f1471",
			1272 => x"09018314",
			1273 => x"03098710",
			1274 => x"0e09070c",
			1275 => x"0705a104",
			1276 => x"045b1471",
			1277 => x"0f082204",
			1278 => x"00e81471",
			1279 => x"033f1471",
			1280 => x"016f1471",
			1281 => x"079d1471",
			1282 => x"fe721471",
			1283 => x"0a021d20",
			1284 => x"0309ef1c",
			1285 => x"02097014",
			1286 => x"0309960c",
			1287 => x"0a01f208",
			1288 => x"0f093d04",
			1289 => x"fe891471",
			1290 => x"01621471",
			1291 => x"fe5e1471",
			1292 => x"0e094004",
			1293 => x"04331471",
			1294 => x"fe741471",
			1295 => x"02098104",
			1296 => x"04491471",
			1297 => x"fe891471",
			1298 => x"09661471",
			1299 => x"0a022308",
			1300 => x"0d085804",
			1301 => x"fe761471",
			1302 => x"01911471",
			1303 => x"0d0a5f04",
			1304 => x"fe5a1471",
			1305 => x"0b086904",
			1306 => x"039d1471",
			1307 => x"fe5f1471",
			1308 => x"0003353c",
			1309 => x"0c065038",
			1310 => x"0802411c",
			1311 => x"0207ed14",
			1312 => x"0100a10c",
			1313 => x"0e060f08",
			1314 => x"0c054304",
			1315 => x"ff7c150d",
			1316 => x"0044150d",
			1317 => x"0166150d",
			1318 => x"0c052804",
			1319 => x"0000150d",
			1320 => x"fecf150d",
			1321 => x"09017604",
			1322 => x"016b150d",
			1323 => x"0000150d",
			1324 => x"03091a08",
			1325 => x"0a01db04",
			1326 => x"0000150d",
			1327 => x"fe34150d",
			1328 => x"0a01e904",
			1329 => x"014b150d",
			1330 => x"03097808",
			1331 => x"0b070104",
			1332 => x"0035150d",
			1333 => x"fe48150d",
			1334 => x"0002ee04",
			1335 => x"0164150d",
			1336 => x"0000150d",
			1337 => x"02cc150d",
			1338 => x"0b06cc04",
			1339 => x"fe68150d",
			1340 => x"0b06dc08",
			1341 => x"0e095104",
			1342 => x"0106150d",
			1343 => x"0000150d",
			1344 => x"0509e304",
			1345 => x"feb3150d",
			1346 => x"0000150d",
			1347 => x"09018344",
			1348 => x"0e087f20",
			1349 => x"0002bf18",
			1350 => x"07058110",
			1351 => x"0c050b04",
			1352 => x"000015a1",
			1353 => x"0d066b04",
			1354 => x"000015a1",
			1355 => x"0c054804",
			1356 => x"005215a1",
			1357 => x"000015a1",
			1358 => x"0d077004",
			1359 => x"fff415a1",
			1360 => x"000015a1",
			1361 => x"08023304",
			1362 => x"000015a1",
			1363 => x"ff3415a1",
			1364 => x"07068520",
			1365 => x"07066c18",
			1366 => x"0b06f00c",
			1367 => x"07065c08",
			1368 => x"00038d04",
			1369 => x"008515a1",
			1370 => x"000015a1",
			1371 => x"000015a1",
			1372 => x"0002dd04",
			1373 => x"000015a1",
			1374 => x"0c061004",
			1375 => x"000015a1",
			1376 => x"ff7915a1",
			1377 => x"03093704",
			1378 => x"000015a1",
			1379 => x"00b815a1",
			1380 => x"000015a1",
			1381 => x"0100ed04",
			1382 => x"000015a1",
			1383 => x"ff7915a1",
			1384 => x"00022e0c",
			1385 => x"01009b08",
			1386 => x"0e059d04",
			1387 => x"0000163d",
			1388 => x"0099163d",
			1389 => x"0000163d",
			1390 => x"0706140c",
			1391 => x"06010804",
			1392 => x"0000163d",
			1393 => x"0c05b804",
			1394 => x"fed9163d",
			1395 => x"0000163d",
			1396 => x"0100e40c",
			1397 => x"06016f08",
			1398 => x"0e07dc04",
			1399 => x"0000163d",
			1400 => x"00da163d",
			1401 => x"0000163d",
			1402 => x"03092e10",
			1403 => x"06013504",
			1404 => x"0000163d",
			1405 => x"07062c04",
			1406 => x"0000163d",
			1407 => x"0c05f504",
			1408 => x"0000163d",
			1409 => x"ff2f163d",
			1410 => x"0c061610",
			1411 => x"06014208",
			1412 => x"0b06d204",
			1413 => x"0000163d",
			1414 => x"00a2163d",
			1415 => x"0d088204",
			1416 => x"fff8163d",
			1417 => x"0000163d",
			1418 => x"02090004",
			1419 => x"0000163d",
			1420 => x"0409b304",
			1421 => x"ff67163d",
			1422 => x"0000163d",
			1423 => x"0003dd40",
			1424 => x"07061614",
			1425 => x"0002cc10",
			1426 => x"0f060a04",
			1427 => x"000016c1",
			1428 => x"0100a608",
			1429 => x"0c050b04",
			1430 => x"000016c1",
			1431 => x"00b716c1",
			1432 => x"000016c1",
			1433 => x"ff2416c1",
			1434 => x"0100eb0c",
			1435 => x"07068508",
			1436 => x"0d086d04",
			1437 => x"010416c1",
			1438 => x"000016c1",
			1439 => x"000016c1",
			1440 => x"0d085704",
			1441 => x"ff7716c1",
			1442 => x"07067210",
			1443 => x"0c061608",
			1444 => x"0b071004",
			1445 => x"00a016c1",
			1446 => x"000016c1",
			1447 => x"07065704",
			1448 => x"000016c1",
			1449 => x"ff4516c1",
			1450 => x"0b06fe04",
			1451 => x"000016c1",
			1452 => x"01013604",
			1453 => x"00a416c1",
			1454 => x"000016c1",
			1455 => x"fec716c1",
			1456 => x"07051a04",
			1457 => x"fe751745",
			1458 => x"0a01d710",
			1459 => x"0207cf0c",
			1460 => x"0b05e908",
			1461 => x"02059a04",
			1462 => x"00001745",
			1463 => x"010c1745",
			1464 => x"fede1745",
			1465 => x"015b1745",
			1466 => x"0507d70c",
			1467 => x"08024104",
			1468 => x"00001745",
			1469 => x"0b06dc04",
			1470 => x"fe921745",
			1471 => x"00001745",
			1472 => x"09014f04",
			1473 => x"fed41745",
			1474 => x"07066f10",
			1475 => x"09018008",
			1476 => x"03096804",
			1477 => x"00101745",
			1478 => x"01951745",
			1479 => x"0d088204",
			1480 => x"ff701745",
			1481 => x"00501745",
			1482 => x"0309ef08",
			1483 => x"08025304",
			1484 => x"00001745",
			1485 => x"fea21745",
			1486 => x"0901ff04",
			1487 => x"01481745",
			1488 => x"ff411745",
			1489 => x"0a020860",
			1490 => x"08025330",
			1491 => x"0207cf1c",
			1492 => x"01009b10",
			1493 => x"0e05e008",
			1494 => x"0600cd04",
			1495 => x"011d1831",
			1496 => x"feaf1831",
			1497 => x"0f061204",
			1498 => x"0c9f1831",
			1499 => x"02001831",
			1500 => x"0801e404",
			1501 => x"fe721831",
			1502 => x"06010a04",
			1503 => x"00f41831",
			1504 => x"fef91831",
			1505 => x"0100ef10",
			1506 => x"0706700c",
			1507 => x"0a01e404",
			1508 => x"01ba1831",
			1509 => x"0e08e104",
			1510 => x"004a1831",
			1511 => x"022f1831",
			1512 => x"00271831",
			1513 => x"fedc1831",
			1514 => x"03097820",
			1515 => x"0a01e908",
			1516 => x"0208db04",
			1517 => x"fe651831",
			1518 => x"01df1831",
			1519 => x"06013908",
			1520 => x"0100d404",
			1521 => x"ff181831",
			1522 => x"01d71831",
			1523 => x"0f091f08",
			1524 => x"05080104",
			1525 => x"fe841831",
			1526 => x"02121831",
			1527 => x"07065804",
			1528 => x"ffdb1831",
			1529 => x"fd2f1831",
			1530 => x"0706850c",
			1531 => x"09018708",
			1532 => x"03098704",
			1533 => x"015b1831",
			1534 => x"03031831",
			1535 => x"ff101831",
			1536 => x"fe7b1831",
			1537 => x"0a023e0c",
			1538 => x"0209ce04",
			1539 => x"fe731831",
			1540 => x"01011504",
			1541 => x"03981831",
			1542 => x"ffe61831",
			1543 => x"0509e304",
			1544 => x"fe691831",
			1545 => x"0f0f4504",
			1546 => x"01901831",
			1547 => x"fe8e1831",
			1548 => x"0003244c",
			1549 => x"0e07dc1c",
			1550 => x"06010718",
			1551 => x"03062104",
			1552 => x"ff0918fd",
			1553 => x"0c054810",
			1554 => x"0c052708",
			1555 => x"0406a304",
			1556 => x"ffd118fd",
			1557 => x"00e218fd",
			1558 => x"0100a604",
			1559 => x"01b118fd",
			1560 => x"000018fd",
			1561 => x"ff1018fd",
			1562 => x"fe6918fd",
			1563 => x"06013808",
			1564 => x"0c061704",
			1565 => x"019218fd",
			1566 => x"000018fd",
			1567 => x"03092e08",
			1568 => x"0c05f504",
			1569 => x"000018fd",
			1570 => x"fe1318fd",
			1571 => x"0c061610",
			1572 => x"06014208",
			1573 => x"09018304",
			1574 => x"01b718fd",
			1575 => x"000018fd",
			1576 => x"03098704",
			1577 => x"ff6818fd",
			1578 => x"014718fd",
			1579 => x"0d087f08",
			1580 => x"0002dd04",
			1581 => x"012b18fd",
			1582 => x"fde218fd",
			1583 => x"0c062e04",
			1584 => x"01b518fd",
			1585 => x"000018fd",
			1586 => x"020b7710",
			1587 => x"0802cc0c",
			1588 => x"0d082504",
			1589 => x"febf18fd",
			1590 => x"0e095104",
			1591 => x"00f818fd",
			1592 => x"ff2f18fd",
			1593 => x"fe6918fd",
			1594 => x"0a029008",
			1595 => x"06019e04",
			1596 => x"02b918fd",
			1597 => x"000018fd",
			1598 => x"fea418fd",
			1599 => x"0a021d44",
			1600 => x"0100f340",
			1601 => x"0e07dc20",
			1602 => x"00028d1c",
			1603 => x"0c052a10",
			1604 => x"0f061208",
			1605 => x"0600cd04",
			1606 => x"01eb19b1",
			1607 => x"fe9919b1",
			1608 => x"01009b04",
			1609 => x"03cf19b1",
			1610 => x"012c19b1",
			1611 => x"0100a108",
			1612 => x"0c054604",
			1613 => x"006119b1",
			1614 => x"000019b1",
			1615 => x"fe7119b1",
			1616 => x"fdf919b1",
			1617 => x"0309a318",
			1618 => x"06013d0c",
			1619 => x"0b06ff04",
			1620 => x"01d319b1",
			1621 => x"0c061304",
			1622 => x"012c19b1",
			1623 => x"008619b1",
			1624 => x"03091a04",
			1625 => x"fc2419b1",
			1626 => x"0100eb04",
			1627 => x"01cc19b1",
			1628 => x"ffbe19b1",
			1629 => x"0b072004",
			1630 => x"03bc19b1",
			1631 => x"016c19b1",
			1632 => x"fe7319b1",
			1633 => x"0a02300c",
			1634 => x"040a6904",
			1635 => x"fe7c19b1",
			1636 => x"0802c704",
			1637 => x"040b19b1",
			1638 => x"ff6619b1",
			1639 => x"0509e304",
			1640 => x"fe6319b1",
			1641 => x"0b086904",
			1642 => x"015919b1",
			1643 => x"fe7b19b1",
			1644 => x"00030c58",
			1645 => x"0802411c",
			1646 => x"0207cf14",
			1647 => x"07058c10",
			1648 => x"0e059d04",
			1649 => x"ffbd1a95",
			1650 => x"0900f304",
			1651 => x"02081a95",
			1652 => x"0d06af04",
			1653 => x"fed21a95",
			1654 => x"01801a95",
			1655 => x"fe441a95",
			1656 => x"06013604",
			1657 => x"018f1a95",
			1658 => x"00001a95",
			1659 => x"0308ff0c",
			1660 => x"0b06cd08",
			1661 => x"02089304",
			1662 => x"fe851a95",
			1663 => x"00001a95",
			1664 => x"fcf31a95",
			1665 => x"02090010",
			1666 => x"0a01ec08",
			1667 => x"09018304",
			1668 => x"01c41a95",
			1669 => x"00001a95",
			1670 => x"03094f04",
			1671 => x"fed81a95",
			1672 => x"00001a95",
			1673 => x"03097810",
			1674 => x"0b06f008",
			1675 => x"09018004",
			1676 => x"00ac1a95",
			1677 => x"00001a95",
			1678 => x"0002ee04",
			1679 => x"fe151a95",
			1680 => x"00001a95",
			1681 => x"0d087208",
			1682 => x"0002f604",
			1683 => x"021c1a95",
			1684 => x"ffaf1a95",
			1685 => x"02095704",
			1686 => x"fee81a95",
			1687 => x"012c1a95",
			1688 => x"020b7710",
			1689 => x"0a02300c",
			1690 => x"040a2804",
			1691 => x"fecb1a95",
			1692 => x"0507c704",
			1693 => x"00001a95",
			1694 => x"00bd1a95",
			1695 => x"fe691a95",
			1696 => x"06019604",
			1697 => x"02aa1a95",
			1698 => x"08031804",
			1699 => x"00001a95",
			1700 => x"feb01a95",
			1701 => x"00030c50",
			1702 => x"08024e18",
			1703 => x"0e059d04",
			1704 => x"ff271b61",
			1705 => x"0100ef10",
			1706 => x"01009204",
			1707 => x"02911b61",
			1708 => x"0b059904",
			1709 => x"feca1b61",
			1710 => x"0f070104",
			1711 => x"00561b61",
			1712 => x"01991b61",
			1713 => x"ff9a1b61",
			1714 => x"03092208",
			1715 => x"04093104",
			1716 => x"fdda1b61",
			1717 => x"00001b61",
			1718 => x"0c061620",
			1719 => x"0f094510",
			1720 => x"08025a08",
			1721 => x"03093704",
			1722 => x"00001b61",
			1723 => x"019b1b61",
			1724 => x"0e090704",
			1725 => x"00001b61",
			1726 => x"feb91b61",
			1727 => x"0002f608",
			1728 => x"0b070104",
			1729 => x"00c71b61",
			1730 => x"02ce1b61",
			1731 => x"0c061004",
			1732 => x"00261b61",
			1733 => x"00001b61",
			1734 => x"0002dd04",
			1735 => x"01731b61",
			1736 => x"05082e04",
			1737 => x"fd5b1b61",
			1738 => x"0c062e04",
			1739 => x"01b21b61",
			1740 => x"ff1b1b61",
			1741 => x"0100d004",
			1742 => x"fe631b61",
			1743 => x"09018b0c",
			1744 => x"0d082504",
			1745 => x"fef41b61",
			1746 => x"030a8104",
			1747 => x"02831b61",
			1748 => x"ffb81b61",
			1749 => x"0509a904",
			1750 => x"fe6e1b61",
			1751 => x"01e61b61",
			1752 => x"00030c58",
			1753 => x"0c061434",
			1754 => x"0f07e314",
			1755 => x"06010a10",
			1756 => x"0c05480c",
			1757 => x"0e059d04",
			1758 => x"ffd01c45",
			1759 => x"0900f304",
			1760 => x"01ac1c45",
			1761 => x"00701c45",
			1762 => x"ff331c45",
			1763 => x"fe451c45",
			1764 => x"09017a04",
			1765 => x"018c1c45",
			1766 => x"07066c10",
			1767 => x"0c060f08",
			1768 => x"0507d704",
			1769 => x"ff471c45",
			1770 => x"013b1c45",
			1771 => x"0a01ec04",
			1772 => x"ffe71c45",
			1773 => x"fe641c45",
			1774 => x"07066f08",
			1775 => x"09018704",
			1776 => x"01f41c45",
			1777 => x"00001c45",
			1778 => x"ffce1c45",
			1779 => x"0e087f04",
			1780 => x"fe1c1c45",
			1781 => x"0f091f08",
			1782 => x"0a01ec04",
			1783 => x"01891c45",
			1784 => x"00001c45",
			1785 => x"0c061608",
			1786 => x"08025f04",
			1787 => x"01191c45",
			1788 => x"00001c45",
			1789 => x"08026f08",
			1790 => x"0c063a04",
			1791 => x"fe3d1c45",
			1792 => x"00001c45",
			1793 => x"0c063004",
			1794 => x"01221c45",
			1795 => x"00001c45",
			1796 => x"0f0b5110",
			1797 => x"0a02300c",
			1798 => x"040a2804",
			1799 => x"fedf1c45",
			1800 => x"0507c704",
			1801 => x"00001c45",
			1802 => x"00951c45",
			1803 => x"fe6b1c45",
			1804 => x"06019b08",
			1805 => x"0003d904",
			1806 => x"00001c45",
			1807 => x"023e1c45",
			1808 => x"fec41c45",
			1809 => x"0505ea04",
			1810 => x"fe781cf1",
			1811 => x"0002e634",
			1812 => x"0309582c",
			1813 => x"0c05f818",
			1814 => x"0f07e30c",
			1815 => x"06010a08",
			1816 => x"0b059904",
			1817 => x"00001cf1",
			1818 => x"00f01cf1",
			1819 => x"fefc1cf1",
			1820 => x"06014108",
			1821 => x"09018304",
			1822 => x"01631cf1",
			1823 => x"00001cf1",
			1824 => x"00001cf1",
			1825 => x"06013504",
			1826 => x"00861cf1",
			1827 => x"0507e608",
			1828 => x"09017204",
			1829 => x"00001cf1",
			1830 => x"fe601cf1",
			1831 => x"0002dd04",
			1832 => x"00d01cf1",
			1833 => x"fee91cf1",
			1834 => x"05080f04",
			1835 => x"00001cf1",
			1836 => x"017b1cf1",
			1837 => x"0309a308",
			1838 => x"0f09b104",
			1839 => x"fee21cf1",
			1840 => x"00001cf1",
			1841 => x"06016a0c",
			1842 => x"09019008",
			1843 => x"05083e04",
			1844 => x"01db1cf1",
			1845 => x"00001cf1",
			1846 => x"00001cf1",
			1847 => x"0d0a5f04",
			1848 => x"fed21cf1",
			1849 => x"0005da04",
			1850 => x"00e51cf1",
			1851 => x"00001cf1",
			1852 => x"07051a04",
			1853 => x"fe801db5",
			1854 => x"07066c38",
			1855 => x"0a01ec24",
			1856 => x"03091a1c",
			1857 => x"08024110",
			1858 => x"0207cf08",
			1859 => x"0900f304",
			1860 => x"00fe1db5",
			1861 => x"ffb31db5",
			1862 => x"09017604",
			1863 => x"01371db5",
			1864 => x"00001db5",
			1865 => x"0002c404",
			1866 => x"00001db5",
			1867 => x"0d083804",
			1868 => x"feda1db5",
			1869 => x"00001db5",
			1870 => x"09018304",
			1871 => x"012a1db5",
			1872 => x"00001db5",
			1873 => x"03097808",
			1874 => x"0f097d04",
			1875 => x"fee01db5",
			1876 => x"00001db5",
			1877 => x"02093504",
			1878 => x"00ab1db5",
			1879 => x"0c05f804",
			1880 => x"ff311db5",
			1881 => x"00001db5",
			1882 => x"07068510",
			1883 => x"0901900c",
			1884 => x"0208dd04",
			1885 => x"00001db5",
			1886 => x"0d084c04",
			1887 => x"00001db5",
			1888 => x"014c1db5",
			1889 => x"fff61db5",
			1890 => x"0d08b308",
			1891 => x"0c061104",
			1892 => x"00001db5",
			1893 => x"ff401db5",
			1894 => x"0901ff0c",
			1895 => x"08031808",
			1896 => x"06019d04",
			1897 => x"00d11db5",
			1898 => x"00001db5",
			1899 => x"00001db5",
			1900 => x"ffcb1db5",
			1901 => x"07051804",
			1902 => x"fed31e53",
			1903 => x"0a01d708",
			1904 => x"0e059d04",
			1905 => x"00001e53",
			1906 => x"00c91e53",
			1907 => x"03097828",
			1908 => x"03091a10",
			1909 => x"0002bf04",
			1910 => x"00001e53",
			1911 => x"07065908",
			1912 => x"0d083804",
			1913 => x"fef51e53",
			1914 => x"00001e53",
			1915 => x"00001e53",
			1916 => x"0d08660c",
			1917 => x"0100ed08",
			1918 => x"07068504",
			1919 => x"00c71e53",
			1920 => x"00001e53",
			1921 => x"00001e53",
			1922 => x"07068308",
			1923 => x"0c062e04",
			1924 => x"fed01e53",
			1925 => x"00001e53",
			1926 => x"00001e53",
			1927 => x"0c05f004",
			1928 => x"ffe61e53",
			1929 => x"09018308",
			1930 => x"07068504",
			1931 => x"01181e53",
			1932 => x"00001e53",
			1933 => x"0309ef08",
			1934 => x"07065604",
			1935 => x"00001e53",
			1936 => x"ffbe1e53",
			1937 => x"01013604",
			1938 => x"008e1e53",
			1939 => x"00001e53",
			1940 => x"00001e55",
			1941 => x"00001e59",
			1942 => x"00001e5d",
			1943 => x"00001e61",
			1944 => x"00001e65",
			1945 => x"00001e69",
			1946 => x"00001e6d",
			1947 => x"00001e71",
			1948 => x"0c052804",
			1949 => x"00001e85",
			1950 => x"0c065004",
			1951 => x"ffef1e85",
			1952 => x"00001e85",
			1953 => x"03098708",
			1954 => x"0305c004",
			1955 => x"00001ea1",
			1956 => x"ffe61ea1",
			1957 => x"030cb804",
			1958 => x"00051ea1",
			1959 => x"00001ea1",
			1960 => x"0002e60c",
			1961 => x"07051804",
			1962 => x"00001ebd",
			1963 => x"0405d204",
			1964 => x"00001ebd",
			1965 => x"00131ebd",
			1966 => x"00001ebd",
			1967 => x"0309870c",
			1968 => x"0900f304",
			1969 => x"00001ed9",
			1970 => x"02097804",
			1971 => x"ffbf1ed9",
			1972 => x"00001ed9",
			1973 => x"00001ed9",
			1974 => x"0508210c",
			1975 => x"07065804",
			1976 => x"00001efd",
			1977 => x"0507c704",
			1978 => x"00001efd",
			1979 => x"ffd11efd",
			1980 => x"07076804",
			1981 => x"00291efd",
			1982 => x"00001efd",
			1983 => x"0900f70c",
			1984 => x"0e059d04",
			1985 => x"00001f21",
			1986 => x"0002b704",
			1987 => x"000f1f21",
			1988 => x"00001f21",
			1989 => x"06013e04",
			1990 => x"ffba1f21",
			1991 => x"00001f21",
			1992 => x"0b06d20c",
			1993 => x"0c052804",
			1994 => x"00001f4d",
			1995 => x"0c061504",
			1996 => x"ffe61f4d",
			1997 => x"00001f4d",
			1998 => x"0100f308",
			1999 => x"07069b04",
			2000 => x"00421f4d",
			2001 => x"00001f4d",
			2002 => x"00001f4d",
			2003 => x"0309780c",
			2004 => x"07065808",
			2005 => x"07054b04",
			2006 => x"00001f79",
			2007 => x"00031f79",
			2008 => x"ffd91f79",
			2009 => x"07066c04",
			2010 => x"00001f79",
			2011 => x"07068504",
			2012 => x"000b1f79",
			2013 => x"00001f79",
			2014 => x"0a021d10",
			2015 => x"0e07dc04",
			2016 => x"00001f9d",
			2017 => x"0b072008",
			2018 => x"0100f104",
			2019 => x"005b1f9d",
			2020 => x"00001f9d",
			2021 => x"00001f9d",
			2022 => x"00001f9d",
			2023 => x"0b071010",
			2024 => x"0b066304",
			2025 => x"00001fc1",
			2026 => x"0100f108",
			2027 => x"0100cd04",
			2028 => x"00001fc1",
			2029 => x"002d1fc1",
			2030 => x"00001fc1",
			2031 => x"00001fc1",
			2032 => x"0002e610",
			2033 => x"0100ef0c",
			2034 => x"07051804",
			2035 => x"00001fe5",
			2036 => x"0405d204",
			2037 => x"00001fe5",
			2038 => x"001e1fe5",
			2039 => x"00001fe5",
			2040 => x"00001fe5",
			2041 => x"06013f10",
			2042 => x"0a01f20c",
			2043 => x"06011f04",
			2044 => x"00002011",
			2045 => x"0a01ec04",
			2046 => x"00442011",
			2047 => x"00002011",
			2048 => x"00002011",
			2049 => x"0a01e904",
			2050 => x"00002011",
			2051 => x"ffde2011",
			2052 => x"0e064304",
			2053 => x"ff5e203d",
			2054 => x"0508210c",
			2055 => x"0506a704",
			2056 => x"0000203d",
			2057 => x"05081204",
			2058 => x"ffda203d",
			2059 => x"0000203d",
			2060 => x"0509d604",
			2061 => x"0007203d",
			2062 => x"0000203d",
			2063 => x"0002c410",
			2064 => x"0d06770c",
			2065 => x"0405d204",
			2066 => x"00002071",
			2067 => x"07055d04",
			2068 => x"00202071",
			2069 => x"00002071",
			2070 => x"00002071",
			2071 => x"07066c08",
			2072 => x"0d088d04",
			2073 => x"ffd62071",
			2074 => x"00002071",
			2075 => x"00002071",
			2076 => x"06013f10",
			2077 => x"0a01f20c",
			2078 => x"0207f304",
			2079 => x"000020a5",
			2080 => x"0a01ec04",
			2081 => x"005420a5",
			2082 => x"000020a5",
			2083 => x"000020a5",
			2084 => x"020c2a08",
			2085 => x"0a01e904",
			2086 => x"000020a5",
			2087 => x"ffce20a5",
			2088 => x"000020a5",
			2089 => x"05088614",
			2090 => x"0802410c",
			2091 => x"0a018404",
			2092 => x"ffef20e1",
			2093 => x"0002cc04",
			2094 => x"000d20e1",
			2095 => x"000020e1",
			2096 => x"0a01d704",
			2097 => x"000020e1",
			2098 => x"ffb320e1",
			2099 => x"06019608",
			2100 => x"01013b04",
			2101 => x"001920e1",
			2102 => x"000020e1",
			2103 => x"000020e1",
			2104 => x"0e064308",
			2105 => x"0600d704",
			2106 => x"00002115",
			2107 => x"ffce2115",
			2108 => x"0a01ec10",
			2109 => x"0601410c",
			2110 => x"09018308",
			2111 => x"0f067a04",
			2112 => x"00002115",
			2113 => x"005e2115",
			2114 => x"00002115",
			2115 => x"00002115",
			2116 => x"00002115",
			2117 => x"0e07dc08",
			2118 => x"0801b004",
			2119 => x"00002149",
			2120 => x"ffd52149",
			2121 => x"0100f810",
			2122 => x"07069b0c",
			2123 => x"06015308",
			2124 => x"0c054c04",
			2125 => x"00002149",
			2126 => x"00602149",
			2127 => x"00002149",
			2128 => x"00002149",
			2129 => x"00002149",
			2130 => x"0002e614",
			2131 => x"0100ef10",
			2132 => x"07051804",
			2133 => x"00002175",
			2134 => x"0c061408",
			2135 => x"0405d204",
			2136 => x"00002175",
			2137 => x"00262175",
			2138 => x"00002175",
			2139 => x"00002175",
			2140 => x"00002175",
			2141 => x"0c05250c",
			2142 => x"0002a708",
			2143 => x"02059a04",
			2144 => x"000021b9",
			2145 => x"005521b9",
			2146 => x"000021b9",
			2147 => x"0706140c",
			2148 => x"0c052804",
			2149 => x"000021b9",
			2150 => x"0c05f404",
			2151 => x"ffa821b9",
			2152 => x"000021b9",
			2153 => x"06014008",
			2154 => x"0c061704",
			2155 => x"002e21b9",
			2156 => x"000021b9",
			2157 => x"000021b9",
			2158 => x"03091a18",
			2159 => x"0900f30c",
			2160 => x"0e059d04",
			2161 => x"00002205",
			2162 => x"0002d504",
			2163 => x"00272205",
			2164 => x"00002205",
			2165 => x"01009304",
			2166 => x"00002205",
			2167 => x"0d083e04",
			2168 => x"ffb72205",
			2169 => x"00002205",
			2170 => x"0a02900c",
			2171 => x"0507d704",
			2172 => x"00002205",
			2173 => x"01013704",
			2174 => x"002b2205",
			2175 => x"00002205",
			2176 => x"00002205",
			2177 => x"0c05280c",
			2178 => x"0207c208",
			2179 => x"0e059d04",
			2180 => x"00002251",
			2181 => x"00622251",
			2182 => x"00002251",
			2183 => x"03097810",
			2184 => x"0c06300c",
			2185 => x"02097808",
			2186 => x"0e092404",
			2187 => x"ff9e2251",
			2188 => x"00002251",
			2189 => x"00002251",
			2190 => x"00002251",
			2191 => x"09019008",
			2192 => x"020bbc04",
			2193 => x"00462251",
			2194 => x"00002251",
			2195 => x"00002251",
			2196 => x"09014f0c",
			2197 => x"0900f304",
			2198 => x"0000229d",
			2199 => x"01009304",
			2200 => x"0000229d",
			2201 => x"ffdc229d",
			2202 => x"0409590c",
			2203 => x"0c05f804",
			2204 => x"0000229d",
			2205 => x"0c062e04",
			2206 => x"ffdf229d",
			2207 => x"0000229d",
			2208 => x"0100f10c",
			2209 => x"0c063208",
			2210 => x"0c05d204",
			2211 => x"0000229d",
			2212 => x"0058229d",
			2213 => x"0000229d",
			2214 => x"0000229d",
			2215 => x"0507f61c",
			2216 => x"0002c40c",
			2217 => x"0f067a04",
			2218 => x"fff822f1",
			2219 => x"03075404",
			2220 => x"003322f1",
			2221 => x"000022f1",
			2222 => x"0b06fc0c",
			2223 => x"0a01db04",
			2224 => x"000022f1",
			2225 => x"0c063304",
			2226 => x"ff2c22f1",
			2227 => x"000022f1",
			2228 => x"000022f1",
			2229 => x"0601960c",
			2230 => x"01013608",
			2231 => x"0b06d204",
			2232 => x"000022f1",
			2233 => x"007322f1",
			2234 => x"000022f1",
			2235 => x"000022f1",
			2236 => x"03091a18",
			2237 => x"0900f30c",
			2238 => x"0e059d04",
			2239 => x"00002345",
			2240 => x"0002d504",
			2241 => x"00232345",
			2242 => x"00002345",
			2243 => x"07053104",
			2244 => x"00002345",
			2245 => x"0d083e04",
			2246 => x"ffbe2345",
			2247 => x"00002345",
			2248 => x"0a029010",
			2249 => x"0901ff0c",
			2250 => x"0d082204",
			2251 => x"00002345",
			2252 => x"0e08ba04",
			2253 => x"00002345",
			2254 => x"00262345",
			2255 => x"00002345",
			2256 => x"00002345",
			2257 => x"09014f14",
			2258 => x"0600d904",
			2259 => x"00002391",
			2260 => x"05064404",
			2261 => x"ff542391",
			2262 => x"07058c08",
			2263 => x"07054b04",
			2264 => x"00002391",
			2265 => x"001a2391",
			2266 => x"ffe62391",
			2267 => x"0100f110",
			2268 => x"0706850c",
			2269 => x"0705a504",
			2270 => x"00002391",
			2271 => x"06016b04",
			2272 => x"007a2391",
			2273 => x"00002391",
			2274 => x"00002391",
			2275 => x"00002391",
			2276 => x"05082118",
			2277 => x"0002dd10",
			2278 => x"0c05280c",
			2279 => x"00028d08",
			2280 => x"0c052504",
			2281 => x"001323e5",
			2282 => x"000023e5",
			2283 => x"000023e5",
			2284 => x"000023e5",
			2285 => x"08025304",
			2286 => x"000023e5",
			2287 => x"fff023e5",
			2288 => x"06019b10",
			2289 => x"0c061004",
			2290 => x"000023e5",
			2291 => x"0100de04",
			2292 => x"000023e5",
			2293 => x"01013704",
			2294 => x"003c23e5",
			2295 => x"000023e5",
			2296 => x"000023e5",
			2297 => x"08032918",
			2298 => x"0e059d04",
			2299 => x"00002419",
			2300 => x"09017d10",
			2301 => x"0706720c",
			2302 => x"07051a04",
			2303 => x"00002419",
			2304 => x"06016b04",
			2305 => x"001f2419",
			2306 => x"00002419",
			2307 => x"00002419",
			2308 => x"00002419",
			2309 => x"00002419",
			2310 => x"0002ee20",
			2311 => x"0f06b50c",
			2312 => x"01009208",
			2313 => x"0e059d04",
			2314 => x"00002465",
			2315 => x"00472465",
			2316 => x"ff0d2465",
			2317 => x"0c061610",
			2318 => x"0601420c",
			2319 => x"0100f108",
			2320 => x"0a018404",
			2321 => x"00002465",
			2322 => x"00672465",
			2323 => x"00002465",
			2324 => x"00002465",
			2325 => x"00002465",
			2326 => x"06013b04",
			2327 => x"00002465",
			2328 => x"ff842465",
			2329 => x"0507e61c",
			2330 => x"0002c40c",
			2331 => x"0f067a04",
			2332 => x"000024c1",
			2333 => x"02074b04",
			2334 => x"001a24c1",
			2335 => x"000024c1",
			2336 => x"0f09150c",
			2337 => x"0d084b08",
			2338 => x"08024104",
			2339 => x"000024c1",
			2340 => x"ff2324c1",
			2341 => x"000024c1",
			2342 => x"000024c1",
			2343 => x"06019610",
			2344 => x"0507f604",
			2345 => x"000024c1",
			2346 => x"01013608",
			2347 => x"0b06d204",
			2348 => x"000024c1",
			2349 => x"006724c1",
			2350 => x"000024c1",
			2351 => x"000024c1",
			2352 => x"03091a18",
			2353 => x"0900f30c",
			2354 => x"0406ea08",
			2355 => x"0e059d04",
			2356 => x"0000251d",
			2357 => x"0031251d",
			2358 => x"0000251d",
			2359 => x"0c052804",
			2360 => x"0000251d",
			2361 => x"0e087f04",
			2362 => x"ffa7251d",
			2363 => x"0000251d",
			2364 => x"09014f04",
			2365 => x"0000251d",
			2366 => x"0901ff10",
			2367 => x"0a02900c",
			2368 => x"0d082204",
			2369 => x"0000251d",
			2370 => x"0c05d204",
			2371 => x"0000251d",
			2372 => x"003c251d",
			2373 => x"0000251d",
			2374 => x"0000251d",
			2375 => x"09014f08",
			2376 => x"0900f304",
			2377 => x"00002571",
			2378 => x"ffe72571",
			2379 => x"04095914",
			2380 => x"0c05f804",
			2381 => x"00002571",
			2382 => x"0c062e0c",
			2383 => x"09017204",
			2384 => x"00002571",
			2385 => x"0a01db04",
			2386 => x"00002571",
			2387 => x"ffbf2571",
			2388 => x"00002571",
			2389 => x"0a02900c",
			2390 => x"0c05d204",
			2391 => x"00002571",
			2392 => x"0901ff04",
			2393 => x"00352571",
			2394 => x"00002571",
			2395 => x"00002571",
			2396 => x"0a01e918",
			2397 => x"0900f710",
			2398 => x"0100970c",
			2399 => x"02059a04",
			2400 => x"000025dd",
			2401 => x"00022e04",
			2402 => x"006425dd",
			2403 => x"000025dd",
			2404 => x"000025dd",
			2405 => x"0207cf04",
			2406 => x"fff625dd",
			2407 => x"000625dd",
			2408 => x"0309780c",
			2409 => x"0f096808",
			2410 => x"0100ef04",
			2411 => x"ffbf25dd",
			2412 => x"000025dd",
			2413 => x"000025dd",
			2414 => x"0c061204",
			2415 => x"000025dd",
			2416 => x"05083e0c",
			2417 => x"0100f108",
			2418 => x"07068504",
			2419 => x"005225dd",
			2420 => x"000025dd",
			2421 => x"000025dd",
			2422 => x"000025dd",
			2423 => x"0e092420",
			2424 => x"0c05f814",
			2425 => x"0c054304",
			2426 => x"00002641",
			2427 => x"0901830c",
			2428 => x"0900ec04",
			2429 => x"00002641",
			2430 => x"00034604",
			2431 => x"00532641",
			2432 => x"00002641",
			2433 => x"00002641",
			2434 => x"07065804",
			2435 => x"00002641",
			2436 => x"0002c404",
			2437 => x"00002641",
			2438 => x"ffaf2641",
			2439 => x"0b06d204",
			2440 => x"00002641",
			2441 => x"0a02900c",
			2442 => x"01013708",
			2443 => x"0507f604",
			2444 => x"00002641",
			2445 => x"00412641",
			2446 => x"00002641",
			2447 => x"00002641",
			2448 => x"0d08661c",
			2449 => x"03062104",
			2450 => x"0000268d",
			2451 => x"0a01f214",
			2452 => x"0c050b04",
			2453 => x"0000268d",
			2454 => x"0100f10c",
			2455 => x"07054704",
			2456 => x"0000268d",
			2457 => x"07067204",
			2458 => x"0057268d",
			2459 => x"0000268d",
			2460 => x"0000268d",
			2461 => x"0000268d",
			2462 => x"0a01f708",
			2463 => x"02092804",
			2464 => x"ffc4268d",
			2465 => x"0000268d",
			2466 => x"0000268d",
			2467 => x"03066908",
			2468 => x"0600d904",
			2469 => x"000026d1",
			2470 => x"ffd926d1",
			2471 => x"0a01ec18",
			2472 => x"06014114",
			2473 => x"0600f204",
			2474 => x"000026d1",
			2475 => x"0b059904",
			2476 => x"000026d1",
			2477 => x"09018308",
			2478 => x"0f067a04",
			2479 => x"000026d1",
			2480 => x"007e26d1",
			2481 => x"000026d1",
			2482 => x"000026d1",
			2483 => x"000026d1",
			2484 => x"05081210",
			2485 => x"06010804",
			2486 => x"00002725",
			2487 => x"0100e808",
			2488 => x"0c063004",
			2489 => x"ffdf2725",
			2490 => x"00002725",
			2491 => x"00002725",
			2492 => x"07066c04",
			2493 => x"00002725",
			2494 => x"06019b14",
			2495 => x"0c061004",
			2496 => x"00002725",
			2497 => x"0b06fc04",
			2498 => x"00002725",
			2499 => x"01013808",
			2500 => x"0100de04",
			2501 => x"00002725",
			2502 => x"00512725",
			2503 => x"00002725",
			2504 => x"00002725",
			2505 => x"0d08661c",
			2506 => x"03062104",
			2507 => x"00002761",
			2508 => x"09018314",
			2509 => x"0c050b04",
			2510 => x"00002761",
			2511 => x"0c06110c",
			2512 => x"0600f204",
			2513 => x"00002761",
			2514 => x"0f067a04",
			2515 => x"00002761",
			2516 => x"00a02761",
			2517 => x"00002761",
			2518 => x"00002761",
			2519 => x"00002761",
			2520 => x"0309962c",
			2521 => x"0a01ec20",
			2522 => x"0f062f0c",
			2523 => x"01009208",
			2524 => x"0e059d04",
			2525 => x"000027cd",
			2526 => x"000c27cd",
			2527 => x"ff4a27cd",
			2528 => x"02090010",
			2529 => x"0100ef0c",
			2530 => x"0e060f04",
			2531 => x"000027cd",
			2532 => x"0b059904",
			2533 => x"000027cd",
			2534 => x"007227cd",
			2535 => x"000027cd",
			2536 => x"000027cd",
			2537 => x"0f09b108",
			2538 => x"0b071004",
			2539 => x"ff9027cd",
			2540 => x"000027cd",
			2541 => x"000027cd",
			2542 => x"0100f808",
			2543 => x"07069b04",
			2544 => x"008d27cd",
			2545 => x"000027cd",
			2546 => x"000027cd",
			2547 => x"0506440c",
			2548 => x"0c054308",
			2549 => x"0600df04",
			2550 => x"00002841",
			2551 => x"fecd2841",
			2552 => x"00002841",
			2553 => x"0309681c",
			2554 => x"0100e410",
			2555 => x"03077c04",
			2556 => x"00002841",
			2557 => x"0c061708",
			2558 => x"0c051104",
			2559 => x"00002841",
			2560 => x"00282841",
			2561 => x"00002841",
			2562 => x"0c05f704",
			2563 => x"00002841",
			2564 => x"0c063004",
			2565 => x"ffb52841",
			2566 => x"00002841",
			2567 => x"09018710",
			2568 => x"030a810c",
			2569 => x"0c063a08",
			2570 => x"03097804",
			2571 => x"00002841",
			2572 => x"004e2841",
			2573 => x"00002841",
			2574 => x"00002841",
			2575 => x"00002841",
			2576 => x"0002e634",
			2577 => x"02088b20",
			2578 => x"0100dc18",
			2579 => x"0c050b08",
			2580 => x"0b053504",
			2581 => x"000028cd",
			2582 => x"ffee28cd",
			2583 => x"0600e804",
			2584 => x"000028cd",
			2585 => x"07054704",
			2586 => x"000028cd",
			2587 => x"07058104",
			2588 => x"008a28cd",
			2589 => x"000028cd",
			2590 => x"0308e704",
			2591 => x"ff9228cd",
			2592 => x"000028cd",
			2593 => x"0f092a0c",
			2594 => x"06014008",
			2595 => x"0100f104",
			2596 => x"009d28cd",
			2597 => x"000028cd",
			2598 => x"000028cd",
			2599 => x"07066c04",
			2600 => x"000028cd",
			2601 => x"000a28cd",
			2602 => x"0f096808",
			2603 => x"03099604",
			2604 => x"ff7328cd",
			2605 => x"000028cd",
			2606 => x"0100f308",
			2607 => x"0100d004",
			2608 => x"000028cd",
			2609 => x"004428cd",
			2610 => x"ff9c28cd",
			2611 => x"06014224",
			2612 => x"040a7b20",
			2613 => x"0c06321c",
			2614 => x"0208dd14",
			2615 => x"07058c0c",
			2616 => x"08022408",
			2617 => x"02059a04",
			2618 => x"00002929",
			2619 => x"002a2929",
			2620 => x"00002929",
			2621 => x"0c061504",
			2622 => x"ffdf2929",
			2623 => x"00002929",
			2624 => x"0100f104",
			2625 => x"004d2929",
			2626 => x"00002929",
			2627 => x"00002929",
			2628 => x"00002929",
			2629 => x"0f0b5108",
			2630 => x"08025a04",
			2631 => x"00002929",
			2632 => x"ffac2929",
			2633 => x"00002929",
			2634 => x"0b06fc2c",
			2635 => x"0a01db20",
			2636 => x"00020a10",
			2637 => x"0100970c",
			2638 => x"02059a04",
			2639 => x"000029ad",
			2640 => x"0900f304",
			2641 => x"004429ad",
			2642 => x"000029ad",
			2643 => x"000029ad",
			2644 => x"0a018404",
			2645 => x"ffdf29ad",
			2646 => x"0f070104",
			2647 => x"000029ad",
			2648 => x"06013804",
			2649 => x"001729ad",
			2650 => x"000029ad",
			2651 => x"03092e08",
			2652 => x"0002c404",
			2653 => x"000029ad",
			2654 => x"ff7929ad",
			2655 => x"000029ad",
			2656 => x"09018714",
			2657 => x"0b073310",
			2658 => x"0c061004",
			2659 => x"000029ad",
			2660 => x"0e08e104",
			2661 => x"000029ad",
			2662 => x"0c063a04",
			2663 => x"007929ad",
			2664 => x"000029ad",
			2665 => x"000029ad",
			2666 => x"000029ad",
			2667 => x"0802792c",
			2668 => x"0e06710c",
			2669 => x"0e060f04",
			2670 => x"fe712a49",
			2671 => x"0d068404",
			2672 => x"04672a49",
			2673 => x"fe932a49",
			2674 => x"0100f118",
			2675 => x"07068814",
			2676 => x"0b072010",
			2677 => x"0e092408",
			2678 => x"06014104",
			2679 => x"02282a49",
			2680 => x"00c62a49",
			2681 => x"0c061404",
			2682 => x"04e72a49",
			2683 => x"02d42a49",
			2684 => x"feb72a49",
			2685 => x"fdb22a49",
			2686 => x"0d089a04",
			2687 => x"fe6d2a49",
			2688 => x"00732a49",
			2689 => x"08029910",
			2690 => x"040a280c",
			2691 => x"0100f508",
			2692 => x"0409a004",
			2693 => x"fef32a49",
			2694 => x"011b2a49",
			2695 => x"fe752a49",
			2696 => x"03502a49",
			2697 => x"0d0a5f0c",
			2698 => x"0802b308",
			2699 => x"0802ae04",
			2700 => x"fe712a49",
			2701 => x"00002a49",
			2702 => x"fe612a49",
			2703 => x"08047204",
			2704 => x"04e02a49",
			2705 => x"fe692a49",
			2706 => x"0c05110c",
			2707 => x"0d069108",
			2708 => x"0a015104",
			2709 => x"00002ad5",
			2710 => x"fef72ad5",
			2711 => x"00002ad5",
			2712 => x"03096824",
			2713 => x"0c061018",
			2714 => x"0d07d810",
			2715 => x"0705750c",
			2716 => x"07054704",
			2717 => x"00002ad5",
			2718 => x"0c054804",
			2719 => x"003f2ad5",
			2720 => x"00002ad5",
			2721 => x"ffd12ad5",
			2722 => x"09018304",
			2723 => x"00b62ad5",
			2724 => x"00002ad5",
			2725 => x"0100e908",
			2726 => x"08024104",
			2727 => x"00002ad5",
			2728 => x"ff202ad5",
			2729 => x"00002ad5",
			2730 => x"0100f108",
			2731 => x"07068504",
			2732 => x"00b22ad5",
			2733 => x"00002ad5",
			2734 => x"0d08da04",
			2735 => x"ffd12ad5",
			2736 => x"0c06de08",
			2737 => x"0e0c3c04",
			2738 => x"00142ad5",
			2739 => x"00002ad5",
			2740 => x"00002ad5",
			2741 => x"0a01f230",
			2742 => x"0e072518",
			2743 => x"0600df08",
			2744 => x"0e059d04",
			2745 => x"fe952b89",
			2746 => x"04da2b89",
			2747 => x"0b059904",
			2748 => x"fe3f2b89",
			2749 => x"09010608",
			2750 => x"05065e04",
			2751 => x"ff292b89",
			2752 => x"03952b89",
			2753 => x"fe792b89",
			2754 => x"09018314",
			2755 => x"07068510",
			2756 => x"0309780c",
			2757 => x"05081f08",
			2758 => x"0e07dc04",
			2759 => x"017b2b89",
			2760 => x"02842b89",
			2761 => x"00602b89",
			2762 => x"04032b89",
			2763 => x"00962b89",
			2764 => x"fe812b89",
			2765 => x"0a021d18",
			2766 => x"0209780c",
			2767 => x"03099604",
			2768 => x"fe622b89",
			2769 => x"07066e04",
			2770 => x"02602b89",
			2771 => x"fe7e2b89",
			2772 => x"09019c08",
			2773 => x"0409ed04",
			2774 => x"027a2b89",
			2775 => x"04dc2b89",
			2776 => x"febe2b89",
			2777 => x"0a022308",
			2778 => x"0d085804",
			2779 => x"fe802b89",
			2780 => x"01332b89",
			2781 => x"0d0a5f04",
			2782 => x"fe5e2b89",
			2783 => x"0b086904",
			2784 => x"024f2b89",
			2785 => x"fe652b89",
			2786 => x"0506440c",
			2787 => x"04065904",
			2788 => x"00002c0d",
			2789 => x"0e067104",
			2790 => x"ff642c0d",
			2791 => x"00002c0d",
			2792 => x"0a01e910",
			2793 => x"0e060f04",
			2794 => x"00002c0d",
			2795 => x"0b059904",
			2796 => x"00002c0d",
			2797 => x"09018304",
			2798 => x"00582c0d",
			2799 => x"00002c0d",
			2800 => x"03099614",
			2801 => x"0507f404",
			2802 => x"00002c0d",
			2803 => x"0a02100c",
			2804 => x"0d084b04",
			2805 => x"00002c0d",
			2806 => x"0b071e04",
			2807 => x"ffb02c0d",
			2808 => x"00002c0d",
			2809 => x"00002c0d",
			2810 => x"0e0a4810",
			2811 => x"0507f604",
			2812 => x"00002c0d",
			2813 => x"0b075f08",
			2814 => x"0a029904",
			2815 => x"00412c0d",
			2816 => x"00002c0d",
			2817 => x"00002c0d",
			2818 => x"00002c0d",
			2819 => x"03091a28",
			2820 => x"0a01db1c",
			2821 => x"0c054814",
			2822 => x"0f067a08",
			2823 => x"0b053504",
			2824 => x"00002cb1",
			2825 => x"fff22cb1",
			2826 => x"0c04e904",
			2827 => x"00002cb1",
			2828 => x"07058c04",
			2829 => x"008d2cb1",
			2830 => x"00002cb1",
			2831 => x"0207ed04",
			2832 => x"ffc72cb1",
			2833 => x"00002cb1",
			2834 => x"08024104",
			2835 => x"00002cb1",
			2836 => x"07065904",
			2837 => x"ff0c2cb1",
			2838 => x"00002cb1",
			2839 => x"09014f04",
			2840 => x"00002cb1",
			2841 => x"0901831c",
			2842 => x"0c061a0c",
			2843 => x"06014208",
			2844 => x"04090804",
			2845 => x"00002cb1",
			2846 => x"00b52cb1",
			2847 => x"00002cb1",
			2848 => x"0d087f08",
			2849 => x"0d086504",
			2850 => x"00002cb1",
			2851 => x"ffd42cb1",
			2852 => x"0d092704",
			2853 => x"00072cb1",
			2854 => x"00002cb1",
			2855 => x"0309ef04",
			2856 => x"fffb2cb1",
			2857 => x"0d088204",
			2858 => x"00002cb1",
			2859 => x"00082cb1",
			2860 => x"0a020030",
			2861 => x"0e06710c",
			2862 => x"0e060f04",
			2863 => x"fe6c2d55",
			2864 => x"0d068404",
			2865 => x"05ba2d55",
			2866 => x"fe8a2d55",
			2867 => x"09018720",
			2868 => x"0b07201c",
			2869 => x"0e092410",
			2870 => x"0a01ec08",
			2871 => x"09011304",
			2872 => x"04c12d55",
			2873 => x"024c2d55",
			2874 => x"09017a04",
			2875 => x"024e2d55",
			2876 => x"ffd92d55",
			2877 => x"0c063208",
			2878 => x"0c061404",
			2879 => x"05b42d55",
			2880 => x"038a2d55",
			2881 => x"ff082d55",
			2882 => x"fe762d55",
			2883 => x"fe6f2d55",
			2884 => x"0a021d10",
			2885 => x"02097808",
			2886 => x"0b071e04",
			2887 => x"fe6f2d55",
			2888 => x"00702d55",
			2889 => x"0100fc04",
			2890 => x"037f2d55",
			2891 => x"febe2d55",
			2892 => x"0d0a5f0c",
			2893 => x"0a023008",
			2894 => x"0a022b04",
			2895 => x"fe6f2d55",
			2896 => x"ffe72d55",
			2897 => x"fe602d55",
			2898 => x"020fc104",
			2899 => x"06532d55",
			2900 => x"fe662d55",
			2901 => x"0c050b08",
			2902 => x"0600df04",
			2903 => x"00002de1",
			2904 => x"ff1c2de1",
			2905 => x"0d086d24",
			2906 => x"06013f18",
			2907 => x"0f07e310",
			2908 => x"0c05450c",
			2909 => x"0600e804",
			2910 => x"00002de1",
			2911 => x"07054704",
			2912 => x"00002de1",
			2913 => x"00852de1",
			2914 => x"ffa02de1",
			2915 => x"09018304",
			2916 => x"00be2de1",
			2917 => x"00002de1",
			2918 => x"05082108",
			2919 => x"0a01e904",
			2920 => x"00002de1",
			2921 => x"ffc62de1",
			2922 => x"00002de1",
			2923 => x"0309a308",
			2924 => x"0d087f04",
			2925 => x"ff4a2de1",
			2926 => x"00002de1",
			2927 => x"06019610",
			2928 => x"0c061304",
			2929 => x"00002de1",
			2930 => x"06015204",
			2931 => x"00002de1",
			2932 => x"0901f604",
			2933 => x"00ab2de1",
			2934 => x"00002de1",
			2935 => x"00002de1",
			2936 => x"07054b10",
			2937 => x"0f061204",
			2938 => x"00002e75",
			2939 => x"05067b08",
			2940 => x"0600e804",
			2941 => x"00002e75",
			2942 => x"ff6b2e75",
			2943 => x"00002e75",
			2944 => x"07065814",
			2945 => x"00030c10",
			2946 => x"0600f204",
			2947 => x"00002e75",
			2948 => x"09018008",
			2949 => x"0f067a04",
			2950 => x"00002e75",
			2951 => x"00982e75",
			2952 => x"00002e75",
			2953 => x"00002e75",
			2954 => x"07066c14",
			2955 => x"0c05f804",
			2956 => x"00002e75",
			2957 => x"040ae80c",
			2958 => x"06013504",
			2959 => x"00002e75",
			2960 => x"0d083204",
			2961 => x"00002e75",
			2962 => x"ff982e75",
			2963 => x"00002e75",
			2964 => x"0c061304",
			2965 => x"00002e75",
			2966 => x"0d085704",
			2967 => x"00002e75",
			2968 => x"06019608",
			2969 => x"05080404",
			2970 => x"00002e75",
			2971 => x"006e2e75",
			2972 => x"00002e75",
			2973 => x"0a020834",
			2974 => x"07054510",
			2975 => x"0b05930c",
			2976 => x"0b058304",
			2977 => x"fea22f21",
			2978 => x"05063504",
			2979 => x"00882f21",
			2980 => x"00002f21",
			2981 => x"fcb42f21",
			2982 => x"01009204",
			2983 => x"0b932f21",
			2984 => x"0901871c",
			2985 => x"0f06de0c",
			2986 => x"01009b08",
			2987 => x"01009904",
			2988 => x"ff792f21",
			2989 => x"00fb2f21",
			2990 => x"fe912f21",
			2991 => x"0c063208",
			2992 => x"0f096804",
			2993 => x"01912f21",
			2994 => x"03782f21",
			2995 => x"08025a04",
			2996 => x"01502f21",
			2997 => x"fe772f21",
			2998 => x"fe9a2f21",
			2999 => x"0a023e10",
			3000 => x"0209e80c",
			3001 => x"0b06cf04",
			3002 => x"fe452f21",
			3003 => x"0b06dc04",
			3004 => x"01262f21",
			3005 => x"fe882f21",
			3006 => x"03012f21",
			3007 => x"0509d30c",
			3008 => x"020b7704",
			3009 => x"fe652f21",
			3010 => x"020b8b04",
			3011 => x"05382f21",
			3012 => x"fe732f21",
			3013 => x"0c06e504",
			3014 => x"043c2f21",
			3015 => x"fe8b2f21",
			3016 => x"0802792c",
			3017 => x"0e060f04",
			3018 => x"fe752fbd",
			3019 => x"0100f120",
			3020 => x"0706881c",
			3021 => x"0e07dc10",
			3022 => x"0c052a08",
			3023 => x"0b059904",
			3024 => x"00742fbd",
			3025 => x"03fa2fbd",
			3026 => x"07057504",
			3027 => x"00202fbd",
			3028 => x"fe332fbd",
			3029 => x"0b072008",
			3030 => x"0e092404",
			3031 => x"02042fbd",
			3032 => x"03732fbd",
			3033 => x"fec22fbd",
			3034 => x"fdb42fbd",
			3035 => x"0d089a04",
			3036 => x"fe712fbd",
			3037 => x"007d2fbd",
			3038 => x"0a021d0c",
			3039 => x"0f097d04",
			3040 => x"fe7a2fbd",
			3041 => x"0100fc04",
			3042 => x"03162fbd",
			3043 => x"feb62fbd",
			3044 => x"0d0a5f10",
			3045 => x"0a02300c",
			3046 => x"0a022b04",
			3047 => x"fe772fbd",
			3048 => x"0802ae04",
			3049 => x"fec22fbd",
			3050 => x"022b2fbd",
			3051 => x"fe622fbd",
			3052 => x"0e0c7e04",
			3053 => x"03df2fbd",
			3054 => x"fe6c2fbd",
			3055 => x"08025f34",
			3056 => x"0f07011c",
			3057 => x"0e064314",
			3058 => x"0600d708",
			3059 => x"0505ea04",
			3060 => x"feb03091",
			3061 => x"08933091",
			3062 => x"0e060f04",
			3063 => x"fe643091",
			3064 => x"0d068504",
			3065 => x"032c3091",
			3066 => x"fe9f3091",
			3067 => x"0600f304",
			3068 => x"14c13091",
			3069 => x"fe773091",
			3070 => x"09018314",
			3071 => x"0b05e504",
			3072 => x"0b613091",
			3073 => x"0207ed04",
			3074 => x"fe833091",
			3075 => x"03097808",
			3076 => x"02091104",
			3077 => x"05483091",
			3078 => x"01793091",
			3079 => x"08ab3091",
			3080 => x"fe6b3091",
			3081 => x"00031a18",
			3082 => x"0100ef0c",
			3083 => x"02094308",
			3084 => x"09017d04",
			3085 => x"045e3091",
			3086 => x"feab3091",
			3087 => x"0e543091",
			3088 => x"0309b004",
			3089 => x"fe603091",
			3090 => x"0b072004",
			3091 => x"070c3091",
			3092 => x"fe8b3091",
			3093 => x"0a02230c",
			3094 => x"0d082504",
			3095 => x"fe603091",
			3096 => x"00032c04",
			3097 => x"fe893091",
			3098 => x"064a3091",
			3099 => x"0d0a5f04",
			3100 => x"fe573091",
			3101 => x"0d0a790c",
			3102 => x"0509f008",
			3103 => x"0509e304",
			3104 => x"ff663091",
			3105 => x"019e3091",
			3106 => x"feb33091",
			3107 => x"fe5b3091",
			3108 => x"0901833c",
			3109 => x"0e087f1c",
			3110 => x"0002bf18",
			3111 => x"07058110",
			3112 => x"0c050b04",
			3113 => x"00003115",
			3114 => x"0d066b04",
			3115 => x"00003115",
			3116 => x"0c054804",
			3117 => x"004e3115",
			3118 => x"00003115",
			3119 => x"0d077004",
			3120 => x"fffb3115",
			3121 => x"00003115",
			3122 => x"ff433115",
			3123 => x"0706851c",
			3124 => x"07066c14",
			3125 => x"07065a0c",
			3126 => x"0d086508",
			3127 => x"00038d04",
			3128 => x"00713115",
			3129 => x"00003115",
			3130 => x"00003115",
			3131 => x"0100eb04",
			3132 => x"00003115",
			3133 => x"ffa43115",
			3134 => x"03093704",
			3135 => x"00003115",
			3136 => x"00b03115",
			3137 => x"00003115",
			3138 => x"0100ed04",
			3139 => x"00003115",
			3140 => x"ff873115",
			3141 => x"0002e630",
			3142 => x"0100f12c",
			3143 => x"07067228",
			3144 => x"0a018418",
			3145 => x"0900f70c",
			3146 => x"0e059d04",
			3147 => x"000031a9",
			3148 => x"01009704",
			3149 => x"009431a9",
			3150 => x"000031a9",
			3151 => x"0600e604",
			3152 => x"000031a9",
			3153 => x"0a017904",
			3154 => x"ff9d31a9",
			3155 => x"000031a9",
			3156 => x"01009f04",
			3157 => x"000031a9",
			3158 => x"09018308",
			3159 => x"0f070104",
			3160 => x"000031a9",
			3161 => x"00c331a9",
			3162 => x"000031a9",
			3163 => x"000031a9",
			3164 => x"000031a9",
			3165 => x"0b06cc08",
			3166 => x"0002f604",
			3167 => x"000031a9",
			3168 => x"fed431a9",
			3169 => x"0b06ec08",
			3170 => x"09018304",
			3171 => x"003a31a9",
			3172 => x"000031a9",
			3173 => x"05088608",
			3174 => x"0c05f404",
			3175 => x"000031a9",
			3176 => x"ff7d31a9",
			3177 => x"000031a9",
			3178 => x"0003354c",
			3179 => x"06014128",
			3180 => x"0e07dc14",
			3181 => x"06010a10",
			3182 => x"0c05480c",
			3183 => x"0e059d04",
			3184 => x"ffd8325d",
			3185 => x"01009204",
			3186 => x"0180325d",
			3187 => x"0094325d",
			3188 => x"ffb0325d",
			3189 => x"fe66325d",
			3190 => x"0a01f210",
			3191 => x"0100f10c",
			3192 => x"0c05f804",
			3193 => x"018d325d",
			3194 => x"0c05f904",
			3195 => x"ff4e325d",
			3196 => x"0134325d",
			3197 => x"ffe8325d",
			3198 => x"fffc325d",
			3199 => x"0309a318",
			3200 => x"04094510",
			3201 => x"0507f508",
			3202 => x"0c05d904",
			3203 => x"0000325d",
			3204 => x"ff0d325d",
			3205 => x"0100ef04",
			3206 => x"011d325d",
			3207 => x"0000325d",
			3208 => x"0100eb04",
			3209 => x"0000325d",
			3210 => x"fea0325d",
			3211 => x"0100f808",
			3212 => x"0c063204",
			3213 => x"015a325d",
			3214 => x"0000325d",
			3215 => x"0000325d",
			3216 => x"020b7704",
			3217 => x"fe6a325d",
			3218 => x"06019d08",
			3219 => x"0100de04",
			3220 => x"0000325d",
			3221 => x"019f325d",
			3222 => x"feeb325d",
			3223 => x"0d066b08",
			3224 => x"0600d704",
			3225 => x"00003301",
			3226 => x"feb43301",
			3227 => x"0a01f220",
			3228 => x"06014114",
			3229 => x"0c050b04",
			3230 => x"00003301",
			3231 => x"03064804",
			3232 => x"00003301",
			3233 => x"0c063208",
			3234 => x"09018304",
			3235 => x"00e23301",
			3236 => x"00003301",
			3237 => x"00003301",
			3238 => x"03097808",
			3239 => x"07065a04",
			3240 => x"00003301",
			3241 => x"ff513301",
			3242 => x"00003301",
			3243 => x"0309a310",
			3244 => x"09017d0c",
			3245 => x"09015304",
			3246 => x"ff613301",
			3247 => x"020a0004",
			3248 => x"004a3301",
			3249 => x"00003301",
			3250 => x"ff233301",
			3251 => x"06015310",
			3252 => x"07069b0c",
			3253 => x"09019c08",
			3254 => x"08026f04",
			3255 => x"00003301",
			3256 => x"00e63301",
			3257 => x"00003301",
			3258 => x"00003301",
			3259 => x"0d0a6c04",
			3260 => x"ff883301",
			3261 => x"0c06fd04",
			3262 => x"00283301",
			3263 => x"00003301",
			3264 => x"0003dd4c",
			3265 => x"0a01f228",
			3266 => x"06014118",
			3267 => x"0600e808",
			3268 => x"01008a04",
			3269 => x"0000339d",
			3270 => x"ffec339d",
			3271 => x"0c050b04",
			3272 => x"0000339d",
			3273 => x"07054704",
			3274 => x"0000339d",
			3275 => x"0100f104",
			3276 => x"00e8339d",
			3277 => x"0000339d",
			3278 => x"0309780c",
			3279 => x"0100eb04",
			3280 => x"0000339d",
			3281 => x"08025304",
			3282 => x"0000339d",
			3283 => x"ff41339d",
			3284 => x"0000339d",
			3285 => x"0309a310",
			3286 => x"0209ce0c",
			3287 => x"0f093308",
			3288 => x"0f091504",
			3289 => x"ffc5339d",
			3290 => x"0000339d",
			3291 => x"ff42339d",
			3292 => x"0000339d",
			3293 => x"0100f80c",
			3294 => x"07069b08",
			3295 => x"08026f04",
			3296 => x"0000339d",
			3297 => x"00d9339d",
			3298 => x"0000339d",
			3299 => x"07073c04",
			3300 => x"ffb2339d",
			3301 => x"001e339d",
			3302 => x"febf339d",
			3303 => x"0003354c",
			3304 => x"09017d18",
			3305 => x"07051804",
			3306 => x"00003449",
			3307 => x"05081f10",
			3308 => x"0706830c",
			3309 => x"0e07dc08",
			3310 => x"0f063b04",
			3311 => x"010f3449",
			3312 => x"ffd43449",
			3313 => x"01143449",
			3314 => x"00003449",
			3315 => x"00003449",
			3316 => x"05081214",
			3317 => x"0002dd08",
			3318 => x"0d084b04",
			3319 => x"ffdc3449",
			3320 => x"00423449",
			3321 => x"04095908",
			3322 => x"07063d04",
			3323 => x"00003449",
			3324 => x"fecb3449",
			3325 => x"00003449",
			3326 => x"07067214",
			3327 => x"04097208",
			3328 => x"0d086504",
			3329 => x"00003449",
			3330 => x"ff373449",
			3331 => x"07066e08",
			3332 => x"07066c04",
			3333 => x"00003449",
			3334 => x"00853449",
			3335 => x"00003449",
			3336 => x"07069b08",
			3337 => x"0100f804",
			3338 => x"00dd3449",
			3339 => x"00003449",
			3340 => x"ffdc3449",
			3341 => x"0f0b5104",
			3342 => x"fe9d3449",
			3343 => x"06018d04",
			3344 => x"00a63449",
			3345 => x"00003449",
			3346 => x"00032444",
			3347 => x"0e07dc18",
			3348 => x"02078014",
			3349 => x"0100aa10",
			3350 => x"0e065a0c",
			3351 => x"01009208",
			3352 => x"0d063f04",
			3353 => x"ff45350d",
			3354 => x"01a9350d",
			3355 => x"fec3350d",
			3356 => x"018c350d",
			3357 => x"fee3350d",
			3358 => x"fe91350d",
			3359 => x"09017a08",
			3360 => x"0b06ff04",
			3361 => x"0196350d",
			3362 => x"ff8c350d",
			3363 => x"03092e08",
			3364 => x"0a01e404",
			3365 => x"fff5350d",
			3366 => x"fdc5350d",
			3367 => x"0c061610",
			3368 => x"0002f608",
			3369 => x"03094f04",
			3370 => x"006b350d",
			3371 => x"01d0350d",
			3372 => x"0e096204",
			3373 => x"ff0c350d",
			3374 => x"0000350d",
			3375 => x"09018004",
			3376 => x"fe2a350d",
			3377 => x"0d087f04",
			3378 => x"fffb350d",
			3379 => x"0166350d",
			3380 => x"020b7714",
			3381 => x"0802cc10",
			3382 => x"0d082504",
			3383 => x"feb5350d",
			3384 => x"0b06dc08",
			3385 => x"0e095104",
			3386 => x"016c350d",
			3387 => x"0000350d",
			3388 => x"ff10350d",
			3389 => x"fe68350d",
			3390 => x"0a029008",
			3391 => x"01016104",
			3392 => x"030d350d",
			3393 => x"0000350d",
			3394 => x"fe9b350d",
			3395 => x"08027948",
			3396 => x"09018740",
			3397 => x"0e07dc28",
			3398 => x"0c052818",
			3399 => x"0b059910",
			3400 => x"0600d908",
			3401 => x"03059904",
			3402 => x"ff3635d1",
			3403 => x"045735d1",
			3404 => x"0d068404",
			3405 => x"fe7c35d1",
			3406 => x"000035d1",
			3407 => x"0600f704",
			3408 => x"050535d1",
			3409 => x"01bd35d1",
			3410 => x"0600fb0c",
			3411 => x"07055f08",
			3412 => x"0b05b404",
			3413 => x"ff1235d1",
			3414 => x"013935d1",
			3415 => x"fe7635d1",
			3416 => x"fdea35d1",
			3417 => x"0309a314",
			3418 => x"0002e60c",
			3419 => x"09018308",
			3420 => x"0e090704",
			3421 => x"01e535d1",
			3422 => x"02f935d1",
			3423 => x"fef135d1",
			3424 => x"09017d04",
			3425 => x"011e35d1",
			3426 => x"fe4635d1",
			3427 => x"042935d1",
			3428 => x"00030c04",
			3429 => x"fe7635d1",
			3430 => x"016a35d1",
			3431 => x"0a023010",
			3432 => x"0209ce0c",
			3433 => x"0b06cf04",
			3434 => x"fe6e35d1",
			3435 => x"0e093304",
			3436 => x"018a35d1",
			3437 => x"fe8435d1",
			3438 => x"03fb35d1",
			3439 => x"0509e304",
			3440 => x"fe6135d1",
			3441 => x"0509f004",
			3442 => x"005735d1",
			3443 => x"fe7435d1",
			3444 => x"00033544",
			3445 => x"08024120",
			3446 => x"0207cf1c",
			3447 => x"0100a110",
			3448 => x"0e059d04",
			3449 => x"ff52368d",
			3450 => x"07055d08",
			3451 => x"0900f304",
			3452 => x"0212368d",
			3453 => x"00ca368d",
			3454 => x"0000368d",
			3455 => x"0c052808",
			3456 => x"07056104",
			3457 => x"ffa3368d",
			3458 => x"0035368d",
			3459 => x"feab368d",
			3460 => x"0194368d",
			3461 => x"0e088604",
			3462 => x"fd51368d",
			3463 => x"0a01e404",
			3464 => x"0193368d",
			3465 => x"02092810",
			3466 => x"0d086608",
			3467 => x"04091d04",
			3468 => x"fe92368d",
			3469 => x"00c2368d",
			3470 => x"0c063204",
			3471 => x"fddd368d",
			3472 => x"00d9368d",
			3473 => x"0a01f204",
			3474 => x"024e368d",
			3475 => x"0100f804",
			3476 => x"00af368d",
			3477 => x"fed9368d",
			3478 => x"0d0a5f14",
			3479 => x"0a023e10",
			3480 => x"0c05f804",
			3481 => x"fe5d368d",
			3482 => x"00035b08",
			3483 => x"0c061604",
			3484 => x"0000368d",
			3485 => x"ff64368d",
			3486 => x"011c368d",
			3487 => x"fe67368d",
			3488 => x"0e0ca304",
			3489 => x"01fa368d",
			3490 => x"ff0c368d",
			3491 => x"07051a04",
			3492 => x"fe723719",
			3493 => x"0002c40c",
			3494 => x"0100e908",
			3495 => x"0e059d04",
			3496 => x"00003719",
			3497 => x"01103719",
			3498 => x"00003719",
			3499 => x"0b06d20c",
			3500 => x"08024104",
			3501 => x"00003719",
			3502 => x"0f09e104",
			3503 => x"fe873719",
			3504 => x"00003719",
			3505 => x"03096810",
			3506 => x"08025308",
			3507 => x"0d083004",
			3508 => x"ffca3719",
			3509 => x"013c3719",
			3510 => x"0100e704",
			3511 => x"00013719",
			3512 => x"fe5f3719",
			3513 => x"0706850c",
			3514 => x"0100f308",
			3515 => x"0309a304",
			3516 => x"00c23719",
			3517 => x"02443719",
			3518 => x"ff103719",
			3519 => x"0d0a5f08",
			3520 => x"0c060f04",
			3521 => x"00003719",
			3522 => x"fec33719",
			3523 => x"07077c04",
			3524 => x"01113719",
			3525 => x"00003719",
			3526 => x"00033554",
			3527 => x"08024120",
			3528 => x"0f07e31c",
			3529 => x"0100a110",
			3530 => x"03064808",
			3531 => x"0600cd04",
			3532 => x"015637f5",
			3533 => x"feed37f5",
			3534 => x"07055d04",
			3535 => x"01ea37f5",
			3536 => x"000037f5",
			3537 => x"0c052808",
			3538 => x"07056104",
			3539 => x"ff8637f5",
			3540 => x"004337f5",
			3541 => x"fe9e37f5",
			3542 => x"019737f5",
			3543 => x"0308f20c",
			3544 => x"07065808",
			3545 => x"0f08bf04",
			3546 => x"fe2237f5",
			3547 => x"000037f5",
			3548 => x"fb2637f5",
			3549 => x"0a01e90c",
			3550 => x"03091a08",
			3551 => x"06013904",
			3552 => x"013e37f5",
			3553 => x"fdfc37f5",
			3554 => x"01a837f5",
			3555 => x"03098710",
			3556 => x"0b071008",
			3557 => x"0f092a04",
			3558 => x"00ba37f5",
			3559 => x"fed337f5",
			3560 => x"0c061a04",
			3561 => x"ff5937f5",
			3562 => x"fb1037f5",
			3563 => x"0c063208",
			3564 => x"09018704",
			3565 => x"021a37f5",
			3566 => x"000037f5",
			3567 => x"feb337f5",
			3568 => x"0d0a5f14",
			3569 => x"0a023e10",
			3570 => x"0c05f804",
			3571 => x"fe5237f5",
			3572 => x"0b06dc08",
			3573 => x"0b06cc04",
			3574 => x"000037f5",
			3575 => x"01a737f5",
			3576 => x"ff3d37f5",
			3577 => x"fe6737f5",
			3578 => x"07077e04",
			3579 => x"021e37f5",
			3580 => x"fef737f5",
			3581 => x"08027950",
			3582 => x"08024120",
			3583 => x"0207cf1c",
			3584 => x"0100a110",
			3585 => x"0e059d04",
			3586 => x"ff3438c9",
			3587 => x"07055d08",
			3588 => x"07051804",
			3589 => x"000038c9",
			3590 => x"01ec38c9",
			3591 => x"000038c9",
			3592 => x"0c052808",
			3593 => x"07056104",
			3594 => x"ff7938c9",
			3595 => x"005b38c9",
			3596 => x"fe8f38c9",
			3597 => x"019a38c9",
			3598 => x"02089008",
			3599 => x"0a01df04",
			3600 => x"fa6438c9",
			3601 => x"ff1038c9",
			3602 => x"0a01e90c",
			3603 => x"03091a08",
			3604 => x"09017a04",
			3605 => x"016038c9",
			3606 => x"fccb38c9",
			3607 => x"01ac38c9",
			3608 => x"02092810",
			3609 => x"0d086608",
			3610 => x"03095804",
			3611 => x"ff8c38c9",
			3612 => x"016738c9",
			3613 => x"0c063204",
			3614 => x"fd5838c9",
			3615 => x"00c638c9",
			3616 => x"0b071008",
			3617 => x"0a01f204",
			3618 => x"029d38c9",
			3619 => x"00dd38c9",
			3620 => x"feca38c9",
			3621 => x"0d0a5f14",
			3622 => x"0a023e10",
			3623 => x"0209e80c",
			3624 => x"0c061504",
			3625 => x"fe4f38c9",
			3626 => x"0c062e04",
			3627 => x"000038c9",
			3628 => x"fee838c9",
			3629 => x"01b538c9",
			3630 => x"fe6738c9",
			3631 => x"09015504",
			3632 => x"fee338c9",
			3633 => x"024a38c9",
			3634 => x"0a023e3c",
			3635 => x"09019038",
			3636 => x"0f096830",
			3637 => x"0002e620",
			3638 => x"0507f410",
			3639 => x"0c061008",
			3640 => x"03077c04",
			3641 => x"00083955",
			3642 => x"00f03955",
			3643 => x"08024104",
			3644 => x"00003955",
			3645 => x"fed33955",
			3646 => x"08025a08",
			3647 => x"03092e04",
			3648 => x"00003955",
			3649 => x"01573955",
			3650 => x"0c061204",
			3651 => x"00003955",
			3652 => x"00443955",
			3653 => x"0309960c",
			3654 => x"0507f408",
			3655 => x"0507ac04",
			3656 => x"ffa03955",
			3657 => x"00263955",
			3658 => x"fefa3955",
			3659 => x"00793955",
			3660 => x"0b072004",
			3661 => x"01883955",
			3662 => x"00003955",
			3663 => x"ff0e3955",
			3664 => x"0d0a5f04",
			3665 => x"fe7f3955",
			3666 => x"07077d04",
			3667 => x"004f3955",
			3668 => x"00003955",
			3669 => x"07051804",
			3670 => x"fedb39e9",
			3671 => x"0a01d708",
			3672 => x"0e059d04",
			3673 => x"000039e9",
			3674 => x"00b639e9",
			3675 => x"03097820",
			3676 => x"03091a0c",
			3677 => x"08024104",
			3678 => x"000039e9",
			3679 => x"0a01db04",
			3680 => x"000039e9",
			3681 => x"fef939e9",
			3682 => x"0d08660c",
			3683 => x"0100ed08",
			3684 => x"07068504",
			3685 => x"00bc39e9",
			3686 => x"000039e9",
			3687 => x"000039e9",
			3688 => x"07068304",
			3689 => x"ff1a39e9",
			3690 => x"000039e9",
			3691 => x"0b06ff08",
			3692 => x"0d086504",
			3693 => x"000039e9",
			3694 => x"ffb739e9",
			3695 => x"07069b0c",
			3696 => x"0100f808",
			3697 => x"07066c04",
			3698 => x"000039e9",
			3699 => x"010939e9",
			3700 => x"000039e9",
			3701 => x"0d0a6c04",
			3702 => x"ffd039e9",
			3703 => x"07079204",
			3704 => x"000139e9",
			3705 => x"000039e9",
			3706 => x"07051804",
			3707 => x"fea93a95",
			3708 => x"0a01d714",
			3709 => x"01009b08",
			3710 => x"0f05ad04",
			3711 => x"00003a95",
			3712 => x"00d43a95",
			3713 => x"0207cf08",
			3714 => x"0c052a04",
			3715 => x"00003a95",
			3716 => x"ff6e3a95",
			3717 => x"00d33a95",
			3718 => x"05081220",
			3719 => x"0c061414",
			3720 => x"07061504",
			3721 => x"fef53a95",
			3722 => x"0c05f508",
			3723 => x"00030c04",
			3724 => x"007c3a95",
			3725 => x"00003a95",
			3726 => x"08025a04",
			3727 => x"00003a95",
			3728 => x"ffb03a95",
			3729 => x"07065804",
			3730 => x"00003a95",
			3731 => x"0c063a04",
			3732 => x"fec13a95",
			3733 => x"00003a95",
			3734 => x"0100f114",
			3735 => x"07068510",
			3736 => x"03097808",
			3737 => x"0f092a04",
			3738 => x"00203a95",
			3739 => x"ffd33a95",
			3740 => x"08025f04",
			3741 => x"00003a95",
			3742 => x"013e3a95",
			3743 => x"00003a95",
			3744 => x"030c9908",
			3745 => x"0b070e04",
			3746 => x"00003a95",
			3747 => x"ff733a95",
			3748 => x"00143a95",
			3749 => x"07051a04",
			3750 => x"fe7a3b41",
			3751 => x"0002e638",
			3752 => x"03095830",
			3753 => x"0c05f818",
			3754 => x"0f07e30c",
			3755 => x"0c054808",
			3756 => x"0b059904",
			3757 => x"00003b41",
			3758 => x"00f93b41",
			3759 => x"ff1a3b41",
			3760 => x"0100f108",
			3761 => x"0c05f604",
			3762 => x"01613b41",
			3763 => x"00003b41",
			3764 => x"00003b41",
			3765 => x"07065808",
			3766 => x"09018004",
			3767 => x"00cb3b41",
			3768 => x"00003b41",
			3769 => x"0100e908",
			3770 => x"09017204",
			3771 => x"00003b41",
			3772 => x"fe843b41",
			3773 => x"0100ed04",
			3774 => x"00c43b41",
			3775 => x"ff593b41",
			3776 => x"05080f04",
			3777 => x"00003b41",
			3778 => x"01623b41",
			3779 => x"0309a308",
			3780 => x"0f09b104",
			3781 => x"ff093b41",
			3782 => x"00003b41",
			3783 => x"0100f80c",
			3784 => x"07068504",
			3785 => x"01b53b41",
			3786 => x"0c063204",
			3787 => x"00193b41",
			3788 => x"ffa53b41",
			3789 => x"05098a04",
			3790 => x"fed53b41",
			3791 => x"009c3b41",
			3792 => x"07051804",
			3793 => x"feb63bf5",
			3794 => x"0a01d710",
			3795 => x"0100dc0c",
			3796 => x"0f05ad04",
			3797 => x"00003bf5",
			3798 => x"0408ea04",
			3799 => x"008a3bf5",
			3800 => x"00003bf5",
			3801 => x"00003bf5",
			3802 => x"03094f1c",
			3803 => x"0706580c",
			3804 => x"0308df04",
			3805 => x"ff5f3bf5",
			3806 => x"06014104",
			3807 => x"006a3bf5",
			3808 => x"00003bf5",
			3809 => x"06013504",
			3810 => x"00003bf5",
			3811 => x"0c05f404",
			3812 => x"00003bf5",
			3813 => x"0c063004",
			3814 => x"feea3bf5",
			3815 => x"00003bf5",
			3816 => x"07066c18",
			3817 => x"0f093d0c",
			3818 => x"07065c08",
			3819 => x"09018704",
			3820 => x"008d3bf5",
			3821 => x"00003bf5",
			3822 => x"00003bf5",
			3823 => x"0d086604",
			3824 => x"00003bf5",
			3825 => x"0d088d04",
			3826 => x"fedc3bf5",
			3827 => x"00003bf5",
			3828 => x"0100f30c",
			3829 => x"07068508",
			3830 => x"0d085804",
			3831 => x"00003bf5",
			3832 => x"00cd3bf5",
			3833 => x"00003bf5",
			3834 => x"030c9904",
			3835 => x"ff963bf5",
			3836 => x"000d3bf5",
			3837 => x"07051a04",
			3838 => x"fe823c9b",
			3839 => x"0a02904c",
			3840 => x"07066c30",
			3841 => x"0a01d714",
			3842 => x"0207cf10",
			3843 => x"01009008",
			3844 => x"0c04ed04",
			3845 => x"01293c9b",
			3846 => x"00003c9b",
			3847 => x"0c052a04",
			3848 => x"00003c9b",
			3849 => x"ff303c9b",
			3850 => x"012d3c9b",
			3851 => x"03091a0c",
			3852 => x"0002c404",
			3853 => x"00003c9b",
			3854 => x"07065904",
			3855 => x"fed33c9b",
			3856 => x"00003c9b",
			3857 => x"0a01ec08",
			3858 => x"09018304",
			3859 => x"01183c9b",
			3860 => x"00003c9b",
			3861 => x"06013e04",
			3862 => x"ff323c9b",
			3863 => x"00003c9b",
			3864 => x"0706850c",
			3865 => x"0100f108",
			3866 => x"0208dd04",
			3867 => x"00003c9b",
			3868 => x"01443c9b",
			3869 => x"00003c9b",
			3870 => x"0e09c104",
			3871 => x"ff553c9b",
			3872 => x"01013908",
			3873 => x"08031804",
			3874 => x"00c83c9b",
			3875 => x"00003c9b",
			3876 => x"00003c9b",
			3877 => x"ff053c9b",
			3878 => x"00003c9d",
			3879 => x"00003ca1",
			3880 => x"00003ca5",
			3881 => x"00003ca9",
			3882 => x"00003cad",
			3883 => x"00003cb1",
			3884 => x"00003cb5",
			3885 => x"00003cb9",
			3886 => x"0801b008",
			3887 => x"0f05ad04",
			3888 => x"00003cd5",
			3889 => x"00143cd5",
			3890 => x"0f08b804",
			3891 => x"ffe83cd5",
			3892 => x"00003cd5",
			3893 => x"03098708",
			3894 => x"0305c004",
			3895 => x"00003cf1",
			3896 => x"ffeb3cf1",
			3897 => x"030cb804",
			3898 => x"00043cf1",
			3899 => x"00003cf1",
			3900 => x"01009204",
			3901 => x"00003d0d",
			3902 => x"0d087f08",
			3903 => x"05081204",
			3904 => x"ffd53d0d",
			3905 => x"00003d0d",
			3906 => x"00003d0d",
			3907 => x"0309870c",
			3908 => x"0900f304",
			3909 => x"00003d29",
			3910 => x"0d087f04",
			3911 => x"ffc83d29",
			3912 => x"00003d29",
			3913 => x"00003d29",
			3914 => x"0508210c",
			3915 => x"07065804",
			3916 => x"00003d4d",
			3917 => x"0507c704",
			3918 => x"00003d4d",
			3919 => x"ffd93d4d",
			3920 => x"07076804",
			3921 => x"00233d4d",
			3922 => x"00003d4d",
			3923 => x"0900f70c",
			3924 => x"0e059d04",
			3925 => x"00003d71",
			3926 => x"0002b704",
			3927 => x"000e3d71",
			3928 => x"00003d71",
			3929 => x"06013e04",
			3930 => x"ffc33d71",
			3931 => x"00003d71",
			3932 => x"0b06d20c",
			3933 => x"0c052804",
			3934 => x"00003d9d",
			3935 => x"0c061504",
			3936 => x"ffe83d9d",
			3937 => x"00003d9d",
			3938 => x"0100f308",
			3939 => x"07069b04",
			3940 => x"00393d9d",
			3941 => x"00003d9d",
			3942 => x"00003d9d",
			3943 => x"0a01ec0c",
			3944 => x"00021b04",
			3945 => x"00003dc9",
			3946 => x"0002f604",
			3947 => x"00323dc9",
			3948 => x"00003dc9",
			3949 => x"0a028308",
			3950 => x"0002e604",
			3951 => x"00003dc9",
			3952 => x"fff33dc9",
			3953 => x"00003dc9",
			3954 => x"0b071010",
			3955 => x"0b066304",
			3956 => x"00003ded",
			3957 => x"06014508",
			3958 => x"0100f104",
			3959 => x"003d3ded",
			3960 => x"00003ded",
			3961 => x"00003ded",
			3962 => x"00003ded",
			3963 => x"0409db10",
			3964 => x"02092004",
			3965 => x"00003e11",
			3966 => x"02097b08",
			3967 => x"08027904",
			3968 => x"003c3e11",
			3969 => x"00003e11",
			3970 => x"00003e11",
			3971 => x"00003e11",
			3972 => x"07066c10",
			3973 => x"07065804",
			3974 => x"00003e35",
			3975 => x"06013504",
			3976 => x"00003e35",
			3977 => x"0d083204",
			3978 => x"00003e35",
			3979 => x"ffcf3e35",
			3980 => x"00003e35",
			3981 => x"06013f10",
			3982 => x"0a01f20c",
			3983 => x"06011f04",
			3984 => x"00003e61",
			3985 => x"0a01ec04",
			3986 => x"00403e61",
			3987 => x"00003e61",
			3988 => x"00003e61",
			3989 => x"0a01e904",
			3990 => x"00003e61",
			3991 => x"ffe43e61",
			3992 => x"0801b00c",
			3993 => x"0900ef08",
			3994 => x"0f05ad04",
			3995 => x"00003e95",
			3996 => x"002b3e95",
			3997 => x"00003e95",
			3998 => x"0b06d204",
			3999 => x"ffda3e95",
			4000 => x"0b071004",
			4001 => x"000b3e95",
			4002 => x"0b086704",
			4003 => x"fff83e95",
			4004 => x"00003e95",
			4005 => x"0a01e910",
			4006 => x"0a014504",
			4007 => x"00003ec9",
			4008 => x"0002e608",
			4009 => x"0a01db04",
			4010 => x"00113ec9",
			4011 => x"00003ec9",
			4012 => x"00003ec9",
			4013 => x"0002dd04",
			4014 => x"00003ec9",
			4015 => x"0a028a04",
			4016 => x"fff13ec9",
			4017 => x"00003ec9",
			4018 => x"0308ff0c",
			4019 => x"0900f304",
			4020 => x"00003efd",
			4021 => x"01009304",
			4022 => x"00003efd",
			4023 => x"ffe83efd",
			4024 => x"0209810c",
			4025 => x"07068508",
			4026 => x"0100f304",
			4027 => x"003f3efd",
			4028 => x"00003efd",
			4029 => x"00003efd",
			4030 => x"00003efd",
			4031 => x"0801b00c",
			4032 => x"01009208",
			4033 => x"0e059d04",
			4034 => x"00003f39",
			4035 => x"00393f39",
			4036 => x"00003f39",
			4037 => x"0100e90c",
			4038 => x"05081208",
			4039 => x"0f09b104",
			4040 => x"ffc13f39",
			4041 => x"00003f39",
			4042 => x"00003f39",
			4043 => x"0100f104",
			4044 => x"00063f39",
			4045 => x"00003f39",
			4046 => x"09014f08",
			4047 => x"0c052804",
			4048 => x"00003f6d",
			4049 => x"ffdb3f6d",
			4050 => x"09017d10",
			4051 => x"0c06660c",
			4052 => x"0100cd04",
			4053 => x"00003f6d",
			4054 => x"0c054c04",
			4055 => x"00003f6d",
			4056 => x"00323f6d",
			4057 => x"00003f6d",
			4058 => x"00003f6d",
			4059 => x"0e07dc08",
			4060 => x"0801b004",
			4061 => x"00003fa1",
			4062 => x"ffd93fa1",
			4063 => x"0100f810",
			4064 => x"07069b0c",
			4065 => x"06015308",
			4066 => x"0c054c04",
			4067 => x"00003fa1",
			4068 => x"00543fa1",
			4069 => x"00003fa1",
			4070 => x"00003fa1",
			4071 => x"00003fa1",
			4072 => x"01009204",
			4073 => x"00003fcd",
			4074 => x"0d087f10",
			4075 => x"0c052504",
			4076 => x"00003fcd",
			4077 => x"0c062e08",
			4078 => x"07068304",
			4079 => x"ffba3fcd",
			4080 => x"00003fcd",
			4081 => x"00003fcd",
			4082 => x"00003fcd",
			4083 => x"0308ff0c",
			4084 => x"0d067704",
			4085 => x"00004009",
			4086 => x"01009004",
			4087 => x"00004009",
			4088 => x"ffeb4009",
			4089 => x"0100d004",
			4090 => x"00004009",
			4091 => x"0b07200c",
			4092 => x"0100f308",
			4093 => x"06016804",
			4094 => x"00524009",
			4095 => x"00004009",
			4096 => x"00004009",
			4097 => x"00004009",
			4098 => x"0b06d210",
			4099 => x"02078004",
			4100 => x"0000404d",
			4101 => x"0c061508",
			4102 => x"07067004",
			4103 => x"ffde404d",
			4104 => x"0000404d",
			4105 => x"0000404d",
			4106 => x"06013e04",
			4107 => x"0000404d",
			4108 => x"0101370c",
			4109 => x"0507e704",
			4110 => x"0000404d",
			4111 => x"06019d04",
			4112 => x"0036404d",
			4113 => x"0000404d",
			4114 => x"0000404d",
			4115 => x"03091a14",
			4116 => x"0900f30c",
			4117 => x"00022e08",
			4118 => x"0e059d04",
			4119 => x"00004099",
			4120 => x"002c4099",
			4121 => x"00004099",
			4122 => x"01009204",
			4123 => x"00004099",
			4124 => x"ffd14099",
			4125 => x"0100d404",
			4126 => x"00004099",
			4127 => x"0101370c",
			4128 => x"0507d704",
			4129 => x"00004099",
			4130 => x"0a029004",
			4131 => x"00364099",
			4132 => x"00004099",
			4133 => x"00004099",
			4134 => x"0e087f14",
			4135 => x"0a01d710",
			4136 => x"01009208",
			4137 => x"0e059d04",
			4138 => x"000040e5",
			4139 => x"004a40e5",
			4140 => x"0600f104",
			4141 => x"ffe640e5",
			4142 => x"000040e5",
			4143 => x"ff8040e5",
			4144 => x"09018310",
			4145 => x"0706710c",
			4146 => x"07061304",
			4147 => x"000040e5",
			4148 => x"0b06ae04",
			4149 => x"000040e5",
			4150 => x"007740e5",
			4151 => x"000040e5",
			4152 => x"000040e5",
			4153 => x"0309781c",
			4154 => x"0c052810",
			4155 => x"0e059d04",
			4156 => x"00004139",
			4157 => x"0c04cd04",
			4158 => x"00004139",
			4159 => x"0e085004",
			4160 => x"00404139",
			4161 => x"00004139",
			4162 => x"0c063008",
			4163 => x"0e092404",
			4164 => x"ffbe4139",
			4165 => x"00004139",
			4166 => x"00004139",
			4167 => x"0c06de0c",
			4168 => x"0c05d404",
			4169 => x"00004139",
			4170 => x"0e0c3c04",
			4171 => x"001b4139",
			4172 => x"00004139",
			4173 => x"00004139",
			4174 => x"07054b0c",
			4175 => x"0f05b604",
			4176 => x"0000417d",
			4177 => x"05067b04",
			4178 => x"ffbf417d",
			4179 => x"0000417d",
			4180 => x"09017d14",
			4181 => x"07069b10",
			4182 => x"0003020c",
			4183 => x"05081f08",
			4184 => x"0f062f04",
			4185 => x"0000417d",
			4186 => x"0053417d",
			4187 => x"0000417d",
			4188 => x"0000417d",
			4189 => x"0000417d",
			4190 => x"0000417d",
			4191 => x"0100cd14",
			4192 => x"0c052810",
			4193 => x"07051a04",
			4194 => x"000041c9",
			4195 => x"0e059d04",
			4196 => x"000041c9",
			4197 => x"0002d504",
			4198 => x"002241c9",
			4199 => x"000041c9",
			4200 => x"ff7a41c9",
			4201 => x"0100f110",
			4202 => x"0706850c",
			4203 => x"0d07a304",
			4204 => x"000041c9",
			4205 => x"0c058104",
			4206 => x"000041c9",
			4207 => x"006241c9",
			4208 => x"000041c9",
			4209 => x"000041c9",
			4210 => x"0b06fc1c",
			4211 => x"0002c410",
			4212 => x"0900f308",
			4213 => x"0e059d04",
			4214 => x"00004225",
			4215 => x"00424225",
			4216 => x"0e06ce04",
			4217 => x"ffef4225",
			4218 => x"00004225",
			4219 => x"03092e08",
			4220 => x"0507e604",
			4221 => x"ff7d4225",
			4222 => x"00004225",
			4223 => x"00004225",
			4224 => x"07069b10",
			4225 => x"0100f80c",
			4226 => x"0c061004",
			4227 => x"00004225",
			4228 => x"0c063404",
			4229 => x"007a4225",
			4230 => x"00004225",
			4231 => x"00004225",
			4232 => x"00004225",
			4233 => x"0100f11c",
			4234 => x"0e07dc08",
			4235 => x"06010804",
			4236 => x"00004261",
			4237 => x"fffd4261",
			4238 => x"07066f10",
			4239 => x"0901830c",
			4240 => x"0d087208",
			4241 => x"06014a04",
			4242 => x"00b44261",
			4243 => x"00004261",
			4244 => x"00004261",
			4245 => x"00004261",
			4246 => x"00004261",
			4247 => x"00004261",
			4248 => x"05081210",
			4249 => x"02078004",
			4250 => x"000042ad",
			4251 => x"0100e808",
			4252 => x"0c063004",
			4253 => x"ffd842ad",
			4254 => x"000042ad",
			4255 => x"000042ad",
			4256 => x"0b070e04",
			4257 => x"000042ad",
			4258 => x"06019b10",
			4259 => x"0c061204",
			4260 => x"000042ad",
			4261 => x"01013b08",
			4262 => x"0100de04",
			4263 => x"000042ad",
			4264 => x"005942ad",
			4265 => x"000042ad",
			4266 => x"000042ad",
			4267 => x"0c052814",
			4268 => x"0e059d04",
			4269 => x"00004309",
			4270 => x"09013d0c",
			4271 => x"0c04cd04",
			4272 => x"00004309",
			4273 => x"0900c604",
			4274 => x"00004309",
			4275 => x"004c4309",
			4276 => x"00004309",
			4277 => x"0309780c",
			4278 => x"0c063008",
			4279 => x"0e092404",
			4280 => x"ffb34309",
			4281 => x"00004309",
			4282 => x"00004309",
			4283 => x"0901900c",
			4284 => x"09014f04",
			4285 => x"00004309",
			4286 => x"0c066a04",
			4287 => x"00434309",
			4288 => x"00004309",
			4289 => x"00004309",
			4290 => x"0309781c",
			4291 => x"0a01e90c",
			4292 => x"02088b08",
			4293 => x"0507d704",
			4294 => x"fff24375",
			4295 => x"00004375",
			4296 => x"00004375",
			4297 => x"0f09680c",
			4298 => x"0002dd04",
			4299 => x"00004375",
			4300 => x"06013904",
			4301 => x"00004375",
			4302 => x"ff734375",
			4303 => x"00004375",
			4304 => x"0c062e10",
			4305 => x"0003350c",
			4306 => x"07066c04",
			4307 => x"00004375",
			4308 => x"0100f804",
			4309 => x"00784375",
			4310 => x"00004375",
			4311 => x"00004375",
			4312 => x"0b086608",
			4313 => x"07065804",
			4314 => x"00004375",
			4315 => x"ffdb4375",
			4316 => x"00004375",
			4317 => x"05082124",
			4318 => x"0002dd14",
			4319 => x"0f062f08",
			4320 => x"01008204",
			4321 => x"000043e1",
			4322 => x"ffcb43e1",
			4323 => x"0100aa08",
			4324 => x"0b059904",
			4325 => x"000043e1",
			4326 => x"005643e1",
			4327 => x"000043e1",
			4328 => x"0d087f0c",
			4329 => x"0507ea04",
			4330 => x"000043e1",
			4331 => x"0d083e04",
			4332 => x"000043e1",
			4333 => x"ff9443e1",
			4334 => x"000043e1",
			4335 => x"0a029010",
			4336 => x"0b06fe04",
			4337 => x"000043e1",
			4338 => x"07066c04",
			4339 => x"000043e1",
			4340 => x"0901f604",
			4341 => x"003f43e1",
			4342 => x"000043e1",
			4343 => x"000043e1",
			4344 => x"0507e61c",
			4345 => x"0002c40c",
			4346 => x"0f067a04",
			4347 => x"00004445",
			4348 => x"0f07d504",
			4349 => x"000f4445",
			4350 => x"00004445",
			4351 => x"0f09150c",
			4352 => x"0d084b08",
			4353 => x"08024104",
			4354 => x"00004445",
			4355 => x"ff314445",
			4356 => x"00004445",
			4357 => x"00004445",
			4358 => x"0a029014",
			4359 => x"01013610",
			4360 => x"0c05d404",
			4361 => x"00004445",
			4362 => x"03091a04",
			4363 => x"00004445",
			4364 => x"06019604",
			4365 => x"005a4445",
			4366 => x"00004445",
			4367 => x"00004445",
			4368 => x"00004445",
			4369 => x"0508211c",
			4370 => x"0c060f10",
			4371 => x"0003020c",
			4372 => x"0a016604",
			4373 => x"000044a9",
			4374 => x"0c050b04",
			4375 => x"000044a9",
			4376 => x"005044a9",
			4377 => x"000044a9",
			4378 => x"08024104",
			4379 => x"000044a9",
			4380 => x"00033e04",
			4381 => x"ffe644a9",
			4382 => x"000044a9",
			4383 => x"06019b14",
			4384 => x"0c061004",
			4385 => x"000044a9",
			4386 => x"0901ff0c",
			4387 => x"0a029308",
			4388 => x"0b06fe04",
			4389 => x"000044a9",
			4390 => x"003b44a9",
			4391 => x"000044a9",
			4392 => x"000044a9",
			4393 => x"000044a9",
			4394 => x"0706141c",
			4395 => x"02078014",
			4396 => x"01009210",
			4397 => x"02059a04",
			4398 => x"0000451d",
			4399 => x"0c04cd04",
			4400 => x"0000451d",
			4401 => x"0405d204",
			4402 => x"0000451d",
			4403 => x"005f451d",
			4404 => x"0000451d",
			4405 => x"0c05f404",
			4406 => x"ff8f451d",
			4407 => x"0000451d",
			4408 => x"03096814",
			4409 => x"0c060f08",
			4410 => x"0100eb04",
			4411 => x"004e451d",
			4412 => x"0000451d",
			4413 => x"08024104",
			4414 => x"0000451d",
			4415 => x"07064304",
			4416 => x"0000451d",
			4417 => x"ffc4451d",
			4418 => x"09018308",
			4419 => x"07068504",
			4420 => x"009a451d",
			4421 => x"0000451d",
			4422 => x"0000451d",
			4423 => x"03066908",
			4424 => x"0600d904",
			4425 => x"00004561",
			4426 => x"ffdf4561",
			4427 => x"0a01ec18",
			4428 => x"06014114",
			4429 => x"0600f204",
			4430 => x"00004561",
			4431 => x"0b059904",
			4432 => x"00004561",
			4433 => x"0f067a04",
			4434 => x"00004561",
			4435 => x"0100f104",
			4436 => x"00714561",
			4437 => x"00004561",
			4438 => x"00004561",
			4439 => x"00004561",
			4440 => x"0a01e914",
			4441 => x"0900f70c",
			4442 => x"01009708",
			4443 => x"0e059d04",
			4444 => x"000045cd",
			4445 => x"005545cd",
			4446 => x"000045cd",
			4447 => x"0207cf04",
			4448 => x"fff745cd",
			4449 => x"000645cd",
			4450 => x"0309780c",
			4451 => x"0100ef08",
			4452 => x"02097804",
			4453 => x"ffc645cd",
			4454 => x"000045cd",
			4455 => x"000045cd",
			4456 => x"0c061204",
			4457 => x"000045cd",
			4458 => x"01013610",
			4459 => x"07065b04",
			4460 => x"000045cd",
			4461 => x"0100d404",
			4462 => x"000045cd",
			4463 => x"05083e04",
			4464 => x"004e45cd",
			4465 => x"000045cd",
			4466 => x"000045cd",
			4467 => x"05082120",
			4468 => x"0002dd18",
			4469 => x"0c061414",
			4470 => x"0a016604",
			4471 => x"00004631",
			4472 => x"0c050b04",
			4473 => x"00004631",
			4474 => x"0a01ec08",
			4475 => x"0c061004",
			4476 => x"00314631",
			4477 => x"00004631",
			4478 => x"00004631",
			4479 => x"00004631",
			4480 => x"0a01e904",
			4481 => x"00004631",
			4482 => x"ffea4631",
			4483 => x"0a029010",
			4484 => x"0c061004",
			4485 => x"00004631",
			4486 => x"01013708",
			4487 => x"07066c04",
			4488 => x"00004631",
			4489 => x"00404631",
			4490 => x"00004631",
			4491 => x"00004631",
			4492 => x"0002ee2c",
			4493 => x"0e06710c",
			4494 => x"01009208",
			4495 => x"0e059d04",
			4496 => x"00004695",
			4497 => x"00494695",
			4498 => x"fee64695",
			4499 => x"0c061614",
			4500 => x"06014210",
			4501 => x"0600f604",
			4502 => x"00004695",
			4503 => x"09018308",
			4504 => x"0e06ce04",
			4505 => x"00004695",
			4506 => x"00764695",
			4507 => x"00004695",
			4508 => x"00004695",
			4509 => x"02090004",
			4510 => x"00004695",
			4511 => x"02091b04",
			4512 => x"ffde4695",
			4513 => x"00004695",
			4514 => x"06013b04",
			4515 => x"00004695",
			4516 => x"ff664695",
			4517 => x"0309962c",
			4518 => x"08025f24",
			4519 => x"0c052810",
			4520 => x"0100a10c",
			4521 => x"0f05ad04",
			4522 => x"00004709",
			4523 => x"01007804",
			4524 => x"00004709",
			4525 => x"004f4709",
			4526 => x"00004709",
			4527 => x"03091a0c",
			4528 => x"01009504",
			4529 => x"00004709",
			4530 => x"0801cb04",
			4531 => x"ff6d4709",
			4532 => x"00004709",
			4533 => x"0100eb04",
			4534 => x"005e4709",
			4535 => x"00004709",
			4536 => x"0f09e104",
			4537 => x"ffbc4709",
			4538 => x"00004709",
			4539 => x"0601960c",
			4540 => x"0c061304",
			4541 => x"00004709",
			4542 => x"01013604",
			4543 => x"00674709",
			4544 => x"00004709",
			4545 => x"00004709",
			4546 => x"0600eb10",
			4547 => x"0100970c",
			4548 => x"0e059d04",
			4549 => x"00004785",
			4550 => x"07051a04",
			4551 => x"00004785",
			4552 => x"00614785",
			4553 => x"00004785",
			4554 => x"0508121c",
			4555 => x"08024104",
			4556 => x"00004785",
			4557 => x"03091a08",
			4558 => x"0a01d704",
			4559 => x"00004785",
			4560 => x"ff424785",
			4561 => x"0a01e904",
			4562 => x"00004785",
			4563 => x"0e08f004",
			4564 => x"00004785",
			4565 => x"0209f704",
			4566 => x"ffc94785",
			4567 => x"00004785",
			4568 => x"07066f0c",
			4569 => x"0100f108",
			4570 => x"08025a04",
			4571 => x"00004785",
			4572 => x"008c4785",
			4573 => x"00004785",
			4574 => x"0d08da04",
			4575 => x"fff94785",
			4576 => x"00004785",
			4577 => x"0b06fc30",
			4578 => x"0a01db20",
			4579 => x"00020a10",
			4580 => x"0100970c",
			4581 => x"02059a04",
			4582 => x"00004809",
			4583 => x"07051a04",
			4584 => x"00004809",
			4585 => x"003d4809",
			4586 => x"00004809",
			4587 => x"0a018404",
			4588 => x"ffe34809",
			4589 => x"0f070104",
			4590 => x"00004809",
			4591 => x"06013804",
			4592 => x"00194809",
			4593 => x"00004809",
			4594 => x"03092e0c",
			4595 => x"0002c404",
			4596 => x"00004809",
			4597 => x"0507e604",
			4598 => x"ff814809",
			4599 => x"00004809",
			4600 => x"00004809",
			4601 => x"07069b10",
			4602 => x"0100f80c",
			4603 => x"0c061004",
			4604 => x"00004809",
			4605 => x"0c063204",
			4606 => x"00764809",
			4607 => x"00004809",
			4608 => x"00004809",
			4609 => x"00004809",
			4610 => x"0002e634",
			4611 => x"0507e724",
			4612 => x"0100dc10",
			4613 => x"0c05f20c",
			4614 => x"02059a04",
			4615 => x"00004885",
			4616 => x"0a01d704",
			4617 => x"00324885",
			4618 => x"00004885",
			4619 => x"00004885",
			4620 => x"09016304",
			4621 => x"00004885",
			4622 => x"0208e90c",
			4623 => x"0c059f04",
			4624 => x"00004885",
			4625 => x"0c061504",
			4626 => x"ffc94885",
			4627 => x"00004885",
			4628 => x"00004885",
			4629 => x"05081f0c",
			4630 => x"0c05f604",
			4631 => x"00004885",
			4632 => x"09018304",
			4633 => x"00634885",
			4634 => x"00004885",
			4635 => x"00004885",
			4636 => x"0f0b5108",
			4637 => x"0a01ec04",
			4638 => x"00004885",
			4639 => x"ffb74885",
			4640 => x"00004885",
			4641 => x"0507f634",
			4642 => x"06013520",
			4643 => x"0e064308",
			4644 => x"0600cd04",
			4645 => x"00004929",
			4646 => x"ffb04929",
			4647 => x"0c056210",
			4648 => x"0b059904",
			4649 => x"00004929",
			4650 => x"0f067a04",
			4651 => x"00004929",
			4652 => x"07058c04",
			4653 => x"007e4929",
			4654 => x"00004929",
			4655 => x"05075604",
			4656 => x"ffbc4929",
			4657 => x"00344929",
			4658 => x"03092e10",
			4659 => x"0002bf04",
			4660 => x"00004929",
			4661 => x"0507e608",
			4662 => x"0d083e04",
			4663 => x"ff004929",
			4664 => x"00004929",
			4665 => x"00004929",
			4666 => x"00004929",
			4667 => x"06013e0c",
			4668 => x"02090004",
			4669 => x"00374929",
			4670 => x"09018004",
			4671 => x"ffb84929",
			4672 => x"00004929",
			4673 => x"07066f08",
			4674 => x"09018304",
			4675 => x"00e64929",
			4676 => x"00004929",
			4677 => x"0309ef04",
			4678 => x"fff74929",
			4679 => x"030cb804",
			4680 => x"00194929",
			4681 => x"00004929",
			4682 => x"0e087f1c",
			4683 => x"0002bf18",
			4684 => x"0a018410",
			4685 => x"0506500c",
			4686 => x"03064804",
			4687 => x"000049c5",
			4688 => x"0600ee04",
			4689 => x"003d49c5",
			4690 => x"000049c5",
			4691 => x"ff6349c5",
			4692 => x"0f070104",
			4693 => x"000049c5",
			4694 => x"005b49c5",
			4695 => x"feb649c5",
			4696 => x"09018324",
			4697 => x"0c061a0c",
			4698 => x"06014208",
			4699 => x"0308ff04",
			4700 => x"000049c5",
			4701 => x"00cb49c5",
			4702 => x"000049c5",
			4703 => x"0e09240c",
			4704 => x"0002dd04",
			4705 => x"002f49c5",
			4706 => x"0b071e04",
			4707 => x"ff3d49c5",
			4708 => x"000049c5",
			4709 => x"09015c04",
			4710 => x"000049c5",
			4711 => x"0c063a04",
			4712 => x"009849c5",
			4713 => x"000049c5",
			4714 => x"0d088204",
			4715 => x"ffb449c5",
			4716 => x"0309a304",
			4717 => x"000049c5",
			4718 => x"05082104",
			4719 => x"000049c5",
			4720 => x"003049c5",
			4721 => x"0802cc34",
			4722 => x"0100f12c",
			4723 => x"03098720",
			4724 => x"0002e614",
			4725 => x"0f092a10",
			4726 => x"0308ff08",
			4727 => x"08024104",
			4728 => x"006f4a41",
			4729 => x"ff454a41",
			4730 => x"09018304",
			4731 => x"01284a41",
			4732 => x"00004a41",
			4733 => x"00004a41",
			4734 => x"0100e908",
			4735 => x"0b06af04",
			4736 => x"ffbd4a41",
			4737 => x"00404a41",
			4738 => x"ff144a41",
			4739 => x"02093004",
			4740 => x"00004a41",
			4741 => x"07068504",
			4742 => x"01634a41",
			4743 => x"00004a41",
			4744 => x"09018704",
			4745 => x"00004a41",
			4746 => x"ff044a41",
			4747 => x"0d0a5f04",
			4748 => x"fe844a41",
			4749 => x"07077d04",
			4750 => x"00264a41",
			4751 => x"00004a41",
			4752 => x"07067138",
			4753 => x"0b06fc2c",
			4754 => x"0a01db18",
			4755 => x"0c054810",
			4756 => x"0002a70c",
			4757 => x"0e059d04",
			4758 => x"00004acd",
			4759 => x"07051a04",
			4760 => x"00004acd",
			4761 => x"00434acd",
			4762 => x"00004acd",
			4763 => x"0207ed04",
			4764 => x"ffca4acd",
			4765 => x"00004acd",
			4766 => x"05080410",
			4767 => x"0f09e10c",
			4768 => x"07066c08",
			4769 => x"0002c404",
			4770 => x"00004acd",
			4771 => x"ff704acd",
			4772 => x"00004acd",
			4773 => x"00004acd",
			4774 => x"00004acd",
			4775 => x"07065504",
			4776 => x"00004acd",
			4777 => x"0100f104",
			4778 => x"00884acd",
			4779 => x"00004acd",
			4780 => x"0d08da0c",
			4781 => x"0002dd04",
			4782 => x"00004acd",
			4783 => x"0b074404",
			4784 => x"ff894acd",
			4785 => x"00004acd",
			4786 => x"00004acd",
			4787 => x"0c050b08",
			4788 => x"0600df04",
			4789 => x"00004b49",
			4790 => x"ff114b49",
			4791 => x"0309ef28",
			4792 => x"08025f20",
			4793 => x"0b06ff18",
			4794 => x"0f07e30c",
			4795 => x"0c054508",
			4796 => x"0600e804",
			4797 => x"00004b49",
			4798 => x"00694b49",
			4799 => x"ff924b49",
			4800 => x"09018008",
			4801 => x"07067104",
			4802 => x"00d74b49",
			4803 => x"00004b49",
			4804 => x"00004b49",
			4805 => x"0100ed04",
			4806 => x"ffee4b49",
			4807 => x"00004b49",
			4808 => x"0f09e104",
			4809 => x"ff9b4b49",
			4810 => x"00004b49",
			4811 => x"0601960c",
			4812 => x"0c061a04",
			4813 => x"00004b49",
			4814 => x"01013804",
			4815 => x"00994b49",
			4816 => x"00004b49",
			4817 => x"00004b49",
			4818 => x"0d067908",
			4819 => x"0600df04",
			4820 => x"00004bb5",
			4821 => x"fe8e4bb5",
			4822 => x"0100f82c",
			4823 => x"03098720",
			4824 => x"0b070118",
			4825 => x"06014510",
			4826 => x"03091a08",
			4827 => x"06013504",
			4828 => x"00734bb5",
			4829 => x"ff3b4bb5",
			4830 => x"06014104",
			4831 => x"01194bb5",
			4832 => x"00004bb5",
			4833 => x"03095804",
			4834 => x"ff764bb5",
			4835 => x"00004bb5",
			4836 => x"02090004",
			4837 => x"00174bb5",
			4838 => x"fe8b4bb5",
			4839 => x"07069b08",
			4840 => x"0b070104",
			4841 => x"00004bb5",
			4842 => x"010a4bb5",
			4843 => x"ffed4bb5",
			4844 => x"ff104bb5",
			4845 => x"0c05250c",
			4846 => x"0002a708",
			4847 => x"0e059d04",
			4848 => x"00004c41",
			4849 => x"00624c41",
			4850 => x"00004c41",
			4851 => x"0706140c",
			4852 => x"0c052804",
			4853 => x"00004c41",
			4854 => x"0c05f404",
			4855 => x"ff9e4c41",
			4856 => x"00004c41",
			4857 => x"06014010",
			4858 => x"0c06170c",
			4859 => x"09018308",
			4860 => x"0d07d804",
			4861 => x"00004c41",
			4862 => x"00444c41",
			4863 => x"00004c41",
			4864 => x"00004c41",
			4865 => x"0e096210",
			4866 => x"0c061104",
			4867 => x"00004c41",
			4868 => x"0208fe04",
			4869 => x"00004c41",
			4870 => x"05083e04",
			4871 => x"ffb54c41",
			4872 => x"00004c41",
			4873 => x"0c061a04",
			4874 => x"00004c41",
			4875 => x"08032908",
			4876 => x"08026f04",
			4877 => x"00004c41",
			4878 => x"002b4c41",
			4879 => x"00004c41",
			4880 => x"0a02082c",
			4881 => x"0705450c",
			4882 => x"0600d908",
			4883 => x"07051b04",
			4884 => x"ff574cdd",
			4885 => x"00604cdd",
			4886 => x"fdf34cdd",
			4887 => x"0901871c",
			4888 => x"0c063214",
			4889 => x"01009204",
			4890 => x"07014cdd",
			4891 => x"0a018408",
			4892 => x"01009b04",
			4893 => x"00fb4cdd",
			4894 => x"fe7d4cdd",
			4895 => x"03098704",
			4896 => x"017a4cdd",
			4897 => x"02a94cdd",
			4898 => x"08025a04",
			4899 => x"01364cdd",
			4900 => x"fe824cdd",
			4901 => x"fea24cdd",
			4902 => x"0100d004",
			4903 => x"fe624cdd",
			4904 => x"09015f10",
			4905 => x"020a2d08",
			4906 => x"0e083c04",
			4907 => x"00004cdd",
			4908 => x"01b94cdd",
			4909 => x"0707ad04",
			4910 => x"0ad54cdd",
			4911 => x"00004cdd",
			4912 => x"0b08350c",
			4913 => x"0100f808",
			4914 => x"0802bb04",
			4915 => x"016c4cdd",
			4916 => x"fed44cdd",
			4917 => x"fe684cdd",
			4918 => x"036d4cdd",
			4919 => x"0d067908",
			4920 => x"0a015104",
			4921 => x"00004d51",
			4922 => x"fe8f4d51",
			4923 => x"09019c30",
			4924 => x"03098720",
			4925 => x"0b070118",
			4926 => x"0002e60c",
			4927 => x"03094008",
			4928 => x"07065804",
			4929 => x"00884d51",
			4930 => x"ff504d51",
			4931 => x"012f4d51",
			4932 => x"03096808",
			4933 => x"0d085804",
			4934 => x"ff994d51",
			4935 => x"00004d51",
			4936 => x"00004d51",
			4937 => x"02090004",
			4938 => x"00364d51",
			4939 => x"fe5f4d51",
			4940 => x"07068508",
			4941 => x"09019004",
			4942 => x"01474d51",
			4943 => x"00004d51",
			4944 => x"0c063004",
			4945 => x"00004d51",
			4946 => x"ff964d51",
			4947 => x"ff074d51",
			4948 => x"0a02082c",
			4949 => x"0705450c",
			4950 => x"0600d908",
			4951 => x"0600d504",
			4952 => x"ff6f4ded",
			4953 => x"00514ded",
			4954 => x"fdff4ded",
			4955 => x"0901871c",
			4956 => x"07068514",
			4957 => x"0f096810",
			4958 => x"0002e608",
			4959 => x"0c050b04",
			4960 => x"ff354ded",
			4961 => x"018c4ded",
			4962 => x"07066c04",
			4963 => x"ff464ded",
			4964 => x"011a4ded",
			4965 => x"03444ded",
			4966 => x"02091104",
			4967 => x"00ea4ded",
			4968 => x"fe8e4ded",
			4969 => x"feaa4ded",
			4970 => x"0100d004",
			4971 => x"fe624ded",
			4972 => x"0100df0c",
			4973 => x"0507c704",
			4974 => x"ff6f4ded",
			4975 => x"0c070704",
			4976 => x"040b4ded",
			4977 => x"00004ded",
			4978 => x"0b083510",
			4979 => x"0100f80c",
			4980 => x"0f0a0304",
			4981 => x"fef84ded",
			4982 => x"040b8504",
			4983 => x"01784ded",
			4984 => x"ffd04ded",
			4985 => x"fe694ded",
			4986 => x"02dc4ded",
			4987 => x"07051a04",
			4988 => x"fe744e71",
			4989 => x"0002c418",
			4990 => x"0100dc10",
			4991 => x"0c05f208",
			4992 => x"0e059d04",
			4993 => x"00004e71",
			4994 => x"01344e71",
			4995 => x"02083f04",
			4996 => x"00004e71",
			4997 => x"00464e71",
			4998 => x"0308bf04",
			4999 => x"ff294e71",
			5000 => x"01064e71",
			5001 => x"0507d70c",
			5002 => x"08024104",
			5003 => x"00004e71",
			5004 => x"0b06dc04",
			5005 => x"fe834e71",
			5006 => x"00004e71",
			5007 => x"0100d404",
			5008 => x"feb74e71",
			5009 => x"0100f30c",
			5010 => x"02097008",
			5011 => x"07066f04",
			5012 => x"00b24e71",
			5013 => x"fec64e71",
			5014 => x"01f54e71",
			5015 => x"0c06dc04",
			5016 => x"feb94e71",
			5017 => x"0601b704",
			5018 => x"00ff4e71",
			5019 => x"00004e71",
			5020 => x"0a02084c",
			5021 => x"0e07dc20",
			5022 => x"01009910",
			5023 => x"0e05e008",
			5024 => x"0600cd04",
			5025 => x"01584f35",
			5026 => x"fe8e4f35",
			5027 => x"0c050a04",
			5028 => x"02394f35",
			5029 => x"067d4f35",
			5030 => x"0c05450c",
			5031 => x"0b05a604",
			5032 => x"fe3e4f35",
			5033 => x"0406a304",
			5034 => x"ff2c4f35",
			5035 => x"01724f35",
			5036 => x"fe5e4f35",
			5037 => x"0100f124",
			5038 => x"07067114",
			5039 => x"04097210",
			5040 => x"06013d08",
			5041 => x"0a01e904",
			5042 => x"01cb4f35",
			5043 => x"012e4f35",
			5044 => x"03092204",
			5045 => x"fc3a4f35",
			5046 => x"00f14f35",
			5047 => x"036e4f35",
			5048 => x"0b071008",
			5049 => x"0002e604",
			5050 => x"01824f35",
			5051 => x"fe074f35",
			5052 => x"0e092404",
			5053 => x"fc354f35",
			5054 => x"fe7e4f35",
			5055 => x"0d089a04",
			5056 => x"fe7e4f35",
			5057 => x"014d4f35",
			5058 => x"0a023e0c",
			5059 => x"0209ce04",
			5060 => x"fe6e4f35",
			5061 => x"01011504",
			5062 => x"04fe4f35",
			5063 => x"fff84f35",
			5064 => x"0509e304",
			5065 => x"fe674f35",
			5066 => x"02100704",
			5067 => x"02164f35",
			5068 => x"fe814f35",
			5069 => x"0a023e3c",
			5070 => x"0100f134",
			5071 => x"03098728",
			5072 => x"0002e61c",
			5073 => x"0507f410",
			5074 => x"07065808",
			5075 => x"03077c04",
			5076 => x"00094fc1",
			5077 => x"00de4fc1",
			5078 => x"06013504",
			5079 => x"00004fc1",
			5080 => x"fef84fc1",
			5081 => x"08025a08",
			5082 => x"03092e04",
			5083 => x"00004fc1",
			5084 => x"01494fc1",
			5085 => x"00004fc1",
			5086 => x"0507f408",
			5087 => x"0d079604",
			5088 => x"ffb44fc1",
			5089 => x"00544fc1",
			5090 => x"ff084fc1",
			5091 => x"02093004",
			5092 => x"00004fc1",
			5093 => x"07068504",
			5094 => x"01754fc1",
			5095 => x"00004fc1",
			5096 => x"09018704",
			5097 => x"00004fc1",
			5098 => x"ff014fc1",
			5099 => x"0d0a5f04",
			5100 => x"fe814fc1",
			5101 => x"07077d04",
			5102 => x"003b4fc1",
			5103 => x"00004fc1",
			5104 => x"07051804",
			5105 => x"feaf5045",
			5106 => x"0a01d710",
			5107 => x"0100dc0c",
			5108 => x"0e059d04",
			5109 => x"00005045",
			5110 => x"0408ea04",
			5111 => x"009f5045",
			5112 => x"00005045",
			5113 => x"00005045",
			5114 => x"05081218",
			5115 => x"07065810",
			5116 => x"07061504",
			5117 => x"ff085045",
			5118 => x"0802b308",
			5119 => x"08023c04",
			5120 => x"00005045",
			5121 => x"004a5045",
			5122 => x"00005045",
			5123 => x"07068304",
			5124 => x"ff155045",
			5125 => x"00005045",
			5126 => x"0100f310",
			5127 => x"0b06fe04",
			5128 => x"00005045",
			5129 => x"07068508",
			5130 => x"03097804",
			5131 => x"00005045",
			5132 => x"00f15045",
			5133 => x"00005045",
			5134 => x"030c9904",
			5135 => x"ff815045",
			5136 => x"000d5045",
			5137 => x"0003353c",
			5138 => x"0c065038",
			5139 => x"0a01d718",
			5140 => x"0207ed14",
			5141 => x"0100a10c",
			5142 => x"0f060a04",
			5143 => x"ff5350e1",
			5144 => x"01008004",
			5145 => x"000050e1",
			5146 => x"016450e1",
			5147 => x"0c052804",
			5148 => x"000050e1",
			5149 => x"fead50e1",
			5150 => x"017650e1",
			5151 => x"03091a10",
			5152 => x"06013508",
			5153 => x"0100d004",
			5154 => x"ff9150e1",
			5155 => x"007950e1",
			5156 => x"0c05f804",
			5157 => x"000050e1",
			5158 => x"fd7a50e1",
			5159 => x"0a01e904",
			5160 => x"015d50e1",
			5161 => x"06013a04",
			5162 => x"fec050e1",
			5163 => x"07066c04",
			5164 => x"ffa350e1",
			5165 => x"00c450e1",
			5166 => x"072750e1",
			5167 => x"0b06cc04",
			5168 => x"fe6450e1",
			5169 => x"0b06dc08",
			5170 => x"0901ce04",
			5171 => x"012350e1",
			5172 => x"000050e1",
			5173 => x"0509e304",
			5174 => x"fea150e1",
			5175 => x"000050e1",
			5176 => x"08025f34",
			5177 => x"0e067114",
			5178 => x"0600d908",
			5179 => x"0a014504",
			5180 => x"fea451b5",
			5181 => x"08f551b5",
			5182 => x"0e060f04",
			5183 => x"fe6651b5",
			5184 => x"0100a104",
			5185 => x"05d051b5",
			5186 => x"fe7751b5",
			5187 => x"0100ef18",
			5188 => x"07057304",
			5189 => x"099d51b5",
			5190 => x"0e073b04",
			5191 => x"fe7e51b5",
			5192 => x"0d086d08",
			5193 => x"07068504",
			5194 => x"03fc51b5",
			5195 => x"027351b5",
			5196 => x"0c061504",
			5197 => x"043251b5",
			5198 => x"013351b5",
			5199 => x"06013d04",
			5200 => x"014d51b5",
			5201 => x"fe6d51b5",
			5202 => x"00031a18",
			5203 => x"0100f314",
			5204 => x"0309b010",
			5205 => x"0c060f04",
			5206 => x"045051b5",
			5207 => x"0a01f704",
			5208 => x"fe7751b5",
			5209 => x"07066f04",
			5210 => x"037151b5",
			5211 => x"feae51b5",
			5212 => x"093e51b5",
			5213 => x"fe6251b5",
			5214 => x"0a02230c",
			5215 => x"040a2804",
			5216 => x"fe6451b5",
			5217 => x"01005e04",
			5218 => x"fe9151b5",
			5219 => x"052e51b5",
			5220 => x"0d0a5f04",
			5221 => x"fe5951b5",
			5222 => x"0d0a790c",
			5223 => x"0509f008",
			5224 => x"0509e304",
			5225 => x"ff7d51b5",
			5226 => x"017751b5",
			5227 => x"fec051b5",
			5228 => x"fe5e51b5",
			5229 => x"0802794c",
			5230 => x"06014128",
			5231 => x"0e07dc14",
			5232 => x"06010a10",
			5233 => x"0c05480c",
			5234 => x"0e059d04",
			5235 => x"ffc85279",
			5236 => x"0900f704",
			5237 => x"01835279",
			5238 => x"007c5279",
			5239 => x"ffa25279",
			5240 => x"fe585279",
			5241 => x"09018310",
			5242 => x"0706850c",
			5243 => x"07066c08",
			5244 => x"07065804",
			5245 => x"01725279",
			5246 => x"00005279",
			5247 => x"01d05279",
			5248 => x"00005279",
			5249 => x"ff8f5279",
			5250 => x"0309a31c",
			5251 => x"04094514",
			5252 => x"0b06ec0c",
			5253 => x"0e08f008",
			5254 => x"08025304",
			5255 => x"00005279",
			5256 => x"ff135279",
			5257 => x"00005279",
			5258 => x"09018004",
			5259 => x"012e5279",
			5260 => x"fff55279",
			5261 => x"0c05f404",
			5262 => x"00005279",
			5263 => x"feb35279",
			5264 => x"0b071e04",
			5265 => x"016d5279",
			5266 => x"fff25279",
			5267 => x"0b071e04",
			5268 => x"fe685279",
			5269 => x"0c063408",
			5270 => x"0100fc04",
			5271 => x"01ea5279",
			5272 => x"ffec5279",
			5273 => x"0d0a5f04",
			5274 => x"fea25279",
			5275 => x"0d0a6c04",
			5276 => x"00005279",
			5277 => x"fff65279",
			5278 => x"0004084c",
			5279 => x"03097830",
			5280 => x"0002dd1c",
			5281 => x"0207cf14",
			5282 => x"0900f30c",
			5283 => x"0e059d04",
			5284 => x"00005315",
			5285 => x"07051a04",
			5286 => x"00005315",
			5287 => x"00815315",
			5288 => x"09011304",
			5289 => x"ff545315",
			5290 => x"00005315",
			5291 => x"06013b04",
			5292 => x"00b45315",
			5293 => x"00005315",
			5294 => x"08025304",
			5295 => x"00005315",
			5296 => x"0a01e904",
			5297 => x"00005315",
			5298 => x"0f096808",
			5299 => x"0c063004",
			5300 => x"ff245315",
			5301 => x"00005315",
			5302 => x"00005315",
			5303 => x"0706850c",
			5304 => x"09019008",
			5305 => x"06014104",
			5306 => x"00005315",
			5307 => x"00fa5315",
			5308 => x"00005315",
			5309 => x"05088604",
			5310 => x"ffa35315",
			5311 => x"0901f408",
			5312 => x"06019904",
			5313 => x"00655315",
			5314 => x"00005315",
			5315 => x"00005315",
			5316 => x"fef75315",
			5317 => x"0a021d4c",
			5318 => x"0100f140",
			5319 => x"0e07dc20",
			5320 => x"00028d1c",
			5321 => x"0c052810",
			5322 => x"0f061208",
			5323 => x"0600cd04",
			5324 => x"026153d9",
			5325 => x"fe9253d9",
			5326 => x"0900fe04",
			5327 => x"04a853d9",
			5328 => x"017353d9",
			5329 => x"07055f08",
			5330 => x"09010f04",
			5331 => x"ff1753d9",
			5332 => x"011853d9",
			5333 => x"fe6753d9",
			5334 => x"fdf053d9",
			5335 => x"0309a318",
			5336 => x"0002e60c",
			5337 => x"09018308",
			5338 => x"0e090704",
			5339 => x"01d053d9",
			5340 => x"02dc53d9",
			5341 => x"fef153d9",
			5342 => x"0c061004",
			5343 => x"029e53d9",
			5344 => x"03098704",
			5345 => x"fe8853d9",
			5346 => x"009b53d9",
			5347 => x"07067204",
			5348 => x"040d53d9",
			5349 => x"023853d9",
			5350 => x"09018708",
			5351 => x"05082e04",
			5352 => x"fee653d9",
			5353 => x"01fc53d9",
			5354 => x"fe6f53d9",
			5355 => x"0a02300c",
			5356 => x"040a6904",
			5357 => x"fe7753d9",
			5358 => x"0003aa04",
			5359 => x"052853d9",
			5360 => x"ff6f53d9",
			5361 => x"0509e304",
			5362 => x"fe6253d9",
			5363 => x"0509f004",
			5364 => x"006253d9",
			5365 => x"fe7953d9",
			5366 => x"0a020850",
			5367 => x"0e07dc2c",
			5368 => x"0600eb18",
			5369 => x"0c054314",
			5370 => x"0e059d04",
			5371 => x"febe54a5",
			5372 => x"01009008",
			5373 => x"0c04f104",
			5374 => x"030a54a5",
			5375 => x"000054a5",
			5376 => x"0900fe04",
			5377 => x"ff0054a5",
			5378 => x"000054a5",
			5379 => x"099354a5",
			5380 => x"0b059904",
			5381 => x"fe4c54a5",
			5382 => x"0c05450c",
			5383 => x"0406a304",
			5384 => x"ff0a54a5",
			5385 => x"0100a604",
			5386 => x"01b054a5",
			5387 => x"000054a5",
			5388 => x"fe6954a5",
			5389 => x"09018720",
			5390 => x"07068514",
			5391 => x"03098710",
			5392 => x"06013b08",
			5393 => x"0d086504",
			5394 => x"01be54a5",
			5395 => x"006e54a5",
			5396 => x"03092204",
			5397 => x"fcb054a5",
			5398 => x"00a754a5",
			5399 => x"034954a5",
			5400 => x"07068808",
			5401 => x"0e091504",
			5402 => x"012254a5",
			5403 => x"fe8454a5",
			5404 => x"fd9454a5",
			5405 => x"fe8a54a5",
			5406 => x"0a023e0c",
			5407 => x"0209ce04",
			5408 => x"fe7054a5",
			5409 => x"0309ef04",
			5410 => x"055954a5",
			5411 => x"017654a5",
			5412 => x"0509e304",
			5413 => x"fe6854a5",
			5414 => x"02100704",
			5415 => x"01ca54a5",
			5416 => x"fe8754a5",
			5417 => x"07051804",
			5418 => x"fee35531",
			5419 => x"0a01d70c",
			5420 => x"0e059d04",
			5421 => x"00005531",
			5422 => x"0c05f204",
			5423 => x"00b15531",
			5424 => x"00005531",
			5425 => x"05081218",
			5426 => x"0d087f14",
			5427 => x"0d086510",
			5428 => x"03091a08",
			5429 => x"08024104",
			5430 => x"00005531",
			5431 => x"ff175531",
			5432 => x"0100eb04",
			5433 => x"00d35531",
			5434 => x"ffee5531",
			5435 => x"fef75531",
			5436 => x"00005531",
			5437 => x"0b070e0c",
			5438 => x"0d086504",
			5439 => x"001e5531",
			5440 => x"0d088204",
			5441 => x"ff8d5531",
			5442 => x"00005531",
			5443 => x"07069b0c",
			5444 => x"0100f108",
			5445 => x"0d086d04",
			5446 => x"00005531",
			5447 => x"00f35531",
			5448 => x"00005531",
			5449 => x"0d0a6c04",
			5450 => x"ffd55531",
			5451 => x"00005531",
			5452 => x"0d067908",
			5453 => x"0a015104",
			5454 => x"000055b5",
			5455 => x"fe9555b5",
			5456 => x"0100f838",
			5457 => x"03098728",
			5458 => x"0b070120",
			5459 => x"03091a10",
			5460 => x"0a01db08",
			5461 => x"0f067a04",
			5462 => x"000055b5",
			5463 => x"009455b5",
			5464 => x"08024104",
			5465 => x"000055b5",
			5466 => x"fefa55b5",
			5467 => x"0100eb08",
			5468 => x"07068504",
			5469 => x"012d55b5",
			5470 => x"000055b5",
			5471 => x"0002e604",
			5472 => x"002a55b5",
			5473 => x"ff9155b5",
			5474 => x"02090004",
			5475 => x"002855b5",
			5476 => x"fe7655b5",
			5477 => x"07069b0c",
			5478 => x"0b070104",
			5479 => x"000055b5",
			5480 => x"07068504",
			5481 => x"013755b5",
			5482 => x"000055b5",
			5483 => x"ffdf55b5",
			5484 => x"ff0455b5",
			5485 => x"00030c54",
			5486 => x"0c061434",
			5487 => x"0e07dc14",
			5488 => x"06010a10",
			5489 => x"0c05480c",
			5490 => x"0e059d04",
			5491 => x"ffc35689",
			5492 => x"0900f304",
			5493 => x"01d55689",
			5494 => x"007f5689",
			5495 => x"ff1e5689",
			5496 => x"fe385689",
			5497 => x"0a01ec08",
			5498 => x"0100ef04",
			5499 => x"017a5689",
			5500 => x"ffec5689",
			5501 => x"0309780c",
			5502 => x"0b06bc04",
			5503 => x"00005689",
			5504 => x"00030204",
			5505 => x"fe955689",
			5506 => x"00005689",
			5507 => x"0002f604",
			5508 => x"01c85689",
			5509 => x"05081304",
			5510 => x"ffeb5689",
			5511 => x"00005689",
			5512 => x"0308e704",
			5513 => x"fdc25689",
			5514 => x"04094508",
			5515 => x"0a01ec04",
			5516 => x"01995689",
			5517 => x"00005689",
			5518 => x"0c061608",
			5519 => x"0002ee04",
			5520 => x"013c5689",
			5521 => x"00005689",
			5522 => x"08026f04",
			5523 => x"fe285689",
			5524 => x"0b071004",
			5525 => x"01355689",
			5526 => x"00005689",
			5527 => x"0d082504",
			5528 => x"fe6a5689",
			5529 => x"06016a08",
			5530 => x"09019004",
			5531 => x"02135689",
			5532 => x"ff0e5689",
			5533 => x"0d0a5f04",
			5534 => x"fe865689",
			5535 => x"0c06e504",
			5536 => x"012c5689",
			5537 => x"ff9d5689",
			5538 => x"00030c60",
			5539 => x"08025320",
			5540 => x"0e059d04",
			5541 => x"ff025775",
			5542 => x"0100920c",
			5543 => x"0b057608",
			5544 => x"0c04ee04",
			5545 => x"02b75775",
			5546 => x"00005775",
			5547 => x"066f5775",
			5548 => x"0b059904",
			5549 => x"feb65775",
			5550 => x"0100ef08",
			5551 => x"06013d04",
			5552 => x"01a05775",
			5553 => x"00995775",
			5554 => x"ff3a5775",
			5555 => x"07066c20",
			5556 => x"07065a10",
			5557 => x"0d084a08",
			5558 => x"0208f004",
			5559 => x"fe635775",
			5560 => x"fffc5775",
			5561 => x"0100f104",
			5562 => x"01875775",
			5563 => x"00005775",
			5564 => x"02091108",
			5565 => x"0507f404",
			5566 => x"000d5775",
			5567 => x"fe975775",
			5568 => x"05082e04",
			5569 => x"fc1c5775",
			5570 => x"00005775",
			5571 => x"07066f10",
			5572 => x"0e092408",
			5573 => x"09018004",
			5574 => x"01a15775",
			5575 => x"ff375775",
			5576 => x"0d087404",
			5577 => x"075c5775",
			5578 => x"02695775",
			5579 => x"06014104",
			5580 => x"017c5775",
			5581 => x"0409b308",
			5582 => x"05081204",
			5583 => x"fffa5775",
			5584 => x"fe1a5775",
			5585 => x"00cc5775",
			5586 => x"0100d004",
			5587 => x"fe625775",
			5588 => x"09015f08",
			5589 => x"06016b04",
			5590 => x"03b25775",
			5591 => x"ff1a5775",
			5592 => x"0509a908",
			5593 => x"06015204",
			5594 => x"00fd5775",
			5595 => x"fe6b5775",
			5596 => x"02975775",
			5597 => x"0003354c",
			5598 => x"0c065048",
			5599 => x"0802411c",
			5600 => x"0e07dc14",
			5601 => x"0100a10c",
			5602 => x"0e060f08",
			5603 => x"0c054304",
			5604 => x"ff5f5831",
			5605 => x"004a5831",
			5606 => x"01895831",
			5607 => x"0c052804",
			5608 => x"00005831",
			5609 => x"feb95831",
			5610 => x"09017604",
			5611 => x"01725831",
			5612 => x"00005831",
			5613 => x"03091a14",
			5614 => x"0c05f80c",
			5615 => x"0d080e08",
			5616 => x"07064004",
			5617 => x"ff5b5831",
			5618 => x"00005831",
			5619 => x"00005831",
			5620 => x"0b06cf04",
			5621 => x"00005831",
			5622 => x"fdbc5831",
			5623 => x"08025308",
			5624 => x"0b06ce04",
			5625 => x"00005831",
			5626 => x"01755831",
			5627 => x"03097808",
			5628 => x"0b070104",
			5629 => x"00005831",
			5630 => x"fe9f5831",
			5631 => x"0002ee04",
			5632 => x"01845831",
			5633 => x"00005831",
			5634 => x"03f35831",
			5635 => x"0b06cc04",
			5636 => x"fe665831",
			5637 => x"0b06dc08",
			5638 => x"0e095104",
			5639 => x"011b5831",
			5640 => x"00005831",
			5641 => x"0509e304",
			5642 => x"feaa5831",
			5643 => x"00005831",
			5644 => x"00032458",
			5645 => x"0e07dc20",
			5646 => x"0207801c",
			5647 => x"07058c18",
			5648 => x"0e065a10",
			5649 => x"0c054308",
			5650 => x"0c04d004",
			5651 => x"00005925",
			5652 => x"fead5925",
			5653 => x"05064404",
			5654 => x"020a5925",
			5655 => x"00005925",
			5656 => x"0c054c04",
			5657 => x"019f5925",
			5658 => x"00005925",
			5659 => x"fed15925",
			5660 => x"fe755925",
			5661 => x"0c061618",
			5662 => x"09018714",
			5663 => x"07068510",
			5664 => x"07066c08",
			5665 => x"09017a04",
			5666 => x"01975925",
			5667 => x"00025925",
			5668 => x"0208dd04",
			5669 => x"00005925",
			5670 => x"025a5925",
			5671 => x"ffe95925",
			5672 => x"feeb5925",
			5673 => x"0d087f14",
			5674 => x"0002dd08",
			5675 => x"03092e04",
			5676 => x"00005925",
			5677 => x"01525925",
			5678 => x"02096008",
			5679 => x"0b06df04",
			5680 => x"00005925",
			5681 => x"fd295925",
			5682 => x"00005925",
			5683 => x"0b071004",
			5684 => x"01e05925",
			5685 => x"0e098704",
			5686 => x"ff6f5925",
			5687 => x"00c65925",
			5688 => x"020b7714",
			5689 => x"0802cc10",
			5690 => x"0d082504",
			5691 => x"fead5925",
			5692 => x"0b06dc08",
			5693 => x"0e095104",
			5694 => x"01875925",
			5695 => x"00005925",
			5696 => x"fefe5925",
			5697 => x"fe685925",
			5698 => x"0a02900c",
			5699 => x"0508c104",
			5700 => x"05715925",
			5701 => x"030bbc04",
			5702 => x"00005925",
			5703 => x"01db5925",
			5704 => x"fe935925",
			5705 => x"08027960",
			5706 => x"08025320",
			5707 => x"0e059d04",
			5708 => x"ff155a19",
			5709 => x"01009204",
			5710 => x"02f45a19",
			5711 => x"0f07010c",
			5712 => x"01009b08",
			5713 => x"07054b04",
			5714 => x"ffaa5a19",
			5715 => x"01905a19",
			5716 => x"fea75a19",
			5717 => x"09017d04",
			5718 => x"019f5a19",
			5719 => x"06013b04",
			5720 => x"01425a19",
			5721 => x"ff835a19",
			5722 => x"07066c20",
			5723 => x"07065a10",
			5724 => x"0d084a08",
			5725 => x"0208f004",
			5726 => x"fe5f5a19",
			5727 => x"00005a19",
			5728 => x"09018304",
			5729 => x"01895a19",
			5730 => x"00005a19",
			5731 => x"02091108",
			5732 => x"0507f404",
			5733 => x"00145a19",
			5734 => x"feb45a19",
			5735 => x"0f094d04",
			5736 => x"fc8e5a19",
			5737 => x"00005a19",
			5738 => x"07066f10",
			5739 => x"03097808",
			5740 => x"09018004",
			5741 => x"01305a19",
			5742 => x"ff345a19",
			5743 => x"0100f104",
			5744 => x"02dd5a19",
			5745 => x"00005a19",
			5746 => x"06014104",
			5747 => x"01555a19",
			5748 => x"0d089a08",
			5749 => x"05081204",
			5750 => x"00005a19",
			5751 => x"fe2f5a19",
			5752 => x"00b85a19",
			5753 => x"0100d004",
			5754 => x"fe625a19",
			5755 => x"09015f08",
			5756 => x"08032904",
			5757 => x"02df5a19",
			5758 => x"ff825a19",
			5759 => x"0509a90c",
			5760 => x"08029108",
			5761 => x"09019c04",
			5762 => x"009c5a19",
			5763 => x"ff2a5a19",
			5764 => x"fe6c5a19",
			5765 => x"022f5a19",
			5766 => x"07051a04",
			5767 => x"fe7d5add",
			5768 => x"07066c3c",
			5769 => x"08024118",
			5770 => x"0207cf10",
			5771 => x"0600d904",
			5772 => x"014d5add",
			5773 => x"0c052808",
			5774 => x"0f067a04",
			5775 => x"ff825add",
			5776 => x"00b35add",
			5777 => x"ff215add",
			5778 => x"09017604",
			5779 => x"01425add",
			5780 => x"00005add",
			5781 => x"0d083814",
			5782 => x"0002c404",
			5783 => x"00005add",
			5784 => x"0f093d08",
			5785 => x"07065904",
			5786 => x"feae5add",
			5787 => x"00005add",
			5788 => x"0507e404",
			5789 => x"ffe45add",
			5790 => x"00005add",
			5791 => x"0a01ec04",
			5792 => x"01255add",
			5793 => x"06013e04",
			5794 => x"fedd5add",
			5795 => x"06014904",
			5796 => x"009b5add",
			5797 => x"00005add",
			5798 => x"07068510",
			5799 => x"0901900c",
			5800 => x"0208dd04",
			5801 => x"00005add",
			5802 => x"0d084c04",
			5803 => x"00005add",
			5804 => x"01645add",
			5805 => x"fff65add",
			5806 => x"0e09c104",
			5807 => x"ff355add",
			5808 => x"0901ff0c",
			5809 => x"08031808",
			5810 => x"06019d04",
			5811 => x"00fa5add",
			5812 => x"00005add",
			5813 => x"00005add",
			5814 => x"ffae5add",
			5815 => x"07051a04",
			5816 => x"fe785b93",
			5817 => x"0a029054",
			5818 => x"0d087f3c",
			5819 => x"0a01ec20",
			5820 => x"0c05f810",
			5821 => x"0207cf08",
			5822 => x"07058c04",
			5823 => x"009c5b93",
			5824 => x"ff015b93",
			5825 => x"0100f104",
			5826 => x"016d5b93",
			5827 => x"00005b93",
			5828 => x"0507e608",
			5829 => x"06013504",
			5830 => x"004f5b93",
			5831 => x"fe9c5b93",
			5832 => x"02090004",
			5833 => x"01225b93",
			5834 => x"ffca5b93",
			5835 => x"0309780c",
			5836 => x"0f096808",
			5837 => x"06013904",
			5838 => x"00005b93",
			5839 => x"fede5b93",
			5840 => x"00005b93",
			5841 => x"02093a08",
			5842 => x"07066e04",
			5843 => x"00d85b93",
			5844 => x"00005b93",
			5845 => x"0209ce04",
			5846 => x"fed45b93",
			5847 => x"00005b93",
			5848 => x"07068508",
			5849 => x"0100f304",
			5850 => x"01bc5b93",
			5851 => x"00005b93",
			5852 => x"030a4904",
			5853 => x"ff225b93",
			5854 => x"01013908",
			5855 => x"0d08da04",
			5856 => x"00005b93",
			5857 => x"010e5b93",
			5858 => x"fffc5b93",
			5859 => x"fee35b93",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1940, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(3878, initial_addr_3'length));
	end generate gen_rom_4;

	gen_rom_5: if SELECT_ROM = 5 generate
		bank <= (
			0 => x"00000005",
			1 => x"00000009",
			2 => x"0000000d",
			3 => x"00000011",
			4 => x"00000015",
			5 => x"00000019",
			6 => x"0000001d",
			7 => x"00000021",
			8 => x"00000025",
			9 => x"00000029",
			10 => x"0000002d",
			11 => x"00000031",
			12 => x"00000035",
			13 => x"00000039",
			14 => x"0000003d",
			15 => x"00000041",
			16 => x"00000045",
			17 => x"00000049",
			18 => x"0000004d",
			19 => x"00000051",
			20 => x"00000055",
			21 => x"00000059",
			22 => x"0000005d",
			23 => x"00000061",
			24 => x"00000065",
			25 => x"00000069",
			26 => x"0000006d",
			27 => x"00000071",
			28 => x"00000075",
			29 => x"00000079",
			30 => x"0000007d",
			31 => x"00000081",
			32 => x"00000085",
			33 => x"040d4204",
			34 => x"ff550091",
			35 => x"00000091",
			36 => x"040d4204",
			37 => x"ff8e009d",
			38 => x"0000009d",
			39 => x"040d4204",
			40 => x"ffd500a9",
			41 => x"000000a9",
			42 => x"07069b04",
			43 => x"fff400b5",
			44 => x"000000b5",
			45 => x"020ac304",
			46 => x"ffcb00c1",
			47 => x"000000c1",
			48 => x"040f7004",
			49 => x"ffc100cd",
			50 => x"000000cd",
			51 => x"0c05f504",
			52 => x"000000d9",
			53 => x"000500d9",
			54 => x"040f7004",
			55 => x"ffea00e5",
			56 => x"000000e5",
			57 => x"040e2304",
			58 => x"fff000f1",
			59 => x"000000f1",
			60 => x"040f7004",
			61 => x"ffe600fd",
			62 => x"000000fd",
			63 => x"0c05f504",
			64 => x"00000109",
			65 => x"00040109",
			66 => x"0c063204",
			67 => x"ff8e011d",
			68 => x"0100de04",
			69 => x"0051011d",
			70 => x"0000011d",
			71 => x"07068604",
			72 => x"ffaf0131",
			73 => x"0100da04",
			74 => x"00300131",
			75 => x"00000131",
			76 => x"0c05f504",
			77 => x"00000145",
			78 => x"0f085c04",
			79 => x"00000145",
			80 => x"000c0145",
			81 => x"07069b08",
			82 => x"04129904",
			83 => x"ff240161",
			84 => x"00000161",
			85 => x"09018304",
			86 => x"00770161",
			87 => x"00000161",
			88 => x"07068608",
			89 => x"0410e104",
			90 => x"ff69017d",
			91 => x"0000017d",
			92 => x"0100ed04",
			93 => x"0074017d",
			94 => x"0000017d",
			95 => x"020bf304",
			96 => x"fe590199",
			97 => x"09019008",
			98 => x"0601a204",
			99 => x"03810199",
			100 => x"02a30199",
			101 => x"fe6f0199",
			102 => x"0c05f504",
			103 => x"fee601b5",
			104 => x"0100d008",
			105 => x"0f085c04",
			106 => x"000001b5",
			107 => x"009b01b5",
			108 => x"000001b5",
			109 => x"0c063204",
			110 => x"ff8601d1",
			111 => x"0100de08",
			112 => x"08051904",
			113 => x"005a01d1",
			114 => x"000001d1",
			115 => x"000001d1",
			116 => x"0c05f504",
			117 => x"ffd401ed",
			118 => x"02096604",
			119 => x"000001ed",
			120 => x"0306a504",
			121 => x"000001ed",
			122 => x"000c01ed",
			123 => x"0c05f504",
			124 => x"fff50209",
			125 => x"02096604",
			126 => x"00000209",
			127 => x"0f085c04",
			128 => x"00000209",
			129 => x"001f0209",
			130 => x"0c05f504",
			131 => x"00000225",
			132 => x"0f085c04",
			133 => x"00000225",
			134 => x"02096604",
			135 => x"00000225",
			136 => x"00130225",
			137 => x"0c05f504",
			138 => x"00000241",
			139 => x"02096604",
			140 => x"00000241",
			141 => x"0306a504",
			142 => x"00000241",
			143 => x"00190241",
			144 => x"020bf30c",
			145 => x"04118b04",
			146 => x"fe6b0265",
			147 => x"0306a504",
			148 => x"fe6d0265",
			149 => x"02b90265",
			150 => x"0100f504",
			151 => x"01a50265",
			152 => x"fed00265",
			153 => x"020bf30c",
			154 => x"07068604",
			155 => x"fe660289",
			156 => x"0b06fc04",
			157 => x"02360289",
			158 => x"fe780289",
			159 => x"0100f504",
			160 => x"019d0289",
			161 => x"ff200289",
			162 => x"0706860c",
			163 => x"020ac304",
			164 => x"fe7102ad",
			165 => x"0004c104",
			166 => x"fffe02ad",
			167 => x"000002ad",
			168 => x"0100d404",
			169 => x"018302ad",
			170 => x"ff1202ad",
			171 => x"0c063208",
			172 => x"0412b204",
			173 => x"fe8202d1",
			174 => x"000002d1",
			175 => x"0100de08",
			176 => x"0006ce04",
			177 => x"014602d1",
			178 => x"000002d1",
			179 => x"ff8d02d1",
			180 => x"0c063208",
			181 => x"0412b204",
			182 => x"feb702f5",
			183 => x"000002f5",
			184 => x"0100ed08",
			185 => x"07067204",
			186 => x"000002f5",
			187 => x"00e302f5",
			188 => x"000002f5",
			189 => x"0c05f504",
			190 => x"fe890319",
			191 => x"0100d008",
			192 => x"07068604",
			193 => x"00000319",
			194 => x"012c0319",
			195 => x"0c06dc04",
			196 => x"ff540319",
			197 => x"00000319",
			198 => x"0c05f504",
			199 => x"fea8033d",
			200 => x"0100d008",
			201 => x"0f085c04",
			202 => x"0000033d",
			203 => x"00e3033d",
			204 => x"00057a04",
			205 => x"ffa7033d",
			206 => x"0000033d",
			207 => x"020cab10",
			208 => x"020c2a08",
			209 => x"020bf304",
			210 => x"d46e0369",
			211 => x"d6430369",
			212 => x"01011f04",
			213 => x"eadb0369",
			214 => x"d4850369",
			215 => x"01013a04",
			216 => x"ec040369",
			217 => x"d4b00369",
			218 => x"040d4204",
			219 => x"feb9038d",
			220 => x"0c05f504",
			221 => x"0000038d",
			222 => x"0100ef08",
			223 => x"01007304",
			224 => x"0000038d",
			225 => x"0090038d",
			226 => x"0000038d",
			227 => x"0c05f504",
			228 => x"feee03b1",
			229 => x"0100d00c",
			230 => x"06015304",
			231 => x"000003b1",
			232 => x"00072404",
			233 => x"009503b1",
			234 => x"000003b1",
			235 => x"000003b1",
			236 => x"040d4204",
			237 => x"ff1a03d5",
			238 => x"0c05f504",
			239 => x"000003d5",
			240 => x"0100ef08",
			241 => x"01007304",
			242 => x"000003d5",
			243 => x"005503d5",
			244 => x"000003d5",
			245 => x"0c05f504",
			246 => x"ff4403f9",
			247 => x"0100ed0c",
			248 => x"02096604",
			249 => x"000003f9",
			250 => x"00072404",
			251 => x"00b903f9",
			252 => x"000003f9",
			253 => x"000003f9",
			254 => x"0c05f504",
			255 => x"0000041d",
			256 => x"0100ed0c",
			257 => x"0f085c04",
			258 => x"0000041d",
			259 => x"02096604",
			260 => x"0000041d",
			261 => x"007e041d",
			262 => x"0000041d",
			263 => x"020bf310",
			264 => x"0c05f504",
			265 => x"fe5f0449",
			266 => x"04118b04",
			267 => x"fe690449",
			268 => x"04182404",
			269 => x"06c70449",
			270 => x"ff040449",
			271 => x"0100f504",
			272 => x"01e90449",
			273 => x"fe8c0449",
			274 => x"020bf310",
			275 => x"0c05f504",
			276 => x"fe670475",
			277 => x"0100cf08",
			278 => x"0f072b04",
			279 => x"00000475",
			280 => x"022a0475",
			281 => x"fe720475",
			282 => x"01011704",
			283 => x"019b0475",
			284 => x"ff300475",
			285 => x"020bf310",
			286 => x"04129904",
			287 => x"fe6804a1",
			288 => x"0005b008",
			289 => x"0c050c04",
			290 => x"000004a1",
			291 => x"016204a1",
			292 => x"fe9204a1",
			293 => x"01011704",
			294 => x"019404a1",
			295 => x"ff5b04a1",
			296 => x"020bf310",
			297 => x"0a02100c",
			298 => x"07069b04",
			299 => x"fec504cd",
			300 => x"0409a004",
			301 => x"000004cd",
			302 => x"014b04cd",
			303 => x"fe6a04cd",
			304 => x"0100f504",
			305 => x"018a04cd",
			306 => x"ffa604cd",
			307 => x"040df508",
			308 => x"0c06aa04",
			309 => x"fe7004f9",
			310 => x"000004f9",
			311 => x"0c05f504",
			312 => x"feee04f9",
			313 => x"0100d008",
			314 => x"01007304",
			315 => x"000004f9",
			316 => x"017e04f9",
			317 => x"000004f9",
			318 => x"0c063210",
			319 => x"020a4604",
			320 => x"fe6b052d",
			321 => x"00058704",
			322 => x"fef6052d",
			323 => x"0a032c04",
			324 => x"0107052d",
			325 => x"0000052d",
			326 => x"0100ed08",
			327 => x"00033504",
			328 => x"0000052d",
			329 => x"0191052d",
			330 => x"feb1052d",
			331 => x"020c2a14",
			332 => x"020bf304",
			333 => x"fe4f0561",
			334 => x"0c068904",
			335 => x"05ed0561",
			336 => x"0c06aa04",
			337 => x"feaa0561",
			338 => x"0c06c304",
			339 => x"017d0561",
			340 => x"ff090561",
			341 => x"01011f04",
			342 => x"063a0561",
			343 => x"fe690561",
			344 => x"0c05f504",
			345 => x"0000058d",
			346 => x"06021810",
			347 => x"06015304",
			348 => x"0000058d",
			349 => x"0306a504",
			350 => x"0000058d",
			351 => x"02096604",
			352 => x"0000058d",
			353 => x"003b058d",
			354 => x"0000058d",
			355 => x"0c05f504",
			356 => x"fe7805c1",
			357 => x"0100d410",
			358 => x"06015304",
			359 => x"000005c1",
			360 => x"01007304",
			361 => x"000005c1",
			362 => x"0100d004",
			363 => x"014905c1",
			364 => x"000005c1",
			365 => x"0c06dc04",
			366 => x"ff0105c1",
			367 => x"000005c1",
			368 => x"020bf318",
			369 => x"0c05f504",
			370 => x"fe6805fd",
			371 => x"0e08f010",
			372 => x"06015304",
			373 => x"fef805fd",
			374 => x"06017008",
			375 => x"02096604",
			376 => x"000005fd",
			377 => x"01d405fd",
			378 => x"000005fd",
			379 => x"fe7905fd",
			380 => x"0901ca04",
			381 => x"019805fd",
			382 => x"ff5005fd",
			383 => x"020bf31c",
			384 => x"0c05f504",
			385 => x"fe5d064b",
			386 => x"0c05f604",
			387 => x"ff5a064b",
			388 => x"0c063a10",
			389 => x"0c063204",
			390 => x"fe72064b",
			391 => x"0c063304",
			392 => x"00fb064b",
			393 => x"0c063404",
			394 => x"feaf064b",
			395 => x"0000064b",
			396 => x"fe5f064b",
			397 => x"0100f508",
			398 => x"0f0c0904",
			399 => x"02eb064b",
			400 => x"0215064b",
			401 => x"fe7d064b",
			402 => x"0000064d",
			403 => x"00000651",
			404 => x"00000655",
			405 => x"00000659",
			406 => x"0000065d",
			407 => x"00000661",
			408 => x"00000665",
			409 => x"00000669",
			410 => x"0000066d",
			411 => x"00000671",
			412 => x"00000675",
			413 => x"00000679",
			414 => x"0000067d",
			415 => x"00000681",
			416 => x"00000685",
			417 => x"00000689",
			418 => x"0000068d",
			419 => x"00000691",
			420 => x"00000695",
			421 => x"00000699",
			422 => x"0000069d",
			423 => x"000006a1",
			424 => x"000006a5",
			425 => x"000006a9",
			426 => x"000006ad",
			427 => x"000006b1",
			428 => x"000006b5",
			429 => x"000006b9",
			430 => x"000006bd",
			431 => x"000006c1",
			432 => x"000006c5",
			433 => x"000006c9",
			434 => x"000006cd",
			435 => x"040d4204",
			436 => x"ff7b06d9",
			437 => x"000006d9",
			438 => x"040d4204",
			439 => x"ffcc06e5",
			440 => x"000006e5",
			441 => x"07069b04",
			442 => x"ffee06f1",
			443 => x"000006f1",
			444 => x"020ac304",
			445 => x"ffc206fd",
			446 => x"000006fd",
			447 => x"07068604",
			448 => x"00000709",
			449 => x"00010709",
			450 => x"040f7004",
			451 => x"ffc70715",
			452 => x"00000715",
			453 => x"07060204",
			454 => x"00000721",
			455 => x"00010721",
			456 => x"040f7004",
			457 => x"ffed072d",
			458 => x"0000072d",
			459 => x"040e2304",
			460 => x"fff30739",
			461 => x"00000739",
			462 => x"040f7004",
			463 => x"ffeb0745",
			464 => x"00000745",
			465 => x"020bf304",
			466 => x"fe670759",
			467 => x"0100f504",
			468 => x"01ce0759",
			469 => x"fe960759",
			470 => x"0c063204",
			471 => x"ff95076d",
			472 => x"0100de04",
			473 => x"0048076d",
			474 => x"0000076d",
			475 => x"07068604",
			476 => x"ffb60781",
			477 => x"0100da04",
			478 => x"002d0781",
			479 => x"00000781",
			480 => x"0c05f504",
			481 => x"00000795",
			482 => x"02096604",
			483 => x"00000795",
			484 => x"00140795",
			485 => x"07069b08",
			486 => x"04129904",
			487 => x"ff2f07b1",
			488 => x"000007b1",
			489 => x"0100ef04",
			490 => x"006f07b1",
			491 => x"000007b1",
			492 => x"020bf304",
			493 => x"fe5307cd",
			494 => x"01011708",
			495 => x"0f0be504",
			496 => x"068607cd",
			497 => x"046a07cd",
			498 => x"fe6007cd",
			499 => x"020bf304",
			500 => x"fe5f07e9",
			501 => x"0100f508",
			502 => x"0f0c0904",
			503 => x"03d607e9",
			504 => x"026407e9",
			505 => x"fe7207e9",
			506 => x"0b068f04",
			507 => x"fef80805",
			508 => x"0100d008",
			509 => x"0507f504",
			510 => x"00000805",
			511 => x"00960805",
			512 => x"00000805",
			513 => x"0c05f504",
			514 => x"ffcb0821",
			515 => x"02096604",
			516 => x"00000821",
			517 => x"0306a504",
			518 => x"00000821",
			519 => x"000f0821",
			520 => x"07060204",
			521 => x"fff5083d",
			522 => x"02096604",
			523 => x"0000083d",
			524 => x"0306a504",
			525 => x"0000083d",
			526 => x"001d083d",
			527 => x"0c05f504",
			528 => x"00000859",
			529 => x"02096604",
			530 => x"00000859",
			531 => x"0d06f904",
			532 => x"00000859",
			533 => x"00180859",
			534 => x"0b063c04",
			535 => x"00000875",
			536 => x"02096604",
			537 => x"00000875",
			538 => x"0f085c04",
			539 => x"00000875",
			540 => x"000d0875",
			541 => x"0b063c04",
			542 => x"00000891",
			543 => x"02096604",
			544 => x"00000891",
			545 => x"0306a504",
			546 => x"00000891",
			547 => x"000f0891",
			548 => x"020bf30c",
			549 => x"07068604",
			550 => x"fe6608b5",
			551 => x"0b06fc04",
			552 => x"02fa08b5",
			553 => x"fe7208b5",
			554 => x"0100f504",
			555 => x"01a008b5",
			556 => x"ff0208b5",
			557 => x"020bf30c",
			558 => x"0a021008",
			559 => x"08029104",
			560 => x"feaf08d9",
			561 => x"019308d9",
			562 => x"fe6908d9",
			563 => x"0100f504",
			564 => x"019008d9",
			565 => x"ff8c08d9",
			566 => x"0c06320c",
			567 => x"020ac304",
			568 => x"fe7308fd",
			569 => x"020ac804",
			570 => x"000008fd",
			571 => x"ffd208fd",
			572 => x"0100de04",
			573 => x"016808fd",
			574 => x"ff1608fd",
			575 => x"0c063208",
			576 => x"0412b204",
			577 => x"fe850921",
			578 => x"00000921",
			579 => x"0100de08",
			580 => x"0006ce04",
			581 => x"013d0921",
			582 => x"00000921",
			583 => x"ff990921",
			584 => x"040f7008",
			585 => x"0f0bc904",
			586 => x"fec60945",
			587 => x"00000945",
			588 => x"0b063c04",
			589 => x"00000945",
			590 => x"01007304",
			591 => x"00000945",
			592 => x"00770945",
			593 => x"0c05f504",
			594 => x"fe8c0969",
			595 => x"0100d008",
			596 => x"07068604",
			597 => x"00000969",
			598 => x"01200969",
			599 => x"0c06dc04",
			600 => x"ff620969",
			601 => x"00000969",
			602 => x"0c05f504",
			603 => x"fead098d",
			604 => x"0100d008",
			605 => x"0f085c04",
			606 => x"0000098d",
			607 => x"00d6098d",
			608 => x"00057a04",
			609 => x"ffb0098d",
			610 => x"0000098d",
			611 => x"040d4204",
			612 => x"fe7809b1",
			613 => x"0c05f504",
			614 => x"ff4f09b1",
			615 => x"0100ef08",
			616 => x"01007304",
			617 => x"000009b1",
			618 => x"014909b1",
			619 => x"000009b1",
			620 => x"040d4204",
			621 => x"fec009d5",
			622 => x"0b063c04",
			623 => x"000009d5",
			624 => x"0100ef08",
			625 => x"01007304",
			626 => x"000009d5",
			627 => x"008709d5",
			628 => x"000009d5",
			629 => x"040d4204",
			630 => x"ff0609f9",
			631 => x"0c05f504",
			632 => x"000009f9",
			633 => x"09019008",
			634 => x"0306a504",
			635 => x"000009f9",
			636 => x"006209f9",
			637 => x"000009f9",
			638 => x"07060204",
			639 => x"ff340a1d",
			640 => x"0100ed0c",
			641 => x"02096604",
			642 => x"00000a1d",
			643 => x"01007304",
			644 => x"00000a1d",
			645 => x"00cc0a1d",
			646 => x"00000a1d",
			647 => x"0c05f504",
			648 => x"ff860a41",
			649 => x"0100ed0c",
			650 => x"06015304",
			651 => x"00000a41",
			652 => x"0006ce04",
			653 => x"00720a41",
			654 => x"00000a41",
			655 => x"00000a41",
			656 => x"0c05f504",
			657 => x"00000a65",
			658 => x"0100ed0c",
			659 => x"0f085c04",
			660 => x"00000a65",
			661 => x"06015304",
			662 => x"00000a65",
			663 => x"00710a65",
			664 => x"00000a65",
			665 => x"020bf310",
			666 => x"0c05f504",
			667 => x"fe640a91",
			668 => x"0100cf08",
			669 => x"03054f04",
			670 => x"ff8c0a91",
			671 => x"03640a91",
			672 => x"fe690a91",
			673 => x"0100f504",
			674 => x"01a80a91",
			675 => x"fec40a91",
			676 => x"0f0bae10",
			677 => x"0c05f504",
			678 => x"fe670abd",
			679 => x"0100cf08",
			680 => x"01007304",
			681 => x"00000abd",
			682 => x"01fa0abd",
			683 => x"fe740abd",
			684 => x"01010b04",
			685 => x"01990abd",
			686 => x"ff050abd",
			687 => x"020bf310",
			688 => x"00058704",
			689 => x"fe690ae9",
			690 => x"0803fa08",
			691 => x"0c045b04",
			692 => x"00000ae9",
			693 => x"01410ae9",
			694 => x"fe980ae9",
			695 => x"01011704",
			696 => x"01920ae9",
			697 => x"ff680ae9",
			698 => x"040df508",
			699 => x"020bf304",
			700 => x"fe6d0b15",
			701 => x"00000b15",
			702 => x"0c05f504",
			703 => x"fed10b15",
			704 => x"0100d408",
			705 => x"01007304",
			706 => x"00000b15",
			707 => x"01850b15",
			708 => x"00000b15",
			709 => x"020bf310",
			710 => x"04118b04",
			711 => x"fe790b41",
			712 => x"0803fa08",
			713 => x"020a2004",
			714 => x"00000b41",
			715 => x"00340b41",
			716 => x"00000b41",
			717 => x"09019004",
			718 => x"01330b41",
			719 => x"00000b41",
			720 => x"0c063210",
			721 => x"020a4604",
			722 => x"fe6c0b75",
			723 => x"00058704",
			724 => x"ff010b75",
			725 => x"0a032c04",
			726 => x"00ed0b75",
			727 => x"00000b75",
			728 => x"0100ed08",
			729 => x"00033504",
			730 => x"00000b75",
			731 => x"018a0b75",
			732 => x"febb0b75",
			733 => x"040d4204",
			734 => x"fe900ba1",
			735 => x"0c05f504",
			736 => x"00000ba1",
			737 => x"0100ef0c",
			738 => x"020a4604",
			739 => x"00000ba1",
			740 => x"0414a404",
			741 => x"00f80ba1",
			742 => x"00000ba1",
			743 => x"00000ba1",
			744 => x"0c05f504",
			745 => x"fe740bd5",
			746 => x"0100d410",
			747 => x"06015304",
			748 => x"00000bd5",
			749 => x"01007304",
			750 => x"00000bd5",
			751 => x"0100d004",
			752 => x"01630bd5",
			753 => x"00000bd5",
			754 => x"0c06dc04",
			755 => x"fee60bd5",
			756 => x"00000bd5",
			757 => x"020bf318",
			758 => x"0c05f504",
			759 => x"fe640c11",
			760 => x"0005870c",
			761 => x"0e08f008",
			762 => x"0f095604",
			763 => x"fe890c11",
			764 => x"03270c11",
			765 => x"fe680c11",
			766 => x"0f06e504",
			767 => x"00000c11",
			768 => x"02ae0c11",
			769 => x"0100f504",
			770 => x"01ac0c11",
			771 => x"fecb0c11",
			772 => x"020bf31c",
			773 => x"0c05f504",
			774 => x"fe630c55",
			775 => x"00058710",
			776 => x"0e08f00c",
			777 => x"03094f04",
			778 => x"fe7e0c55",
			779 => x"0e08e104",
			780 => x"00000c55",
			781 => x"070b0c55",
			782 => x"fe660c55",
			783 => x"0f06e504",
			784 => x"ffd70c55",
			785 => x"040a0c55",
			786 => x"0100f504",
			787 => x"01b60c55",
			788 => x"feb60c55",
			789 => x"020bf320",
			790 => x"0c05f504",
			791 => x"fe640ca3",
			792 => x"00058714",
			793 => x"0b06dd10",
			794 => x"0b06dc04",
			795 => x"fe7a0ca3",
			796 => x"0a021008",
			797 => x"0408f804",
			798 => x"00000ca3",
			799 => x"06900ca3",
			800 => x"ff8a0ca3",
			801 => x"fe680ca3",
			802 => x"0f06e504",
			803 => x"fff20ca3",
			804 => x"03370ca3",
			805 => x"0100f504",
			806 => x"01b10ca3",
			807 => x"fec00ca3",
			808 => x"00000ca5",
			809 => x"00000ca9",
			810 => x"00000cad",
			811 => x"00000cb1",
			812 => x"00000cb5",
			813 => x"00000cb9",
			814 => x"00000cbd",
			815 => x"00000cc1",
			816 => x"00000cc5",
			817 => x"00000cc9",
			818 => x"00000ccd",
			819 => x"00000cd1",
			820 => x"00000cd5",
			821 => x"00000cd9",
			822 => x"00000cdd",
			823 => x"00000ce1",
			824 => x"00000ce5",
			825 => x"00000ce9",
			826 => x"00000ced",
			827 => x"00000cf1",
			828 => x"00000cf5",
			829 => x"00000cf9",
			830 => x"00000cfd",
			831 => x"00000d01",
			832 => x"00000d05",
			833 => x"00000d09",
			834 => x"00000d0d",
			835 => x"00000d11",
			836 => x"00000d15",
			837 => x"00000d19",
			838 => x"00000d1d",
			839 => x"00000d21",
			840 => x"040d4204",
			841 => x"ff420d2d",
			842 => x"00000d2d",
			843 => x"040d4204",
			844 => x"ff860d39",
			845 => x"00000d39",
			846 => x"040d4204",
			847 => x"ffd00d45",
			848 => x"00000d45",
			849 => x"07069b04",
			850 => x"fff10d51",
			851 => x"00000d51",
			852 => x"040d4204",
			853 => x"ffc70d5d",
			854 => x"00000d5d",
			855 => x"07068604",
			856 => x"00000d69",
			857 => x"00000d69",
			858 => x"040f7004",
			859 => x"ffcd0d75",
			860 => x"00000d75",
			861 => x"040f7004",
			862 => x"ffe50d81",
			863 => x"00000d81",
			864 => x"040e2304",
			865 => x"ffeb0d8d",
			866 => x"00000d8d",
			867 => x"040f7004",
			868 => x"ffe20d99",
			869 => x"00000d99",
			870 => x"0c05f504",
			871 => x"00000da5",
			872 => x"00050da5",
			873 => x"020bf304",
			874 => x"fe690db9",
			875 => x"09019004",
			876 => x"01c40db9",
			877 => x"fe9d0db9",
			878 => x"07068604",
			879 => x"ffa70dcd",
			880 => x"0100da04",
			881 => x"00340dcd",
			882 => x"00000dcd",
			883 => x"0c05f504",
			884 => x"00000de1",
			885 => x"0f085c04",
			886 => x"00000de1",
			887 => x"00100de1",
			888 => x"020bf308",
			889 => x"0005a804",
			890 => x"fe970dfd",
			891 => x"00000dfd",
			892 => x"01011704",
			893 => x"00bd0dfd",
			894 => x"00000dfd",
			895 => x"07069b08",
			896 => x"04129904",
			897 => x"ff3a0e19",
			898 => x"00000e19",
			899 => x"0100ef04",
			900 => x"00680e19",
			901 => x"00000e19",
			902 => x"020bf304",
			903 => x"fe570e35",
			904 => x"0100f508",
			905 => x"0601a204",
			906 => x"041a0e35",
			907 => x"02fc0e35",
			908 => x"fe6a0e35",
			909 => x"0c05fc04",
			910 => x"febf0e51",
			911 => x"0100d408",
			912 => x"0414cb04",
			913 => x"00d50e51",
			914 => x"00000e51",
			915 => x"00000e51",
			916 => x"0005080c",
			917 => x"0c06a408",
			918 => x"020cab04",
			919 => x"ff4c0e6d",
			920 => x"00000e6d",
			921 => x"00000e6d",
			922 => x"00000e6d",
			923 => x"0c05f504",
			924 => x"ffd00e89",
			925 => x"02096604",
			926 => x"00000e89",
			927 => x"0306a504",
			928 => x"00000e89",
			929 => x"000d0e89",
			930 => x"0c05f504",
			931 => x"fff30ea5",
			932 => x"02096604",
			933 => x"00000ea5",
			934 => x"0306a504",
			935 => x"00000ea5",
			936 => x"00200ea5",
			937 => x"0c05f504",
			938 => x"00000ec1",
			939 => x"0f085c04",
			940 => x"00000ec1",
			941 => x"02096604",
			942 => x"00000ec1",
			943 => x"00160ec1",
			944 => x"0c05f504",
			945 => x"00000edd",
			946 => x"0f085c04",
			947 => x"00000edd",
			948 => x"02096604",
			949 => x"00000edd",
			950 => x"00110edd",
			951 => x"020bf30c",
			952 => x"0c05f504",
			953 => x"fe620f01",
			954 => x"0c05f604",
			955 => x"00000f01",
			956 => x"fe820f01",
			957 => x"0100f504",
			958 => x"01bc0f01",
			959 => x"fea40f01",
			960 => x"020bf30c",
			961 => x"07068604",
			962 => x"fe660f25",
			963 => x"0b06fc04",
			964 => x"028a0f25",
			965 => x"fe750f25",
			966 => x"0100f504",
			967 => x"019e0f25",
			968 => x"ff110f25",
			969 => x"0c06320c",
			970 => x"020ac304",
			971 => x"fe700f49",
			972 => x"020ac804",
			973 => x"00000f49",
			974 => x"ffc90f49",
			975 => x"0100de04",
			976 => x"017b0f49",
			977 => x"fefa0f49",
			978 => x"0c063208",
			979 => x"0412b204",
			980 => x"fe7f0f6d",
			981 => x"00000f6d",
			982 => x"0100de08",
			983 => x"0006ce04",
			984 => x"01520f6d",
			985 => x"00000f6d",
			986 => x"ff7c0f6d",
			987 => x"07068608",
			988 => x"04129904",
			989 => x"fe8d0f91",
			990 => x"00000f91",
			991 => x"0100ed08",
			992 => x"00033504",
			993 => x"00000f91",
			994 => x"01160f91",
			995 => x"ffec0f91",
			996 => x"07068608",
			997 => x"04129904",
			998 => x"feec0fb5",
			999 => x"00000fb5",
			1000 => x"09018308",
			1001 => x"00033504",
			1002 => x"00000fb5",
			1003 => x"00a90fb5",
			1004 => x"00000fb5",
			1005 => x"0c05f504",
			1006 => x"fea20fd9",
			1007 => x"0100d008",
			1008 => x"0f085c04",
			1009 => x"00000fd9",
			1010 => x"00f30fd9",
			1011 => x"020f1004",
			1012 => x"ff9b0fd9",
			1013 => x"00000fd9",
			1014 => x"0c05fc04",
			1015 => x"feb20ffd",
			1016 => x"09015a08",
			1017 => x"0414cb04",
			1018 => x"00e60ffd",
			1019 => x"00000ffd",
			1020 => x"09018304",
			1021 => x"00000ffd",
			1022 => x"fffa0ffd",
			1023 => x"040d4204",
			1024 => x"fe7c1021",
			1025 => x"0c05f504",
			1026 => x"ff6d1021",
			1027 => x"0100ef08",
			1028 => x"01007304",
			1029 => x"00001021",
			1030 => x"01351021",
			1031 => x"00001021",
			1032 => x"0c05f504",
			1033 => x"fedd1045",
			1034 => x"0100d00c",
			1035 => x"06015304",
			1036 => x"00001045",
			1037 => x"00072404",
			1038 => x"00ac1045",
			1039 => x"00001045",
			1040 => x"00001045",
			1041 => x"040d4204",
			1042 => x"ff101069",
			1043 => x"07060204",
			1044 => x"00001069",
			1045 => x"0100ef08",
			1046 => x"01007304",
			1047 => x"00001069",
			1048 => x"005b1069",
			1049 => x"00001069",
			1050 => x"0c05f504",
			1051 => x"ff3a108d",
			1052 => x"0100ed0c",
			1053 => x"02096604",
			1054 => x"0000108d",
			1055 => x"00072404",
			1056 => x"00c3108d",
			1057 => x"0000108d",
			1058 => x"0000108d",
			1059 => x"0c05f504",
			1060 => x"ff9710b1",
			1061 => x"0100ed0c",
			1062 => x"00033504",
			1063 => x"000010b1",
			1064 => x"01007304",
			1065 => x"000010b1",
			1066 => x"006910b1",
			1067 => x"000010b1",
			1068 => x"020bf310",
			1069 => x"0c05f504",
			1070 => x"fe5e10dd",
			1071 => x"00053e04",
			1072 => x"fe6710dd",
			1073 => x"08050404",
			1074 => x"0da910dd",
			1075 => x"ff1410dd",
			1076 => x"0100f504",
			1077 => x"01fd10dd",
			1078 => x"fe8610dd",
			1079 => x"020bf310",
			1080 => x"0c05f504",
			1081 => x"fe651109",
			1082 => x"0100cf08",
			1083 => x"06015304",
			1084 => x"ffd41109",
			1085 => x"02a91109",
			1086 => x"fe6b1109",
			1087 => x"0100f504",
			1088 => x"01a21109",
			1089 => x"fedd1109",
			1090 => x"020bf310",
			1091 => x"04129904",
			1092 => x"fe681135",
			1093 => x"08040208",
			1094 => x"0207bc04",
			1095 => x"00001135",
			1096 => x"01791135",
			1097 => x"fe8b1135",
			1098 => x"01011704",
			1099 => x"01961135",
			1100 => x"ff4f1135",
			1101 => x"020bf310",
			1102 => x"0a02100c",
			1103 => x"07069b04",
			1104 => x"feba1161",
			1105 => x"0409a004",
			1106 => x"00001161",
			1107 => x"01781161",
			1108 => x"fe6a1161",
			1109 => x"0100f504",
			1110 => x"018d1161",
			1111 => x"ff9a1161",
			1112 => x"020bf310",
			1113 => x"0803be04",
			1114 => x"fe6e118d",
			1115 => x"0c05f504",
			1116 => x"fedd118d",
			1117 => x"020a3a04",
			1118 => x"0000118d",
			1119 => x"0120118d",
			1120 => x"0100f504",
			1121 => x"0177118d",
			1122 => x"ffc2118d",
			1123 => x"07068608",
			1124 => x"04129904",
			1125 => x"fef611b9",
			1126 => x"000011b9",
			1127 => x"0c063204",
			1128 => x"000011b9",
			1129 => x"06022408",
			1130 => x"00033504",
			1131 => x"000011b9",
			1132 => x"004211b9",
			1133 => x"000011b9",
			1134 => x"0c063210",
			1135 => x"020a4604",
			1136 => x"fe6c11ed",
			1137 => x"0412b204",
			1138 => x"ff0b11ed",
			1139 => x"0a033404",
			1140 => x"00d611ed",
			1141 => x"000011ed",
			1142 => x"0100da04",
			1143 => x"018611ed",
			1144 => x"0100ed04",
			1145 => x"000011ed",
			1146 => x"fec711ed",
			1147 => x"040d4204",
			1148 => x"fe941219",
			1149 => x"0c05f504",
			1150 => x"00001219",
			1151 => x"0100ef0c",
			1152 => x"020a4604",
			1153 => x"00001219",
			1154 => x"0414a404",
			1155 => x"00e81219",
			1156 => x"00001219",
			1157 => x"00001219",
			1158 => x"0c05f504",
			1159 => x"fe76124d",
			1160 => x"0100d410",
			1161 => x"06015304",
			1162 => x"0000124d",
			1163 => x"01007304",
			1164 => x"0000124d",
			1165 => x"0100d004",
			1166 => x"0157124d",
			1167 => x"0000124d",
			1168 => x"0c06dc04",
			1169 => x"fef4124d",
			1170 => x"0000124d",
			1171 => x"0f0bae18",
			1172 => x"040f7004",
			1173 => x"fe631289",
			1174 => x"0f085c04",
			1175 => x"fe641289",
			1176 => x"06017304",
			1177 => x"05ff1289",
			1178 => x"0100a104",
			1179 => x"01d71289",
			1180 => x"00051504",
			1181 => x"00001289",
			1182 => x"ff751289",
			1183 => x"0100f504",
			1184 => x"01d91289",
			1185 => x"fe7d1289",
			1186 => x"020bf31c",
			1187 => x"0c05f504",
			1188 => x"fe5c12d5",
			1189 => x"0c05f604",
			1190 => x"ff4012d5",
			1191 => x"0c063a10",
			1192 => x"0c063204",
			1193 => x"fe6e12d5",
			1194 => x"0c063304",
			1195 => x"011112d5",
			1196 => x"0c063404",
			1197 => x"fea412d5",
			1198 => x"000012d5",
			1199 => x"fe5e12d5",
			1200 => x"09019008",
			1201 => x"0f0c0904",
			1202 => x"035112d5",
			1203 => x"023712d5",
			1204 => x"fe7712d5",
			1205 => x"030ba628",
			1206 => x"030b6320",
			1207 => x"06019914",
			1208 => x"0d097510",
			1209 => x"030b2304",
			1210 => x"fe551333",
			1211 => x"030b3208",
			1212 => x"030b2a04",
			1213 => x"ff2c1333",
			1214 => x"ffc61333",
			1215 => x"fe5a1333",
			1216 => x"006f1333",
			1217 => x"0100cd08",
			1218 => x"030a2804",
			1219 => x"feac1333",
			1220 => x"03e91333",
			1221 => x"fe551333",
			1222 => x"00048204",
			1223 => x"fe5d1333",
			1224 => x"038c1333",
			1225 => x"01011304",
			1226 => x"03851333",
			1227 => x"fe5f1333",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(402, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(808, initial_addr_3'length));
	end generate gen_rom_5;

	gen_rom_6: if SELECT_ROM = 6 generate
		bank <= (
			0 => x"00000005",
			1 => x"00000009",
			2 => x"0000000d",
			3 => x"00000011",
			4 => x"00000015",
			5 => x"00000019",
			6 => x"0000001d",
			7 => x"00000021",
			8 => x"00000025",
			9 => x"00000029",
			10 => x"0000002d",
			11 => x"00000031",
			12 => x"00000035",
			13 => x"00000039",
			14 => x"0000003d",
			15 => x"00000041",
			16 => x"00000045",
			17 => x"00000049",
			18 => x"0000004d",
			19 => x"00000051",
			20 => x"00000055",
			21 => x"00000059",
			22 => x"0000005d",
			23 => x"00000061",
			24 => x"00000065",
			25 => x"00000069",
			26 => x"0000006d",
			27 => x"00000071",
			28 => x"00000075",
			29 => x"00000079",
			30 => x"0207f804",
			31 => x"00000085",
			32 => x"fff90085",
			33 => x"03039404",
			34 => x"00000091",
			35 => x"ffd20091",
			36 => x"0207eb04",
			37 => x"0000009d",
			38 => x"ffe8009d",
			39 => x"0207eb04",
			40 => x"000000a9",
			41 => x"fffc00a9",
			42 => x"06013e08",
			43 => x"06011204",
			44 => x"000000bd",
			45 => x"002100bd",
			46 => x"000000bd",
			47 => x"06013e08",
			48 => x"06011204",
			49 => x"000000d1",
			50 => x"001e00d1",
			51 => x"000000d1",
			52 => x"040f7008",
			53 => x"0d063704",
			54 => x"ffa400e5",
			55 => x"000000e5",
			56 => x"000000e5",
			57 => x"06013608",
			58 => x"06011204",
			59 => x"000000f9",
			60 => x"001300f9",
			61 => x"000000f9",
			62 => x"06013e08",
			63 => x"06011204",
			64 => x"0000010d",
			65 => x"0010010d",
			66 => x"0000010d",
			67 => x"0207eb04",
			68 => x"00000121",
			69 => x"0303a004",
			70 => x"00000121",
			71 => x"ffe80121",
			72 => x"06013e08",
			73 => x"06011204",
			74 => x"00000135",
			75 => x"00100135",
			76 => x"00000135",
			77 => x"06013e08",
			78 => x"06011204",
			79 => x"00000149",
			80 => x"001f0149",
			81 => x"00000149",
			82 => x"06013e08",
			83 => x"06011204",
			84 => x"0000015d",
			85 => x"000d015d",
			86 => x"0000015d",
			87 => x"06013e08",
			88 => x"06011204",
			89 => x"00000171",
			90 => x"001b0171",
			91 => x"00000171",
			92 => x"06013508",
			93 => x"06011204",
			94 => x"0000018d",
			95 => x"0018018d",
			96 => x"0207f804",
			97 => x"0000018d",
			98 => x"ffc0018d",
			99 => x"06013e0c",
			100 => x"0207f808",
			101 => x"06011204",
			102 => x"000001a9",
			103 => x"003a01a9",
			104 => x"000001a9",
			105 => x"ffd401a9",
			106 => x"0207f80c",
			107 => x"06013e08",
			108 => x"06011204",
			109 => x"000001cd",
			110 => x"004501cd",
			111 => x"000001cd",
			112 => x"02099d04",
			113 => x"ff9401cd",
			114 => x"000001cd",
			115 => x"0d063708",
			116 => x"03037b04",
			117 => x"000001f1",
			118 => x"ffc301f1",
			119 => x"0e055204",
			120 => x"000001f1",
			121 => x"0e094004",
			122 => x"003b01f1",
			123 => x"000001f1",
			124 => x"040d5504",
			125 => x"ff5b0215",
			126 => x"0c050b0c",
			127 => x"06013e08",
			128 => x"06011f04",
			129 => x"00000215",
			130 => x"006e0215",
			131 => x"00000215",
			132 => x"00000215",
			133 => x"06013e10",
			134 => x"0305f904",
			135 => x"00000239",
			136 => x"06011204",
			137 => x"00000239",
			138 => x"0d063704",
			139 => x"00000239",
			140 => x"00600239",
			141 => x"00000239",
			142 => x"06013510",
			143 => x"06011204",
			144 => x"00000265",
			145 => x"08048f08",
			146 => x"08027904",
			147 => x"00000265",
			148 => x"00270265",
			149 => x"00000265",
			150 => x"03036b04",
			151 => x"00000265",
			152 => x"ffbb0265",
			153 => x"06013610",
			154 => x"0305f908",
			155 => x"0410bb04",
			156 => x"fff20299",
			157 => x"00000299",
			158 => x"040a6904",
			159 => x"00000299",
			160 => x"007c0299",
			161 => x"04120c08",
			162 => x"05065d04",
			163 => x"ff6b0299",
			164 => x"00000299",
			165 => x"00000299",
			166 => x"0e02ea10",
			167 => x"0804d30c",
			168 => x"0f05ad08",
			169 => x"0411ca04",
			170 => x"025202d5",
			171 => x"037e02d5",
			172 => x"fe6602d5",
			173 => x"fe6102d5",
			174 => x"0f05ad0c",
			175 => x"0704aa08",
			176 => x"01002504",
			177 => x"039f02d5",
			178 => x"fe9202d5",
			179 => x"fe5c02d5",
			180 => x"fe5a02d5",
			181 => x"0207f814",
			182 => x"01005c10",
			183 => x"06013e0c",
			184 => x"06011204",
			185 => x"00000309",
			186 => x"00076604",
			187 => x"00280309",
			188 => x"00000309",
			189 => x"00000309",
			190 => x"00000309",
			191 => x"0303a004",
			192 => x"00000309",
			193 => x"ffb40309",
			194 => x"040d5504",
			195 => x"fe7c0335",
			196 => x"06013e10",
			197 => x"07055f0c",
			198 => x"06011904",
			199 => x"00000335",
			200 => x"02090004",
			201 => x"01160335",
			202 => x"00000335",
			203 => x"fff70335",
			204 => x"ff100335",
			205 => x"06013e14",
			206 => x"0d05b504",
			207 => x"00000361",
			208 => x"0207df04",
			209 => x"00000361",
			210 => x"0304c704",
			211 => x"00000361",
			212 => x"0b06cc04",
			213 => x"007a0361",
			214 => x"00000361",
			215 => x"00000361",
			216 => x"01003214",
			217 => x"0505df10",
			218 => x"06013e0c",
			219 => x"06011f04",
			220 => x"000003a5",
			221 => x"0208ad04",
			222 => x"014503a5",
			223 => x"000003a5",
			224 => x"000003a5",
			225 => x"ffbd03a5",
			226 => x"0d067804",
			227 => x"fe8103a5",
			228 => x"0c04ee08",
			229 => x"0e070104",
			230 => x"013d03a5",
			231 => x"000003a5",
			232 => x"fef803a5",
			233 => x"040d5504",
			234 => x"fede03d9",
			235 => x"0c050b14",
			236 => x"0b04c30c",
			237 => x"09003908",
			238 => x"0f05e004",
			239 => x"003a03d9",
			240 => x"000003d9",
			241 => x"ffe603d9",
			242 => x"06014a04",
			243 => x"00c303d9",
			244 => x"000003d9",
			245 => x"000003d9",
			246 => x"040f7018",
			247 => x"08028708",
			248 => x"02098e04",
			249 => x"fee30425",
			250 => x"01db0425",
			251 => x"040d8804",
			252 => x"fe6e0425",
			253 => x"0d063704",
			254 => x"fed00425",
			255 => x"0d06c704",
			256 => x"00f80425",
			257 => x"00000425",
			258 => x"0b05040c",
			259 => x"02089308",
			260 => x"06011904",
			261 => x"00000425",
			262 => x"01780425",
			263 => x"00000425",
			264 => x"feca0425",
			265 => x"0d063718",
			266 => x"040f7008",
			267 => x"0f051204",
			268 => x"00000471",
			269 => x"ff130471",
			270 => x"0208930c",
			271 => x"0a038508",
			272 => x"0a02d404",
			273 => x"00000471",
			274 => x"00370471",
			275 => x"00000471",
			276 => x"00000471",
			277 => x"0a028e0c",
			278 => x"040a6904",
			279 => x"00000471",
			280 => x"0100b704",
			281 => x"00ab0471",
			282 => x"00000471",
			283 => x"00000471",
			284 => x"06013e1c",
			285 => x"0d05b510",
			286 => x"0f05e00c",
			287 => x"040df504",
			288 => x"000004ad",
			289 => x"06011904",
			290 => x"000004ad",
			291 => x"005604ad",
			292 => x"ff4504ad",
			293 => x"09004f04",
			294 => x"000004ad",
			295 => x"040a6904",
			296 => x"000004ad",
			297 => x"013b04ad",
			298 => x"ff1604ad",
			299 => x"06013e1c",
			300 => x"0d05b50c",
			301 => x"0f05da08",
			302 => x"0a02c904",
			303 => x"000004e9",
			304 => x"002d04e9",
			305 => x"ff7d04e9",
			306 => x"040aa904",
			307 => x"000004e9",
			308 => x"09004f04",
			309 => x"000004e9",
			310 => x"06013104",
			311 => x"000004e9",
			312 => x"00b004e9",
			313 => x"ff5404e9",
			314 => x"0601321c",
			315 => x"0303a008",
			316 => x"06011f04",
			317 => x"0000053d",
			318 => x"0087053d",
			319 => x"0305f90c",
			320 => x"0f052f04",
			321 => x"0000053d",
			322 => x"01001704",
			323 => x"0000053d",
			324 => x"ff4c053d",
			325 => x"0a020804",
			326 => x"0000053d",
			327 => x"0098053d",
			328 => x"0506a608",
			329 => x"03036b04",
			330 => x"0000053d",
			331 => x"feb4053d",
			332 => x"0b05c704",
			333 => x"0000053d",
			334 => x"ffac053d",
			335 => x"040d550c",
			336 => x"08028708",
			337 => x"00032c04",
			338 => x"ff410581",
			339 => x"01140581",
			340 => x"fe780581",
			341 => x"06013e14",
			342 => x"07055f10",
			343 => x"06011f04",
			344 => x"00000581",
			345 => x"01003204",
			346 => x"015d0581",
			347 => x"040da904",
			348 => x"00c60581",
			349 => x"ff7b0581",
			350 => x"ffc00581",
			351 => x"fefe0581",
			352 => x"040d5504",
			353 => x"ff6d05b5",
			354 => x"0c050b14",
			355 => x"06013e10",
			356 => x"06011904",
			357 => x"000005b5",
			358 => x"02092e08",
			359 => x"08049304",
			360 => x"006905b5",
			361 => x"000005b5",
			362 => x"000005b5",
			363 => x"000005b5",
			364 => x"000005b5",
			365 => x"06013a1c",
			366 => x"0305f914",
			367 => x"01003210",
			368 => x"0506080c",
			369 => x"06011904",
			370 => x"000005f1",
			371 => x"02089304",
			372 => x"00f205f1",
			373 => x"000005f1",
			374 => x"000005f1",
			375 => x"fedb05f1",
			376 => x"040a6904",
			377 => x"000005f1",
			378 => x"014805f1",
			379 => x"fea205f1",
			380 => x"0b054514",
			381 => x"04112a08",
			382 => x"01002504",
			383 => x"00000645",
			384 => x"fe870645",
			385 => x"02089308",
			386 => x"0804a304",
			387 => x"01010645",
			388 => x"00000645",
			389 => x"00000645",
			390 => x"0c059c14",
			391 => x"0a029310",
			392 => x"040a6904",
			393 => x"00000645",
			394 => x"0100b708",
			395 => x"0c04d104",
			396 => x"00000645",
			397 => x"017b0645",
			398 => x"00000645",
			399 => x"ff990645",
			400 => x"ff300645",
			401 => x"06013e20",
			402 => x"0305f914",
			403 => x"0a02c904",
			404 => x"ff520689",
			405 => x"0100320c",
			406 => x"0505f908",
			407 => x"0f067404",
			408 => x"00970689",
			409 => x"00000689",
			410 => x"00000689",
			411 => x"00000689",
			412 => x"040a6904",
			413 => x"00000689",
			414 => x"0505ce04",
			415 => x"00000689",
			416 => x"00fe0689",
			417 => x"ff2e0689",
			418 => x"06013e20",
			419 => x"0305f914",
			420 => x"01003210",
			421 => x"0505f90c",
			422 => x"02089308",
			423 => x"0a02c904",
			424 => x"000006cd",
			425 => x"006906cd",
			426 => x"000006cd",
			427 => x"000006cd",
			428 => x"ff8806cd",
			429 => x"040a6904",
			430 => x"000006cd",
			431 => x"0505cc04",
			432 => x"000006cd",
			433 => x"00a406cd",
			434 => x"ff7506cd",
			435 => x"0e02ea18",
			436 => x"06013910",
			437 => x"0208930c",
			438 => x"06011904",
			439 => x"00000729",
			440 => x"0804a304",
			441 => x"019d0729",
			442 => x"00000729",
			443 => x"00000729",
			444 => x"06013a04",
			445 => x"00000729",
			446 => x"ff420729",
			447 => x"040d5504",
			448 => x"fe680729",
			449 => x"06013e10",
			450 => x"0e04bb0c",
			451 => x"0207eb08",
			452 => x"040f7004",
			453 => x"ff480729",
			454 => x"01120729",
			455 => x"fec90729",
			456 => x"01e90729",
			457 => x"fe830729",
			458 => x"01003214",
			459 => x"0505df10",
			460 => x"06013e0c",
			461 => x"06011904",
			462 => x"ffc80785",
			463 => x"02089304",
			464 => x"019e0785",
			465 => x"00000785",
			466 => x"ff5c0785",
			467 => x"fec90785",
			468 => x"08028708",
			469 => x"0409ed04",
			470 => x"fec70785",
			471 => x"02d00785",
			472 => x"040d5504",
			473 => x"fe6b0785",
			474 => x"040d6e0c",
			475 => x"0d06e204",
			476 => x"fff20785",
			477 => x"0506c404",
			478 => x"00f90785",
			479 => x"00000785",
			480 => x"fef90785",
			481 => x"040d550c",
			482 => x"08028708",
			483 => x"00033504",
			484 => x"fee707d1",
			485 => x"020807d1",
			486 => x"fe6d07d1",
			487 => x"06013e18",
			488 => x"07055f14",
			489 => x"06011904",
			490 => x"000007d1",
			491 => x"01003608",
			492 => x"02089304",
			493 => x"019507d1",
			494 => x"000007d1",
			495 => x"01004704",
			496 => x"ffbb07d1",
			497 => x"00e907d1",
			498 => x"ff5707d1",
			499 => x"feaf07d1",
			500 => x"0303a010",
			501 => x"06013a0c",
			502 => x"0f05ad08",
			503 => x"0804b204",
			504 => x"02620835",
			505 => x"011e0835",
			506 => x"00090835",
			507 => x"fe780835",
			508 => x"0f05c310",
			509 => x"0505b10c",
			510 => x"01002508",
			511 => x"05051404",
			512 => x"02430835",
			513 => x"03aa0835",
			514 => x"fe930835",
			515 => x"fe610835",
			516 => x"040d5504",
			517 => x"fe5b0835",
			518 => x"06013e0c",
			519 => x"06012b04",
			520 => x"fe660835",
			521 => x"04138704",
			522 => x"0a050835",
			523 => x"fe780835",
			524 => x"fe5d0835",
			525 => x"040d550c",
			526 => x"08028708",
			527 => x"0409db04",
			528 => x"ff520889",
			529 => x"01000889",
			530 => x"fe7a0889",
			531 => x"06013e1c",
			532 => x"07055f18",
			533 => x"0100320c",
			534 => x"06011f04",
			535 => x"00000889",
			536 => x"02089304",
			537 => x"01620889",
			538 => x"00000889",
			539 => x"08035e08",
			540 => x"0600fb04",
			541 => x"00000889",
			542 => x"01290889",
			543 => x"ff3b0889",
			544 => x"ffd40889",
			545 => x"ff0b0889",
			546 => x"0303a00c",
			547 => x"06013a08",
			548 => x"0f05da04",
			549 => x"01ca08fd",
			550 => x"ff9908fd",
			551 => x"fe9b08fd",
			552 => x"0f05e014",
			553 => x"0505b110",
			554 => x"040f7004",
			555 => x"fea808fd",
			556 => x"07049408",
			557 => x"0504f204",
			558 => x"ff9a08fd",
			559 => x"019f08fd",
			560 => x"03da08fd",
			561 => x"fe6b08fd",
			562 => x"040d550c",
			563 => x"06011408",
			564 => x"06011204",
			565 => x"fe7908fd",
			566 => x"01d808fd",
			567 => x"fe6508fd",
			568 => x"06013e0c",
			569 => x"05059204",
			570 => x"fe6708fd",
			571 => x"0b05c704",
			572 => x"065308fd",
			573 => x"fe9d08fd",
			574 => x"fe6508fd",
			575 => x"0303ac14",
			576 => x"06013a10",
			577 => x"06011904",
			578 => x"fe880981",
			579 => x"02089108",
			580 => x"00081204",
			581 => x"01b40981",
			582 => x"ff8c0981",
			583 => x"06250981",
			584 => x"feb50981",
			585 => x"01003220",
			586 => x"0207f80c",
			587 => x"03041608",
			588 => x"06013504",
			589 => x"01440981",
			590 => x"ff440981",
			591 => x"03380981",
			592 => x"09004f0c",
			593 => x"02081b08",
			594 => x"02081504",
			595 => x"ff0d0981",
			596 => x"00c40981",
			597 => x"fe660981",
			598 => x"0c045b04",
			599 => x"00000981",
			600 => x"020e0981",
			601 => x"040d8804",
			602 => x"fe680981",
			603 => x"06013908",
			604 => x"06012404",
			605 => x"00000981",
			606 => x"01810981",
			607 => x"fe6a0981",
			608 => x"040d5510",
			609 => x"0601140c",
			610 => x"0207df04",
			611 => x"000009e5",
			612 => x"0305a704",
			613 => x"000009e5",
			614 => x"004609e5",
			615 => x"fe8809e5",
			616 => x"06013e20",
			617 => x"07055f1c",
			618 => x"040df50c",
			619 => x"08032308",
			620 => x"0a025704",
			621 => x"000009e5",
			622 => x"007f09e5",
			623 => x"ffa909e5",
			624 => x"06011904",
			625 => x"000009e5",
			626 => x"02090008",
			627 => x"08049e04",
			628 => x"011509e5",
			629 => x"000009e5",
			630 => x"000009e5",
			631 => x"000009e5",
			632 => x"ff4009e5",
			633 => x"0303a00c",
			634 => x"06013a08",
			635 => x"06011c04",
			636 => x"00000a61",
			637 => x"01a60a61",
			638 => x"ff090a61",
			639 => x"040d550c",
			640 => x"08028708",
			641 => x"00032c04",
			642 => x"fe780a61",
			643 => x"05b90a61",
			644 => x"fe650a61",
			645 => x"02080918",
			646 => x"06013e14",
			647 => x"0c04b30c",
			648 => x"01003208",
			649 => x"06012304",
			650 => x"00000a61",
			651 => x"01ba0a61",
			652 => x"fee70a61",
			653 => x"01001304",
			654 => x"00000a61",
			655 => x"02cf0a61",
			656 => x"ff1a0a61",
			657 => x"06013a0c",
			658 => x"06013104",
			659 => x"fe920a61",
			660 => x"0414a404",
			661 => x"019a0a61",
			662 => x"ff7d0a61",
			663 => x"fe6d0a61",
			664 => x"0e02f114",
			665 => x"06013a10",
			666 => x"0f05da0c",
			667 => x"0007f608",
			668 => x"04118b04",
			669 => x"00000aed",
			670 => x"01a20aed",
			671 => x"00000aed",
			672 => x"ff820aed",
			673 => x"fefc0aed",
			674 => x"040d550c",
			675 => x"06011408",
			676 => x"06011204",
			677 => x"fea00aed",
			678 => x"00680aed",
			679 => x"fe670aed",
			680 => x"08035b0c",
			681 => x"0305f904",
			682 => x"fffa0aed",
			683 => x"0c052504",
			684 => x"02740aed",
			685 => x"00000aed",
			686 => x"0207df0c",
			687 => x"01002508",
			688 => x"00081204",
			689 => x"01900aed",
			690 => x"00000aed",
			691 => x"ff0d0aed",
			692 => x"06013a0c",
			693 => x"06013904",
			694 => x"feea0aed",
			695 => x"05065004",
			696 => x"00960aed",
			697 => x"00000aed",
			698 => x"fe770aed",
			699 => x"0303ac14",
			700 => x"06013a10",
			701 => x"06011904",
			702 => x"fe7e0b83",
			703 => x"00081208",
			704 => x"02088904",
			705 => x"01d80b83",
			706 => x"00030b83",
			707 => x"ff340b83",
			708 => x"fe7f0b83",
			709 => x"0f05e010",
			710 => x"0d055a0c",
			711 => x"01002a08",
			712 => x"05050304",
			713 => x"00000b83",
			714 => x"02ea0b83",
			715 => x"fea40b83",
			716 => x"fe690b83",
			717 => x"040d550c",
			718 => x"06011408",
			719 => x"06011204",
			720 => x"fe760b83",
			721 => x"01eb0b83",
			722 => x"fe610b83",
			723 => x"0207f808",
			724 => x"06013e04",
			725 => x"019d0b83",
			726 => x"ff7e0b83",
			727 => x"02090010",
			728 => x"0208f708",
			729 => x"04120c04",
			730 => x"fe6d0b83",
			731 => x"ff710b83",
			732 => x"040f0204",
			733 => x"04610b83",
			734 => x"fee70b83",
			735 => x"fe640b83",
			736 => x"00000b85",
			737 => x"00000b89",
			738 => x"00000b8d",
			739 => x"00000b91",
			740 => x"00000b95",
			741 => x"00000b99",
			742 => x"00000b9d",
			743 => x"00000ba1",
			744 => x"00000ba5",
			745 => x"00000ba9",
			746 => x"00000bad",
			747 => x"00000bb1",
			748 => x"00000bb5",
			749 => x"00000bb9",
			750 => x"00000bbd",
			751 => x"00000bc1",
			752 => x"00000bc5",
			753 => x"00000bc9",
			754 => x"00000bcd",
			755 => x"00000bd1",
			756 => x"00000bd5",
			757 => x"00000bd9",
			758 => x"00000bdd",
			759 => x"00000be1",
			760 => x"00000be5",
			761 => x"00000be9",
			762 => x"00000bed",
			763 => x"00000bf1",
			764 => x"00000bf5",
			765 => x"040d5504",
			766 => x"ffab0c01",
			767 => x"00000c01",
			768 => x"0207f804",
			769 => x"00000c0d",
			770 => x"fffa0c0d",
			771 => x"03039404",
			772 => x"00000c19",
			773 => x"ffd80c19",
			774 => x"0207eb04",
			775 => x"00000c25",
			776 => x"ffeb0c25",
			777 => x"06013e08",
			778 => x"06012004",
			779 => x"00000c39",
			780 => x"00140c39",
			781 => x"ffe00c39",
			782 => x"06013e08",
			783 => x"06011204",
			784 => x"00000c4d",
			785 => x"001c0c4d",
			786 => x"00000c4d",
			787 => x"06013e08",
			788 => x"06011204",
			789 => x"00000c61",
			790 => x"00170c61",
			791 => x"00000c61",
			792 => x"040f7008",
			793 => x"0305f904",
			794 => x"ffbe0c75",
			795 => x"00000c75",
			796 => x"00000c75",
			797 => x"06013608",
			798 => x"06011204",
			799 => x"00000c89",
			800 => x"000f0c89",
			801 => x"00000c89",
			802 => x"06013e08",
			803 => x"06011204",
			804 => x"00000c9d",
			805 => x"00110c9d",
			806 => x"00000c9d",
			807 => x"0207eb04",
			808 => x"00000cb1",
			809 => x"0303a004",
			810 => x"00000cb1",
			811 => x"ffea0cb1",
			812 => x"06013e08",
			813 => x"06011204",
			814 => x"00000cc5",
			815 => x"000e0cc5",
			816 => x"00000cc5",
			817 => x"06013e08",
			818 => x"06011204",
			819 => x"00000cd9",
			820 => x"001c0cd9",
			821 => x"00000cd9",
			822 => x"06013e08",
			823 => x"06011204",
			824 => x"00000ced",
			825 => x"000c0ced",
			826 => x"00000ced",
			827 => x"06013e08",
			828 => x"06011204",
			829 => x"00000d01",
			830 => x"00180d01",
			831 => x"00000d01",
			832 => x"04112a0c",
			833 => x"0f051204",
			834 => x"00000d1d",
			835 => x"05064404",
			836 => x"ff290d1d",
			837 => x"00000d1d",
			838 => x"00000d1d",
			839 => x"06013a0c",
			840 => x"06011204",
			841 => x"00000d39",
			842 => x"06013604",
			843 => x"002b0d39",
			844 => x"00000d39",
			845 => x"ffe00d39",
			846 => x"0207f80c",
			847 => x"06013e08",
			848 => x"06011204",
			849 => x"00000d5d",
			850 => x"00410d5d",
			851 => x"00000d5d",
			852 => x"02099d04",
			853 => x"ff9c0d5d",
			854 => x"00000d5d",
			855 => x"06013610",
			856 => x"0305f904",
			857 => x"00000d81",
			858 => x"00033504",
			859 => x"00000d81",
			860 => x"0d060f04",
			861 => x"00000d81",
			862 => x"00630d81",
			863 => x"ff9d0d81",
			864 => x"040d5504",
			865 => x"ff640da5",
			866 => x"0c050b0c",
			867 => x"02090008",
			868 => x"08048f04",
			869 => x"00490da5",
			870 => x"00000da5",
			871 => x"00000da5",
			872 => x"00000da5",
			873 => x"0207f810",
			874 => x"01005c0c",
			875 => x"040a6904",
			876 => x"00000dd1",
			877 => x"0417c304",
			878 => x"000f0dd1",
			879 => x"00000dd1",
			880 => x"00000dd1",
			881 => x"0303a004",
			882 => x"00000dd1",
			883 => x"ffc10dd1",
			884 => x"06013510",
			885 => x"06011204",
			886 => x"00000dfd",
			887 => x"00033504",
			888 => x"00000dfd",
			889 => x"08048f04",
			890 => x"00240dfd",
			891 => x"00000dfd",
			892 => x"03036b04",
			893 => x"00000dfd",
			894 => x"ffc10dfd",
			895 => x"0303a00c",
			896 => x"06013908",
			897 => x"0f05d204",
			898 => x"045a0e31",
			899 => x"fe990e31",
			900 => x"fe670e31",
			901 => x"0f05ad0c",
			902 => x"0505b108",
			903 => x"01002504",
			904 => x"04650e31",
			905 => x"fe840e31",
			906 => x"fe590e31",
			907 => x"fe560e31",
			908 => x"0303a010",
			909 => x"06013a0c",
			910 => x"0f05d208",
			911 => x"0a037204",
			912 => x"02f90e6d",
			913 => x"00ef0e6d",
			914 => x"fec60e6d",
			915 => x"fe670e6d",
			916 => x"0f05ad0c",
			917 => x"0b04b108",
			918 => x"01002504",
			919 => x"02f20e6d",
			920 => x"fe9d0e6d",
			921 => x"fe5e0e6d",
			922 => x"fe5d0e6d",
			923 => x"0207f814",
			924 => x"01005c10",
			925 => x"06013e0c",
			926 => x"06011204",
			927 => x"00000ea1",
			928 => x"0417c304",
			929 => x"00250ea1",
			930 => x"00000ea1",
			931 => x"00000ea1",
			932 => x"00000ea1",
			933 => x"0303a004",
			934 => x"00000ea1",
			935 => x"ffbb0ea1",
			936 => x"040d5504",
			937 => x"fed60ecd",
			938 => x"07054910",
			939 => x"06013e0c",
			940 => x"06011f04",
			941 => x"00000ecd",
			942 => x"08049e04",
			943 => x"00a10ecd",
			944 => x"00000ecd",
			945 => x"00000ecd",
			946 => x"00000ecd",
			947 => x"0303a010",
			948 => x"06013a0c",
			949 => x"0f05d208",
			950 => x"0d051904",
			951 => x"02a00f11",
			952 => x"00bb0f11",
			953 => x"fedb0f11",
			954 => x"fe6f0f11",
			955 => x"0f05ad0c",
			956 => x"0b04b108",
			957 => x"01002504",
			958 => x"02980f11",
			959 => x"fea60f11",
			960 => x"fe600f11",
			961 => x"06013e04",
			962 => x"fe710f11",
			963 => x"fe5a0f11",
			964 => x"040d5508",
			965 => x"06011404",
			966 => x"00000f55",
			967 => x"fec30f55",
			968 => x"0207f810",
			969 => x"06013e0c",
			970 => x"0417c308",
			971 => x"06011c04",
			972 => x"00000f55",
			973 => x"00da0f55",
			974 => x"00000f55",
			975 => x"00000f55",
			976 => x"08034204",
			977 => x"00000f55",
			978 => x"0303a004",
			979 => x"00000f55",
			980 => x"ff9a0f55",
			981 => x"0303940c",
			982 => x"0a038808",
			983 => x"09003004",
			984 => x"06150fa1",
			985 => x"043d0fa1",
			986 => x"fea90fa1",
			987 => x"0303ac0c",
			988 => x"00062f08",
			989 => x"0504f204",
			990 => x"fe840fa1",
			991 => x"07610fa1",
			992 => x"fe5f0fa1",
			993 => x"0f05ad0c",
			994 => x"0b04b108",
			995 => x"09004204",
			996 => x"06360fa1",
			997 => x"fe840fa1",
			998 => x"fe560fa1",
			999 => x"fe520fa1",
			1000 => x"01003214",
			1001 => x"0505df10",
			1002 => x"06013e0c",
			1003 => x"06011f04",
			1004 => x"00000fed",
			1005 => x"02089304",
			1006 => x"01820fed",
			1007 => x"00000fed",
			1008 => x"ffa40fed",
			1009 => x"ff140fed",
			1010 => x"08028708",
			1011 => x"02098e04",
			1012 => x"fefb0fed",
			1013 => x"01770fed",
			1014 => x"0d063704",
			1015 => x"fe710fed",
			1016 => x"0d063804",
			1017 => x"00950fed",
			1018 => x"fed20fed",
			1019 => x"06013a1c",
			1020 => x"0305f910",
			1021 => x"00050804",
			1022 => x"fec81029",
			1023 => x"0207f808",
			1024 => x"0007e504",
			1025 => x"00e71029",
			1026 => x"00001029",
			1027 => x"00001029",
			1028 => x"00033504",
			1029 => x"00001029",
			1030 => x"0d062b04",
			1031 => x"00001029",
			1032 => x"016d1029",
			1033 => x"fe971029",
			1034 => x"06013e1c",
			1035 => x"0d05b510",
			1036 => x"0900420c",
			1037 => x"0f05e008",
			1038 => x"06011904",
			1039 => x"00001065",
			1040 => x"00501065",
			1041 => x"00001065",
			1042 => x"ff4e1065",
			1043 => x"09004f04",
			1044 => x"00001065",
			1045 => x"040a6904",
			1046 => x"00001065",
			1047 => x"012b1065",
			1048 => x"ff211065",
			1049 => x"06013e1c",
			1050 => x"0d05b50c",
			1051 => x"09004208",
			1052 => x"0a02c904",
			1053 => x"000010a1",
			1054 => x"000e10a1",
			1055 => x"ff9b10a1",
			1056 => x"040aa904",
			1057 => x"000010a1",
			1058 => x"09004f04",
			1059 => x"000010a1",
			1060 => x"06013104",
			1061 => x"000010a1",
			1062 => x"009110a1",
			1063 => x"ff6710a1",
			1064 => x"0900621c",
			1065 => x"03037b08",
			1066 => x"0f057204",
			1067 => x"015e10f5",
			1068 => x"000010f5",
			1069 => x"05050e08",
			1070 => x"09002f04",
			1071 => x"000010f5",
			1072 => x"ff3110f5",
			1073 => x"0505df08",
			1074 => x"0a02cc04",
			1075 => x"000010f5",
			1076 => x"013510f5",
			1077 => x"ff5f10f5",
			1078 => x"0d067804",
			1079 => x"fe7410f5",
			1080 => x"06013e08",
			1081 => x"00032c04",
			1082 => x"ffdc10f5",
			1083 => x"01a010f5",
			1084 => x"feb110f5",
			1085 => x"0d06370c",
			1086 => x"0410bb08",
			1087 => x"09003404",
			1088 => x"00001139",
			1089 => x"ff261139",
			1090 => x"00001139",
			1091 => x"0c059c14",
			1092 => x"0a029310",
			1093 => x"040a6904",
			1094 => x"00001139",
			1095 => x"0100b708",
			1096 => x"0c04d104",
			1097 => x"00001139",
			1098 => x"009a1139",
			1099 => x"00001139",
			1100 => x"00001139",
			1101 => x"00001139",
			1102 => x"040d5504",
			1103 => x"fe7e1175",
			1104 => x"0c050b18",
			1105 => x"0d05b510",
			1106 => x"04112a08",
			1107 => x"01002504",
			1108 => x"00001175",
			1109 => x"fef71175",
			1110 => x"0f05e004",
			1111 => x"012d1175",
			1112 => x"00001175",
			1113 => x"02090004",
			1114 => x"015b1175",
			1115 => x"00001175",
			1116 => x"ff4f1175",
			1117 => x"06013e20",
			1118 => x"05059210",
			1119 => x"0f05e00c",
			1120 => x"0a02c904",
			1121 => x"000011b9",
			1122 => x"06011c04",
			1123 => x"000011b9",
			1124 => x"00bc11b9",
			1125 => x"fef111b9",
			1126 => x"040a6904",
			1127 => x"000011b9",
			1128 => x"01002d04",
			1129 => x"000011b9",
			1130 => x"0b04f104",
			1131 => x"000011b9",
			1132 => x"015311b9",
			1133 => x"fec811b9",
			1134 => x"0e02d910",
			1135 => x"0f05da0c",
			1136 => x"04117604",
			1137 => x"0000120d",
			1138 => x"0a038804",
			1139 => x"00a0120d",
			1140 => x"0000120d",
			1141 => x"0000120d",
			1142 => x"0d067808",
			1143 => x"01002304",
			1144 => x"0000120d",
			1145 => x"fea1120d",
			1146 => x"0c059c10",
			1147 => x"0a02750c",
			1148 => x"040aa904",
			1149 => x"0000120d",
			1150 => x"0100da04",
			1151 => x"00f7120d",
			1152 => x"0000120d",
			1153 => x"0000120d",
			1154 => x"ff96120d",
			1155 => x"06013e20",
			1156 => x"0305f914",
			1157 => x"0a02c904",
			1158 => x"ff5c1251",
			1159 => x"0207f80c",
			1160 => x"040f7004",
			1161 => x"00001251",
			1162 => x"00076604",
			1163 => x"007b1251",
			1164 => x"00001251",
			1165 => x"00001251",
			1166 => x"040a6904",
			1167 => x"00001251",
			1168 => x"0505ce04",
			1169 => x"00001251",
			1170 => x"00f11251",
			1171 => x"ff381251",
			1172 => x"0303a00c",
			1173 => x"0804d308",
			1174 => x"06011c04",
			1175 => x"00f212ad",
			1176 => x"023512ad",
			1177 => x"fe8112ad",
			1178 => x"0f05c310",
			1179 => x"0c04b90c",
			1180 => x"04100804",
			1181 => x"fe9c12ad",
			1182 => x"06013004",
			1183 => x"020f12ad",
			1184 => x"037912ad",
			1185 => x"fe6312ad",
			1186 => x"040d5504",
			1187 => x"fe5d12ad",
			1188 => x"06013e0c",
			1189 => x"06012b04",
			1190 => x"fe6912ad",
			1191 => x"04138704",
			1192 => x"051112ad",
			1193 => x"fe7f12ad",
			1194 => x"fe5f12ad",
			1195 => x"0e02ea18",
			1196 => x"06013910",
			1197 => x"0f05da0c",
			1198 => x"04117604",
			1199 => x"00001309",
			1200 => x"0804a304",
			1201 => x"019a1309",
			1202 => x"00001309",
			1203 => x"ffd31309",
			1204 => x"06013a04",
			1205 => x"00001309",
			1206 => x"ff551309",
			1207 => x"040d5504",
			1208 => x"fe681309",
			1209 => x"06013e10",
			1210 => x"03054f0c",
			1211 => x"0f05c308",
			1212 => x"04151804",
			1213 => x"00fa1309",
			1214 => x"00001309",
			1215 => x"febc1309",
			1216 => x"01cf1309",
			1217 => x"fe881309",
			1218 => x"0d063718",
			1219 => x"0410bb08",
			1220 => x"01002104",
			1221 => x"00001365",
			1222 => x"fe9a1365",
			1223 => x"0208930c",
			1224 => x"04112a04",
			1225 => x"00001365",
			1226 => x"0505ea04",
			1227 => x"00cc1365",
			1228 => x"00001365",
			1229 => x"00001365",
			1230 => x"0c059c14",
			1231 => x"0a029310",
			1232 => x"040a6904",
			1233 => x"00001365",
			1234 => x"0100b708",
			1235 => x"0c04d104",
			1236 => x"00001365",
			1237 => x"012e1365",
			1238 => x"00001365",
			1239 => x"00001365",
			1240 => x"ff9f1365",
			1241 => x"040d550c",
			1242 => x"08028708",
			1243 => x"00032404",
			1244 => x"ff2313b1",
			1245 => x"017713b1",
			1246 => x"fe7213b1",
			1247 => x"06013e18",
			1248 => x"07055f14",
			1249 => x"06011904",
			1250 => x"000013b1",
			1251 => x"01003208",
			1252 => x"02089304",
			1253 => x"018313b1",
			1254 => x"000013b1",
			1255 => x"01004704",
			1256 => x"ffaa13b1",
			1257 => x"00cd13b1",
			1258 => x"fff513b1",
			1259 => x"fed013b1",
			1260 => x"01003214",
			1261 => x"0505df10",
			1262 => x"040f7004",
			1263 => x"ffcf1415",
			1264 => x"0a02cc04",
			1265 => x"00001415",
			1266 => x"0f067404",
			1267 => x"01671415",
			1268 => x"00001415",
			1269 => x"ff001415",
			1270 => x"0802870c",
			1271 => x"0f098b04",
			1272 => x"fef01415",
			1273 => x"0d088d04",
			1274 => x"01aa1415",
			1275 => x"00001415",
			1276 => x"040d8804",
			1277 => x"fe6f1415",
			1278 => x"040da904",
			1279 => x"004e1415",
			1280 => x"040e2308",
			1281 => x"040df504",
			1282 => x"ffeb1415",
			1283 => x"00001415",
			1284 => x"feed1415",
			1285 => x"0303a00c",
			1286 => x"06013a08",
			1287 => x"06011c04",
			1288 => x"00001481",
			1289 => x"01a91481",
			1290 => x"fefa1481",
			1291 => x"040d550c",
			1292 => x"08028708",
			1293 => x"0409ed04",
			1294 => x"fe751481",
			1295 => x"08711481",
			1296 => x"fe651481",
			1297 => x"02080910",
			1298 => x"0b04bf08",
			1299 => x"0f05b604",
			1300 => x"01581481",
			1301 => x"feb81481",
			1302 => x"09002304",
			1303 => x"ff641481",
			1304 => x"02f71481",
			1305 => x"06013a0c",
			1306 => x"06013104",
			1307 => x"fe881481",
			1308 => x"0414a404",
			1309 => x"01cd1481",
			1310 => x"ff601481",
			1311 => x"fe6b1481",
			1312 => x"0303a010",
			1313 => x"06013908",
			1314 => x"06011c04",
			1315 => x"000014f5",
			1316 => x"01a314f5",
			1317 => x"03039404",
			1318 => x"000014f5",
			1319 => x"ff0014f5",
			1320 => x"040d550c",
			1321 => x"00033e08",
			1322 => x"040a2804",
			1323 => x"fe7714f5",
			1324 => x"046414f5",
			1325 => x"fe6614f5",
			1326 => x"00042d08",
			1327 => x"0c052e04",
			1328 => x"034414f5",
			1329 => x"000014f5",
			1330 => x"06013a14",
			1331 => x"06013008",
			1332 => x"0f05b604",
			1333 => x"008814f5",
			1334 => x"fe9414f5",
			1335 => x"07057308",
			1336 => x"0704a504",
			1337 => x"000014f5",
			1338 => x"01ca14f5",
			1339 => x"ff3b14f5",
			1340 => x"fe6f14f5",
			1341 => x"0303a014",
			1342 => x"0601390c",
			1343 => x"06011c04",
			1344 => x"00001569",
			1345 => x"0a036704",
			1346 => x"01a41569",
			1347 => x"00001569",
			1348 => x"03039404",
			1349 => x"00001569",
			1350 => x"ff0e1569",
			1351 => x"06013e24",
			1352 => x"0d067818",
			1353 => x"0a02e408",
			1354 => x"0f054604",
			1355 => x"00001569",
			1356 => x"fe681569",
			1357 => x"0005ea0c",
			1358 => x"0f05ee04",
			1359 => x"01661569",
			1360 => x"0f066d04",
			1361 => x"ff8b1569",
			1362 => x"00cd1569",
			1363 => x"ff7b1569",
			1364 => x"00033504",
			1365 => x"fe911569",
			1366 => x"0f06d904",
			1367 => x"ff701569",
			1368 => x"03641569",
			1369 => x"fe671569",
			1370 => x"0303ac18",
			1371 => x"06011904",
			1372 => x"fe9d15e5",
			1373 => x"06013a10",
			1374 => x"0419260c",
			1375 => x"0f05e608",
			1376 => x"0d050d04",
			1377 => x"01aa15e5",
			1378 => x"02fc15e5",
			1379 => x"000015e5",
			1380 => x"ffd415e5",
			1381 => x"fece15e5",
			1382 => x"0f05e010",
			1383 => x"0c04b90c",
			1384 => x"01002a08",
			1385 => x"06012304",
			1386 => x"000015e5",
			1387 => x"022b15e5",
			1388 => x"feda15e5",
			1389 => x"fe7915e5",
			1390 => x"040d8804",
			1391 => x"fe6a15e5",
			1392 => x"06013e10",
			1393 => x"09004f04",
			1394 => x"fe7615e5",
			1395 => x"0f065904",
			1396 => x"fea615e5",
			1397 => x"06011404",
			1398 => x"000015e5",
			1399 => x"02d515e5",
			1400 => x"fe6c15e5",
			1401 => x"0303ac14",
			1402 => x"0804d310",
			1403 => x"04112a04",
			1404 => x"ff141669",
			1405 => x"0f05da08",
			1406 => x"0b049d04",
			1407 => x"01ae1669",
			1408 => x"03031669",
			1409 => x"ff711669",
			1410 => x"fece1669",
			1411 => x"0f05e010",
			1412 => x"0c04b90c",
			1413 => x"01002a08",
			1414 => x"0c045904",
			1415 => x"00001669",
			1416 => x"02491669",
			1417 => x"fed01669",
			1418 => x"fe751669",
			1419 => x"040d8804",
			1420 => x"fe691669",
			1421 => x"040da90c",
			1422 => x"09009504",
			1423 => x"ff1b1669",
			1424 => x"01008804",
			1425 => x"03311669",
			1426 => x"00001669",
			1427 => x"040e230c",
			1428 => x"0900c204",
			1429 => x"feaa1669",
			1430 => x"09015c04",
			1431 => x"01901669",
			1432 => x"ff511669",
			1433 => x"fe971669",
			1434 => x"0e02ea14",
			1435 => x"06013a10",
			1436 => x"06011904",
			1437 => x"ffc816e5",
			1438 => x"0208ab08",
			1439 => x"0007f604",
			1440 => x"01a016e5",
			1441 => x"000016e5",
			1442 => x"000016e5",
			1443 => x"ff2216e5",
			1444 => x"040d550c",
			1445 => x"06011408",
			1446 => x"06011204",
			1447 => x"fea816e5",
			1448 => x"005316e5",
			1449 => x"fe6716e5",
			1450 => x"06013e1c",
			1451 => x"0e04bb18",
			1452 => x"0410bb0c",
			1453 => x"03041d08",
			1454 => x"0e032004",
			1455 => x"000016e5",
			1456 => x"001f16e5",
			1457 => x"feae16e5",
			1458 => x"05061508",
			1459 => x"07047e04",
			1460 => x"000016e5",
			1461 => x"019216e5",
			1462 => x"ff3816e5",
			1463 => x"024216e5",
			1464 => x"fe7a16e5",
			1465 => x"0303a010",
			1466 => x"06013a0c",
			1467 => x"0f05da08",
			1468 => x"0c04ce04",
			1469 => x"01b9177b",
			1470 => x"0083177b",
			1471 => x"ffe8177b",
			1472 => x"feae177b",
			1473 => x"0f05e014",
			1474 => x"0505b110",
			1475 => x"040f7004",
			1476 => x"febb177b",
			1477 => x"0504f204",
			1478 => x"ffd7177b",
			1479 => x"0f058504",
			1480 => x"017a177b",
			1481 => x"0333177b",
			1482 => x"fe6f177b",
			1483 => x"040d550c",
			1484 => x"06011408",
			1485 => x"06011204",
			1486 => x"fe82177b",
			1487 => x"0176177b",
			1488 => x"fe67177b",
			1489 => x"08035b0c",
			1490 => x"01005804",
			1491 => x"fed4177b",
			1492 => x"0b05c704",
			1493 => x"042d177b",
			1494 => x"ff2d177b",
			1495 => x"06013e0c",
			1496 => x"05059204",
			1497 => x"fe72177b",
			1498 => x"05067904",
			1499 => x"028e177b",
			1500 => x"feb6177b",
			1501 => x"fe67177b",
			1502 => x"0000177d",
			1503 => x"00001781",
			1504 => x"00001785",
			1505 => x"00001789",
			1506 => x"0000178d",
			1507 => x"00001791",
			1508 => x"00001795",
			1509 => x"00001799",
			1510 => x"0000179d",
			1511 => x"000017a1",
			1512 => x"000017a5",
			1513 => x"000017a9",
			1514 => x"000017ad",
			1515 => x"000017b1",
			1516 => x"000017b5",
			1517 => x"000017b9",
			1518 => x"000017bd",
			1519 => x"000017c1",
			1520 => x"000017c5",
			1521 => x"000017c9",
			1522 => x"000017cd",
			1523 => x"000017d1",
			1524 => x"000017d5",
			1525 => x"000017d9",
			1526 => x"000017dd",
			1527 => x"000017e1",
			1528 => x"000017e5",
			1529 => x"000017e9",
			1530 => x"000017ed",
			1531 => x"0207f804",
			1532 => x"000017f9",
			1533 => x"fff617f9",
			1534 => x"0e02af04",
			1535 => x"00001805",
			1536 => x"ffd71805",
			1537 => x"0207eb04",
			1538 => x"00001811",
			1539 => x"ffe61811",
			1540 => x"0207eb04",
			1541 => x"0000181d",
			1542 => x"fff9181d",
			1543 => x"06013e08",
			1544 => x"06012004",
			1545 => x"00001831",
			1546 => x"00131831",
			1547 => x"ffe61831",
			1548 => x"01003204",
			1549 => x"00001845",
			1550 => x"0d063704",
			1551 => x"ff881845",
			1552 => x"00001845",
			1553 => x"06013e08",
			1554 => x"06011204",
			1555 => x"00001859",
			1556 => x"00161859",
			1557 => x"00001859",
			1558 => x"040f7008",
			1559 => x"0305f904",
			1560 => x"ffc5186d",
			1561 => x"0000186d",
			1562 => x"0000186d",
			1563 => x"06013608",
			1564 => x"06011204",
			1565 => x"00001881",
			1566 => x"000f1881",
			1567 => x"00001881",
			1568 => x"0207eb04",
			1569 => x"00001895",
			1570 => x"0303a004",
			1571 => x"00001895",
			1572 => x"ffe41895",
			1573 => x"06013e08",
			1574 => x"06011204",
			1575 => x"000018a9",
			1576 => x"000f18a9",
			1577 => x"000018a9",
			1578 => x"06013e08",
			1579 => x"06011204",
			1580 => x"000018bd",
			1581 => x"002218bd",
			1582 => x"000018bd",
			1583 => x"06013e08",
			1584 => x"06011204",
			1585 => x"000018d1",
			1586 => x"000f18d1",
			1587 => x"000018d1",
			1588 => x"06013e08",
			1589 => x"06011204",
			1590 => x"000018e5",
			1591 => x"001d18e5",
			1592 => x"000018e5",
			1593 => x"0207f808",
			1594 => x"02078004",
			1595 => x"00001901",
			1596 => x"000d1901",
			1597 => x"02099d04",
			1598 => x"ffb51901",
			1599 => x"00001901",
			1600 => x"04112a0c",
			1601 => x"0f051204",
			1602 => x"0000191d",
			1603 => x"05064404",
			1604 => x"ff3c191d",
			1605 => x"0000191d",
			1606 => x"0000191d",
			1607 => x"06013a0c",
			1608 => x"06011204",
			1609 => x"00001939",
			1610 => x"06013604",
			1611 => x"00271939",
			1612 => x"00001939",
			1613 => x"ffe21939",
			1614 => x"0207f80c",
			1615 => x"06011204",
			1616 => x"0000195d",
			1617 => x"06013e04",
			1618 => x"0022195d",
			1619 => x"0000195d",
			1620 => x"02099d04",
			1621 => x"ffbe195d",
			1622 => x"0000195d",
			1623 => x"04112a10",
			1624 => x"02069d04",
			1625 => x"00001981",
			1626 => x"0b058308",
			1627 => x"01001d04",
			1628 => x"00001981",
			1629 => x"ff351981",
			1630 => x"00001981",
			1631 => x"00001981",
			1632 => x"040d5504",
			1633 => x"ffa419a5",
			1634 => x"0705450c",
			1635 => x"06013e08",
			1636 => x"06011904",
			1637 => x"000019a5",
			1638 => x"003219a5",
			1639 => x"000019a5",
			1640 => x"000019a5",
			1641 => x"06013510",
			1642 => x"040a6904",
			1643 => x"000019d1",
			1644 => x"06011204",
			1645 => x"000019d1",
			1646 => x"08048f04",
			1647 => x"002f19d1",
			1648 => x"000019d1",
			1649 => x"04120c04",
			1650 => x"ffa919d1",
			1651 => x"000019d1",
			1652 => x"0d063708",
			1653 => x"03037b04",
			1654 => x"000019fd",
			1655 => x"ffbf19fd",
			1656 => x"06013e0c",
			1657 => x"0305f904",
			1658 => x"000019fd",
			1659 => x"06011204",
			1660 => x"000019fd",
			1661 => x"006d19fd",
			1662 => x"000019fd",
			1663 => x"040d550c",
			1664 => x"08028708",
			1665 => x"0409ed04",
			1666 => x"fed41a31",
			1667 => x"02691a31",
			1668 => x"fe6c1a31",
			1669 => x"06013e0c",
			1670 => x"07055f08",
			1671 => x"06011904",
			1672 => x"ffe81a31",
			1673 => x"01771a31",
			1674 => x"ff341a31",
			1675 => x"fe9e1a31",
			1676 => x"040d5508",
			1677 => x"06011404",
			1678 => x"00001a65",
			1679 => x"fed21a65",
			1680 => x"06013e10",
			1681 => x"0c05250c",
			1682 => x"06011f04",
			1683 => x"00001a65",
			1684 => x"08049e04",
			1685 => x"00c71a65",
			1686 => x"00001a65",
			1687 => x"00001a65",
			1688 => x"00001a65",
			1689 => x"040d5504",
			1690 => x"fe7a1a91",
			1691 => x"06013e10",
			1692 => x"07055f0c",
			1693 => x"06011904",
			1694 => x"00001a91",
			1695 => x"02090004",
			1696 => x"01291a91",
			1697 => x"00001a91",
			1698 => x"ffeb1a91",
			1699 => x"ff051a91",
			1700 => x"040d5504",
			1701 => x"fee71abd",
			1702 => x"0c050b10",
			1703 => x"06013e0c",
			1704 => x"06011f04",
			1705 => x"00001abd",
			1706 => x"08049e04",
			1707 => x"00931abd",
			1708 => x"00001abd",
			1709 => x"00001abd",
			1710 => x"00001abd",
			1711 => x"03039408",
			1712 => x"06013a04",
			1713 => x"eca31af9",
			1714 => x"d3311af9",
			1715 => x"0303a008",
			1716 => x"0005ff04",
			1717 => x"e5fe1af9",
			1718 => x"d2e11af9",
			1719 => x"0f05ad0c",
			1720 => x"0b04b108",
			1721 => x"01002504",
			1722 => x"ebb91af9",
			1723 => x"d3011af9",
			1724 => x"d2d41af9",
			1725 => x"d2d51af9",
			1726 => x"040d5508",
			1727 => x"06011404",
			1728 => x"00001b3d",
			1729 => x"fecb1b3d",
			1730 => x"0207f810",
			1731 => x"06013e0c",
			1732 => x"00076608",
			1733 => x"06011c04",
			1734 => x"00001b3d",
			1735 => x"00ce1b3d",
			1736 => x"00001b3d",
			1737 => x"00001b3d",
			1738 => x"08034204",
			1739 => x"00001b3d",
			1740 => x"0303a004",
			1741 => x"00001b3d",
			1742 => x"ffa71b3d",
			1743 => x"01003214",
			1744 => x"0505df10",
			1745 => x"06013e0c",
			1746 => x"06011904",
			1747 => x"ff8b1b89",
			1748 => x"02089304",
			1749 => x"01a71b89",
			1750 => x"00001b89",
			1751 => x"ff4f1b89",
			1752 => x"feae1b89",
			1753 => x"08028708",
			1754 => x"0409ed04",
			1755 => x"feb21b89",
			1756 => x"03c41b89",
			1757 => x"040d5504",
			1758 => x"fe6a1b89",
			1759 => x"040d6e04",
			1760 => x"00351b89",
			1761 => x"fee61b89",
			1762 => x"040d550c",
			1763 => x"08028708",
			1764 => x"0409db04",
			1765 => x"00001bd5",
			1766 => x"00ab1bd5",
			1767 => x"febb1bd5",
			1768 => x"0e047810",
			1769 => x"0f05e00c",
			1770 => x"0505ea08",
			1771 => x"01002704",
			1772 => x"00981bd5",
			1773 => x"00001bd5",
			1774 => x"00001bd5",
			1775 => x"ff921bd5",
			1776 => x"0208f908",
			1777 => x"0803b404",
			1778 => x"01171bd5",
			1779 => x"00001bd5",
			1780 => x"00001bd5",
			1781 => x"06013e1c",
			1782 => x"0d05b510",
			1783 => x"0f05e00c",
			1784 => x"0a02c904",
			1785 => x"00001c11",
			1786 => x"06011c04",
			1787 => x"00001c11",
			1788 => x"00ac1c11",
			1789 => x"ff021c11",
			1790 => x"040a6904",
			1791 => x"00001c11",
			1792 => x"04117604",
			1793 => x"013f1c11",
			1794 => x"00001c11",
			1795 => x"fed71c11",
			1796 => x"06013e1c",
			1797 => x"0d05b510",
			1798 => x"0f05da0c",
			1799 => x"09004208",
			1800 => x"06011904",
			1801 => x"00001c4d",
			1802 => x"00401c4d",
			1803 => x"00001c4d",
			1804 => x"ff6b1c4d",
			1805 => x"09004f04",
			1806 => x"00001c4d",
			1807 => x"040a6904",
			1808 => x"00001c4d",
			1809 => x"00ff1c4d",
			1810 => x"ff431c4d",
			1811 => x"040d550c",
			1812 => x"08028708",
			1813 => x"00032c04",
			1814 => x"ff351ca1",
			1815 => x"012d1ca1",
			1816 => x"fe761ca1",
			1817 => x"0207f810",
			1818 => x"040f7008",
			1819 => x"0004d204",
			1820 => x"00761ca1",
			1821 => x"ffae1ca1",
			1822 => x"00076604",
			1823 => x"015c1ca1",
			1824 => x"00001ca1",
			1825 => x"00042508",
			1826 => x"0d06e204",
			1827 => x"00001ca1",
			1828 => x"00921ca1",
			1829 => x"0303a004",
			1830 => x"00001ca1",
			1831 => x"ff121ca1",
			1832 => x"06013220",
			1833 => x"0303a00c",
			1834 => x"06011f04",
			1835 => x"00001cfd",
			1836 => x"0006ad04",
			1837 => x"007b1cfd",
			1838 => x"00001cfd",
			1839 => x"0305f90c",
			1840 => x"0f052f04",
			1841 => x"00001cfd",
			1842 => x"01001704",
			1843 => x"00001cfd",
			1844 => x"ff561cfd",
			1845 => x"00033504",
			1846 => x"00001cfd",
			1847 => x"00911cfd",
			1848 => x"0d06e208",
			1849 => x"03036b04",
			1850 => x"00001cfd",
			1851 => x"febb1cfd",
			1852 => x"0506a704",
			1853 => x"00001cfd",
			1854 => x"ffbd1cfd",
			1855 => x"040d550c",
			1856 => x"08028708",
			1857 => x"0409ed04",
			1858 => x"ff4c1d49",
			1859 => x"012c1d49",
			1860 => x"fe741d49",
			1861 => x"0c050b18",
			1862 => x"040f700c",
			1863 => x"07051a08",
			1864 => x"01002104",
			1865 => x"00001d49",
			1866 => x"ff031d49",
			1867 => x"01261d49",
			1868 => x"02089308",
			1869 => x"0a02cc04",
			1870 => x"00001d49",
			1871 => x"014b1d49",
			1872 => x"00001d49",
			1873 => x"ff121d49",
			1874 => x"06013a1c",
			1875 => x"0305f914",
			1876 => x"01003210",
			1877 => x"0506080c",
			1878 => x"06011904",
			1879 => x"00001d85",
			1880 => x"02089304",
			1881 => x"01001d85",
			1882 => x"00001d85",
			1883 => x"00001d85",
			1884 => x"fed31d85",
			1885 => x"040a6904",
			1886 => x"00001d85",
			1887 => x"01571d85",
			1888 => x"fe9d1d85",
			1889 => x"06013e20",
			1890 => x"0d05b510",
			1891 => x"0900420c",
			1892 => x"02089308",
			1893 => x"0a02c904",
			1894 => x"00001dc9",
			1895 => x"00291dc9",
			1896 => x"00001dc9",
			1897 => x"ff951dc9",
			1898 => x"040aa904",
			1899 => x"00001dc9",
			1900 => x"09004f04",
			1901 => x"00001dc9",
			1902 => x"06013104",
			1903 => x"00001dc9",
			1904 => x"009d1dc9",
			1905 => x"ff5e1dc9",
			1906 => x"06013e20",
			1907 => x"0d05b514",
			1908 => x"0f05e010",
			1909 => x"0a02c904",
			1910 => x"00001e0d",
			1911 => x"06013508",
			1912 => x"06011c04",
			1913 => x"00001e0d",
			1914 => x"00511e0d",
			1915 => x"00001e0d",
			1916 => x"ff3c1e0d",
			1917 => x"09004f04",
			1918 => x"00001e0d",
			1919 => x"040a6904",
			1920 => x"00001e0d",
			1921 => x"014b1e0d",
			1922 => x"ff0b1e0d",
			1923 => x"06013e20",
			1924 => x"0305f914",
			1925 => x"01003210",
			1926 => x"0505f90c",
			1927 => x"02089308",
			1928 => x"0a02c904",
			1929 => x"00001e51",
			1930 => x"00741e51",
			1931 => x"00001e51",
			1932 => x"00001e51",
			1933 => x"ff741e51",
			1934 => x"00033504",
			1935 => x"00001e51",
			1936 => x"0d062b04",
			1937 => x"00001e51",
			1938 => x"00bb1e51",
			1939 => x"ff631e51",
			1940 => x"0e02ea0c",
			1941 => x"0a03aa08",
			1942 => x"0f05b604",
			1943 => x"02131ead",
			1944 => x"fe7f1ead",
			1945 => x"fe741ead",
			1946 => x"0f05c310",
			1947 => x"0c04b90c",
			1948 => x"0410e104",
			1949 => x"fe611ead",
			1950 => x"07049304",
			1951 => x"02001ead",
			1952 => x"03431ead",
			1953 => x"fe661ead",
			1954 => x"040d5504",
			1955 => x"fe5e1ead",
			1956 => x"06013e0c",
			1957 => x"06012b04",
			1958 => x"fe6f1ead",
			1959 => x"04138704",
			1960 => x"03751ead",
			1961 => x"fe861ead",
			1962 => x"fe601ead",
			1963 => x"0e02ea18",
			1964 => x"06013910",
			1965 => x"0f05da0c",
			1966 => x"06011c04",
			1967 => x"00001f09",
			1968 => x"0804a304",
			1969 => x"01981f09",
			1970 => x"00001f09",
			1971 => x"ffed1f09",
			1972 => x"06013a04",
			1973 => x"00001f09",
			1974 => x"ff6a1f09",
			1975 => x"040d5504",
			1976 => x"fe691f09",
			1977 => x"06013e10",
			1978 => x"0e04bb0c",
			1979 => x"0f05c308",
			1980 => x"04151804",
			1981 => x"00e51f09",
			1982 => x"00001f09",
			1983 => x"fec81f09",
			1984 => x"01b61f09",
			1985 => x"fe8d1f09",
			1986 => x"040d550c",
			1987 => x"08028708",
			1988 => x"00033504",
			1989 => x"fedb1f55",
			1990 => x"02471f55",
			1991 => x"fe6c1f55",
			1992 => x"06013e18",
			1993 => x"07055f14",
			1994 => x"06011904",
			1995 => x"00001f55",
			1996 => x"01003608",
			1997 => x"02089304",
			1998 => x"01991f55",
			1999 => x"00001f55",
			2000 => x"01004704",
			2001 => x"ffaf1f55",
			2002 => x"00fd1f55",
			2003 => x"ff431f55",
			2004 => x"fea61f55",
			2005 => x"06013a24",
			2006 => x"0305f918",
			2007 => x"04100808",
			2008 => x"09003604",
			2009 => x"00001fa1",
			2010 => x"febe1fa1",
			2011 => x"0505f90c",
			2012 => x"06011f04",
			2013 => x"00001fa1",
			2014 => x"0006ad04",
			2015 => x"01051fa1",
			2016 => x"00001fa1",
			2017 => x"00001fa1",
			2018 => x"040a6904",
			2019 => x"00001fa1",
			2020 => x"0d061104",
			2021 => x"00001fa1",
			2022 => x"017f1fa1",
			2023 => x"fe931fa1",
			2024 => x"0303a010",
			2025 => x"0411de04",
			2026 => x"ff6a1ffd",
			2027 => x"0a038808",
			2028 => x"06011c04",
			2029 => x"00001ffd",
			2030 => x"01901ffd",
			2031 => x"00001ffd",
			2032 => x"0a021008",
			2033 => x"040a6904",
			2034 => x"febd1ffd",
			2035 => x"03501ffd",
			2036 => x"040d5504",
			2037 => x"fe6b1ffd",
			2038 => x"06013e10",
			2039 => x"0e04780c",
			2040 => x"0f05d208",
			2041 => x"0207e504",
			2042 => x"00fe1ffd",
			2043 => x"00001ffd",
			2044 => x"fec51ffd",
			2045 => x"01c51ffd",
			2046 => x"fe961ffd",
			2047 => x"040d5510",
			2048 => x"0601140c",
			2049 => x"0207df04",
			2050 => x"00002059",
			2051 => x"0305a704",
			2052 => x"00002059",
			2053 => x"00602059",
			2054 => x"fe852059",
			2055 => x"06013e1c",
			2056 => x"07055f18",
			2057 => x"040df50c",
			2058 => x"0a027508",
			2059 => x"0a026904",
			2060 => x"00002059",
			2061 => x"00872059",
			2062 => x"ffa72059",
			2063 => x"06011904",
			2064 => x"00002059",
			2065 => x"02090004",
			2066 => x"01202059",
			2067 => x"00002059",
			2068 => x"00002059",
			2069 => x"ff332059",
			2070 => x"0e02d910",
			2071 => x"0f05da0c",
			2072 => x"06013a08",
			2073 => x"0303a004",
			2074 => x"019e20c5",
			2075 => x"000020c5",
			2076 => x"000020c5",
			2077 => x"ffe720c5",
			2078 => x"040d550c",
			2079 => x"06011408",
			2080 => x"06011204",
			2081 => x"feb120c5",
			2082 => x"005220c5",
			2083 => x"fe6820c5",
			2084 => x"06013e18",
			2085 => x"0e04bb14",
			2086 => x"0f05d208",
			2087 => x"00067104",
			2088 => x"016b20c5",
			2089 => x"ffda20c5",
			2090 => x"04120c04",
			2091 => x"feae20c5",
			2092 => x"0208b404",
			2093 => x"009b20c5",
			2094 => x"ffc720c5",
			2095 => x"021c20c5",
			2096 => x"fe7c20c5",
			2097 => x"0303a010",
			2098 => x"06013908",
			2099 => x"06011c04",
			2100 => x"00002141",
			2101 => x"01a02141",
			2102 => x"03039404",
			2103 => x"00002141",
			2104 => x"ff1d2141",
			2105 => x"040d550c",
			2106 => x"08028708",
			2107 => x"00032c04",
			2108 => x"fe832141",
			2109 => x"03042141",
			2110 => x"fe672141",
			2111 => x"08035b10",
			2112 => x"0208f90c",
			2113 => x"0f06d904",
			2114 => x"00002141",
			2115 => x"0504e504",
			2116 => x"00002141",
			2117 => x"02822141",
			2118 => x"ffd72141",
			2119 => x"06013a10",
			2120 => x"0803c704",
			2121 => x"feb32141",
			2122 => x"02087608",
			2123 => x"00062f04",
			2124 => x"014c2141",
			2125 => x"00002141",
			2126 => x"ff442141",
			2127 => x"fe732141",
			2128 => x"0e02f110",
			2129 => x"06013a0c",
			2130 => x"0f05b608",
			2131 => x"00080104",
			2132 => x"01c221c5",
			2133 => x"ff2321c5",
			2134 => x"fea821c5",
			2135 => x"fe8121c5",
			2136 => x"0f05e00c",
			2137 => x"0505b108",
			2138 => x"040f7004",
			2139 => x"fe9b21c5",
			2140 => x"02d621c5",
			2141 => x"fe6e21c5",
			2142 => x"040d550c",
			2143 => x"06011408",
			2144 => x"06011204",
			2145 => x"fe7d21c5",
			2146 => x"019921c5",
			2147 => x"fe6621c5",
			2148 => x"08035b0c",
			2149 => x"05064404",
			2150 => x"fec321c5",
			2151 => x"0b05c704",
			2152 => x"054721c5",
			2153 => x"ff1b21c5",
			2154 => x"06013e0c",
			2155 => x"05059204",
			2156 => x"fe6f21c5",
			2157 => x"05067904",
			2158 => x"031021c5",
			2159 => x"feaa21c5",
			2160 => x"fe6621c5",
			2161 => x"0303a014",
			2162 => x"0411de04",
			2163 => x"ffc02251",
			2164 => x"0a03880c",
			2165 => x"0c04b108",
			2166 => x"0f05d204",
			2167 => x"01a72251",
			2168 => x"00002251",
			2169 => x"02f02251",
			2170 => x"ff4d2251",
			2171 => x"040d550c",
			2172 => x"0a021008",
			2173 => x"040a6904",
			2174 => x"fe722251",
			2175 => x"10c42251",
			2176 => x"fe652251",
			2177 => x"02080910",
			2178 => x"0b04bf08",
			2179 => x"0f05b604",
			2180 => x"016b2251",
			2181 => x"fead2251",
			2182 => x"0c054604",
			2183 => x"035b2251",
			2184 => x"ff4a2251",
			2185 => x"02088314",
			2186 => x"0208740c",
			2187 => x"02081b08",
			2188 => x"0c047704",
			2189 => x"ffb42251",
			2190 => x"001b2251",
			2191 => x"fe792251",
			2192 => x"0a030804",
			2193 => x"024a2251",
			2194 => x"00002251",
			2195 => x"fe6b2251",
			2196 => x"0e02ea10",
			2197 => x"06013a0c",
			2198 => x"0f05b608",
			2199 => x"0007f604",
			2200 => x"01e722dd",
			2201 => x"fefe22dd",
			2202 => x"fe8a22dd",
			2203 => x"fe7522dd",
			2204 => x"0f05e010",
			2205 => x"0704aa0c",
			2206 => x"01002508",
			2207 => x"0f058504",
			2208 => x"01d322dd",
			2209 => x"03f122dd",
			2210 => x"fe6622dd",
			2211 => x"fe6822dd",
			2212 => x"040d550c",
			2213 => x"06011408",
			2214 => x"06011204",
			2215 => x"fe7322dd",
			2216 => x"024f22dd",
			2217 => x"fe6022dd",
			2218 => x"0207f808",
			2219 => x"06013e04",
			2220 => x"020022dd",
			2221 => x"ff6d22dd",
			2222 => x"02090010",
			2223 => x"0208f708",
			2224 => x"04120c04",
			2225 => x"fe6a22dd",
			2226 => x"ffab22dd",
			2227 => x"040f0204",
			2228 => x"065a22dd",
			2229 => x"fee522dd",
			2230 => x"fe6322dd",
			2231 => x"0303ac14",
			2232 => x"06013a10",
			2233 => x"06011904",
			2234 => x"fe56237b",
			2235 => x"00081208",
			2236 => x"0f05ad04",
			2237 => x"01fb237b",
			2238 => x"0032237b",
			2239 => x"ff00237b",
			2240 => x"fe72237b",
			2241 => x"0f05e010",
			2242 => x"0d055a0c",
			2243 => x"01002a08",
			2244 => x"0f05ad04",
			2245 => x"01e3237b",
			2246 => x"0707237b",
			2247 => x"fe93237b",
			2248 => x"fe66237b",
			2249 => x"040d550c",
			2250 => x"06011408",
			2251 => x"06011204",
			2252 => x"fe6f237b",
			2253 => x"02ea237b",
			2254 => x"fe5f237b",
			2255 => x"0207f808",
			2256 => x"06013e04",
			2257 => x"026d237b",
			2258 => x"ff5a237b",
			2259 => x"040d6e0c",
			2260 => x"0208f704",
			2261 => x"fec3237b",
			2262 => x"06016804",
			2263 => x"04a7237b",
			2264 => x"ff55237b",
			2265 => x"06013a08",
			2266 => x"06013404",
			2267 => x"fe68237b",
			2268 => x"016e237b",
			2269 => x"fe62237b",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(736, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(1502, initial_addr_3'length));
	end generate gen_rom_6;

	gen_rom_7: if SELECT_ROM = 7 generate
		bank <= (
			0 => x"040eab68",
			1 => x"09014f38",
			2 => x"0f08f928",
			3 => x"04097208",
			4 => x"07049204",
			5 => x"00000115",
			6 => x"fe0f0115",
			7 => x"09008f10",
			8 => x"0c049608",
			9 => x"09007104",
			10 => x"ffb50115",
			11 => x"00270115",
			12 => x"0e048804",
			13 => x"ffdc0115",
			14 => x"fe780115",
			15 => x"01005708",
			16 => x"0e052604",
			17 => x"01d40115",
			18 => x"ff7b0115",
			19 => x"06012104",
			20 => x"013a0115",
			21 => x"00250115",
			22 => x"05066a08",
			23 => x"09010f04",
			24 => x"02020115",
			25 => x"fe480115",
			26 => x"020bf304",
			27 => x"02530115",
			28 => x"ff2d0115",
			29 => x"0601bb1c",
			30 => x"0a029204",
			31 => x"fe640115",
			32 => x"0c05f70c",
			33 => x"020b4908",
			34 => x"06018804",
			35 => x"ffb90115",
			36 => x"fe4a0115",
			37 => x"00000115",
			38 => x"0f0b2608",
			39 => x"040d0004",
			40 => x"01290115",
			41 => x"ff3e0115",
			42 => x"fe700115",
			43 => x"0e0b770c",
			44 => x"040c2604",
			45 => x"ff140115",
			46 => x"0c061504",
			47 => x"00aa0115",
			48 => x"02020115",
			49 => x"0c06c704",
			50 => x"fe860115",
			51 => x"00d20115",
			52 => x"0601670c",
			53 => x"040fc604",
			54 => x"fdc30115",
			55 => x"04108904",
			56 => x"00000115",
			57 => x"fe6f0115",
			58 => x"02091108",
			59 => x"01001604",
			60 => x"ffcd0115",
			61 => x"01920115",
			62 => x"0a03150c",
			63 => x"0803e604",
			64 => x"febe0115",
			65 => x"04112a04",
			66 => x"01f90115",
			67 => x"00000115",
			68 => x"fe8f0115",
			69 => x"07058b3c",
			70 => x"01002a08",
			71 => x"06016b04",
			72 => x"fe610219",
			73 => x"ff950219",
			74 => x"06010a04",
			75 => x"fe600219",
			76 => x"06018520",
			77 => x"0e048810",
			78 => x"05053108",
			79 => x"03049f04",
			80 => x"00ea0219",
			81 => x"00540219",
			82 => x"06012b04",
			83 => x"01af0219",
			84 => x"00e10219",
			85 => x"0f06e308",
			86 => x"06012504",
			87 => x"010c0219",
			88 => x"ff5b0219",
			89 => x"0c04d404",
			90 => x"00630219",
			91 => x"00e30219",
			92 => x"0c05280c",
			93 => x"0a031e08",
			94 => x"0b05ca04",
			95 => x"fe3e0219",
			96 => x"ff160219",
			97 => x"010c0219",
			98 => x"017e0219",
			99 => x"08032610",
			100 => x"0100c30c",
			101 => x"0100bc04",
			102 => x"fe7a0219",
			103 => x"0506c504",
			104 => x"fee90219",
			105 => x"02a90219",
			106 => x"fe5d0219",
			107 => x"0803fa2c",
			108 => x"0e0a2a14",
			109 => x"0901db10",
			110 => x"0f091508",
			111 => x"0d06c504",
			112 => x"01740219",
			113 => x"fe4c0219",
			114 => x"06018a04",
			115 => x"03230219",
			116 => x"00ee0219",
			117 => x"fe580219",
			118 => x"0601b708",
			119 => x"08032804",
			120 => x"00860219",
			121 => x"fe4c0219",
			122 => x"0c06a108",
			123 => x"0a02d104",
			124 => x"fe390219",
			125 => x"00130219",
			126 => x"0f0be504",
			127 => x"03700219",
			128 => x"ffea0219",
			129 => x"08045308",
			130 => x"08044e04",
			131 => x"fe6b0219",
			132 => x"01400219",
			133 => x"fe5f0219",
			134 => x"0c057f60",
			135 => x"01003210",
			136 => x"02076708",
			137 => x"06012d04",
			138 => x"fecb033d",
			139 => x"01e3033d",
			140 => x"06016f04",
			141 => x"fe61033d",
			142 => x"0000033d",
			143 => x"0409b310",
			144 => x"0e04f004",
			145 => x"ff82033d",
			146 => x"0b056904",
			147 => x"fe17033d",
			148 => x"0b057404",
			149 => x"0000033d",
			150 => x"fe6d033d",
			151 => x"0c04b220",
			152 => x"0c049610",
			153 => x"0c049408",
			154 => x"03049704",
			155 => x"00be033d",
			156 => x"0029033d",
			157 => x"040d6e04",
			158 => x"00ed033d",
			159 => x"fe0e033d",
			160 => x"040c7208",
			161 => x"0c049704",
			162 => x"ff24033d",
			163 => x"fffa033d",
			164 => x"0c049904",
			165 => x"0000033d",
			166 => x"014b033d",
			167 => x"0c04b410",
			168 => x"0a029008",
			169 => x"0208c704",
			170 => x"0171033d",
			171 => x"03a6033d",
			172 => x"040bb204",
			173 => x"feb1033d",
			174 => x"00f3033d",
			175 => x"0c04b508",
			176 => x"0f072504",
			177 => x"005c033d",
			178 => x"fdcd033d",
			179 => x"0e050704",
			180 => x"0104033d",
			181 => x"004c033d",
			182 => x"08032608",
			183 => x"0e06ac04",
			184 => x"0157033d",
			185 => x"fe6a033d",
			186 => x"040eab28",
			187 => x"08034c10",
			188 => x"020b1c0c",
			189 => x"040c0408",
			190 => x"040bb004",
			191 => x"ff97033d",
			192 => x"039f033d",
			193 => x"fe8a033d",
			194 => x"fe67033d",
			195 => x"040ce10c",
			196 => x"040bf104",
			197 => x"ffbc033d",
			198 => x"0c05d404",
			199 => x"00db033d",
			200 => x"0253033d",
			201 => x"08037304",
			202 => x"fe29033d",
			203 => x"06019e04",
			204 => x"fe4a033d",
			205 => x"011f033d",
			206 => x"fe64033d",
			207 => x"07057764",
			208 => x"040e2348",
			209 => x"06010a08",
			210 => x"06010604",
			211 => x"fe500481",
			212 => x"ffac0481",
			213 => x"0e04e220",
			214 => x"0b04c010",
			215 => x"0304d808",
			216 => x"07047804",
			217 => x"008a0481",
			218 => x"01ab0481",
			219 => x"0f070504",
			220 => x"00b30481",
			221 => x"01960481",
			222 => x"040bec08",
			223 => x"06014104",
			224 => x"01be0481",
			225 => x"003c0481",
			226 => x"09009904",
			227 => x"01c10481",
			228 => x"025d0481",
			229 => x"040bb210",
			230 => x"0704ec08",
			231 => x"06014a04",
			232 => x"00490481",
			233 => x"fef40481",
			234 => x"09013104",
			235 => x"012f0481",
			236 => x"fea40481",
			237 => x"06017008",
			238 => x"0900b304",
			239 => x"00e60481",
			240 => x"01b50481",
			241 => x"07051f04",
			242 => x"ff2b0481",
			243 => x"01530481",
			244 => x"06014108",
			245 => x"0d054d04",
			246 => x"fe480481",
			247 => x"ff5c0481",
			248 => x"0505a00c",
			249 => x"06014a04",
			250 => x"ff670481",
			251 => x"00057a04",
			252 => x"00d20481",
			253 => x"02710481",
			254 => x"0f08d404",
			255 => x"fe3a0481",
			256 => x"01a90481",
			257 => x"0803260c",
			258 => x"0705a908",
			259 => x"0705a504",
			260 => x"fe590481",
			261 => x"02040481",
			262 => x"fe470481",
			263 => x"040e6330",
			264 => x"08035218",
			265 => x"0f0ad90c",
			266 => x"040c6008",
			267 => x"040ba404",
			268 => x"ff9e0481",
			269 => x"046e0481",
			270 => x"fe580481",
			271 => x"08032804",
			272 => x"00000481",
			273 => x"07073804",
			274 => x"fe460481",
			275 => x"ffea0481",
			276 => x"0f0c3910",
			277 => x"040c1208",
			278 => x"0a02c704",
			279 => x"00680481",
			280 => x"fe3f0481",
			281 => x"00043904",
			282 => x"050c0481",
			283 => x"019e0481",
			284 => x"0601d004",
			285 => x"fe150481",
			286 => x"01b60481",
			287 => x"fe4b0481",
			288 => x"07056164",
			289 => x"040eab44",
			290 => x"06010a04",
			291 => x"fe6305cd",
			292 => x"040c5e20",
			293 => x"0a02ac10",
			294 => x"0208ce08",
			295 => x"06014104",
			296 => x"008f05cd",
			297 => x"001e05cd",
			298 => x"06015204",
			299 => x"01fc05cd",
			300 => x"009105cd",
			301 => x"0208b908",
			302 => x"0900b304",
			303 => x"fff805cd",
			304 => x"019005cd",
			305 => x"0c04d404",
			306 => x"ff0505cd",
			307 => x"009605cd",
			308 => x"09008010",
			309 => x"0304ef08",
			310 => x"03043704",
			311 => x"016305cd",
			312 => x"005805cd",
			313 => x"0b049004",
			314 => x"010805cd",
			315 => x"fea505cd",
			316 => x"0505bf08",
			317 => x"03050004",
			318 => x"016d05cd",
			319 => x"00db05cd",
			320 => x"0f08c604",
			321 => x"ff9105cd",
			322 => x"01d805cd",
			323 => x"01005618",
			324 => x"09005514",
			325 => x"01002504",
			326 => x"fe6105cd",
			327 => x"0504e708",
			328 => x"04108904",
			329 => x"fe1405cd",
			330 => x"000005cd",
			331 => x"02087404",
			332 => x"014205cd",
			333 => x"fee805cd",
			334 => x"fd7a05cd",
			335 => x"040f0204",
			336 => x"006305cd",
			337 => x"fe7005cd",
			338 => x"08032610",
			339 => x"0100c30c",
			340 => x"0100bc04",
			341 => x"fe3905cd",
			342 => x"0b05f904",
			343 => x"fef105cd",
			344 => x"027b05cd",
			345 => x"fe5f05cd",
			346 => x"040e6324",
			347 => x"0a02e81c",
			348 => x"06018a0c",
			349 => x"06018308",
			350 => x"0100ad04",
			351 => x"01b905cd",
			352 => x"fe9d05cd",
			353 => x"02ec05cd",
			354 => x"07068808",
			355 => x"08032b04",
			356 => x"003505cd",
			357 => x"fe8005cd",
			358 => x"040c4704",
			359 => x"01fc05cd",
			360 => x"ff6705cd",
			361 => x"0a02fd04",
			362 => x"00f005cd",
			363 => x"021405cd",
			364 => x"0411030c",
			365 => x"08044e04",
			366 => x"feaf05cd",
			367 => x"0a037204",
			368 => x"018205cd",
			369 => x"fed305cd",
			370 => x"fe6005cd",
			371 => x"0705617c",
			372 => x"01003210",
			373 => x"02076708",
			374 => x"04117604",
			375 => x"01750759",
			376 => x"febe0759",
			377 => x"0a038504",
			378 => x"fe5f0759",
			379 => x"00000759",
			380 => x"0704913c",
			381 => x"0304af20",
			382 => x"0504e710",
			383 => x"03045e08",
			384 => x"0004b804",
			385 => x"fff80759",
			386 => x"01760759",
			387 => x"0504e404",
			388 => x"ff750759",
			389 => x"fd4b0759",
			390 => x"0a02d408",
			391 => x"09006204",
			392 => x"00000759",
			393 => x"015c0759",
			394 => x"0e03a604",
			395 => x"00690759",
			396 => x"fd910759",
			397 => x"0900770c",
			398 => x"0c048f08",
			399 => x"0e040e04",
			400 => x"000a0759",
			401 => x"fdc30759",
			402 => x"011d0759",
			403 => x"0304f708",
			404 => x"0b048004",
			405 => x"fe820759",
			406 => x"00880759",
			407 => x"02089004",
			408 => x"fee10759",
			409 => x"003c0759",
			410 => x"0409b310",
			411 => x"0e04f004",
			412 => x"fffe0759",
			413 => x"07052f04",
			414 => x"fe060759",
			415 => x"07053104",
			416 => x"00470759",
			417 => x"fe7a0759",
			418 => x"0a024710",
			419 => x"0d054108",
			420 => x"0e046104",
			421 => x"009b0759",
			422 => x"fcc70759",
			423 => x"040a0104",
			424 => x"006f0759",
			425 => x"01d80759",
			426 => x"0e04f708",
			427 => x"09009c04",
			428 => x"00780759",
			429 => x"012f0759",
			430 => x"02086204",
			431 => x"ffba0759",
			432 => x"00680759",
			433 => x"0a029218",
			434 => x"0e068d0c",
			435 => x"0d06d408",
			436 => x"0e060f04",
			437 => x"00000759",
			438 => x"fe530759",
			439 => x"02100759",
			440 => x"09013108",
			441 => x"09012704",
			442 => x"fe0e0759",
			443 => x"00d70759",
			444 => x"fe650759",
			445 => x"040f0228",
			446 => x"0a02e81c",
			447 => x"020a460c",
			448 => x"040d5508",
			449 => x"0f091f04",
			450 => x"00a80759",
			451 => x"02d80759",
			452 => x"fe400759",
			453 => x"07068808",
			454 => x"0901a104",
			455 => x"ffc00759",
			456 => x"fe490759",
			457 => x"0f0bae04",
			458 => x"01420759",
			459 => x"ff320759",
			460 => x"0a030808",
			461 => x"0f0c3904",
			462 => x"01b10759",
			463 => x"fe990759",
			464 => x"03040759",
			465 => x"04110308",
			466 => x"0410e104",
			467 => x"fe720759",
			468 => x"00000759",
			469 => x"fe620759",
			470 => x"040df598",
			471 => x"0505f93c",
			472 => x"07051b28",
			473 => x"01009520",
			474 => x"0f06e310",
			475 => x"0e043608",
			476 => x"0b049104",
			477 => x"ffe80905",
			478 => x"007d0905",
			479 => x"0a029e04",
			480 => x"ffe60905",
			481 => x"ff310905",
			482 => x"06014108",
			483 => x"0505a104",
			484 => x"00440905",
			485 => x"01610905",
			486 => x"0c045b04",
			487 => x"01640905",
			488 => x"00030905",
			489 => x"040ae204",
			490 => x"02f40905",
			491 => x"000e0905",
			492 => x"0f080e0c",
			493 => x"06015108",
			494 => x"0e057804",
			495 => x"01630905",
			496 => x"feb20905",
			497 => x"01fe0905",
			498 => x"0c04ed04",
			499 => x"fee40905",
			500 => x"01a80905",
			501 => x"0a028d2c",
			502 => x"0208521c",
			503 => x"0208240c",
			504 => x"0f071708",
			505 => x"0f06ed04",
			506 => x"feef0905",
			507 => x"00e60905",
			508 => x"fe5f0905",
			509 => x"02083708",
			510 => x"06012504",
			511 => x"00000905",
			512 => x"02970905",
			513 => x"02084d04",
			514 => x"fec30905",
			515 => x"021f0905",
			516 => x"05060804",
			517 => x"fdbc0905",
			518 => x"05061504",
			519 => x"01940905",
			520 => x"08032e04",
			521 => x"fef00905",
			522 => x"fcab0905",
			523 => x"0c04ec14",
			524 => x"0e065a04",
			525 => x"fdf30905",
			526 => x"06017908",
			527 => x"0100a104",
			528 => x"01040905",
			529 => x"fe9a0905",
			530 => x"0f091504",
			531 => x"fe5a0905",
			532 => x"002f0905",
			533 => x"00040810",
			534 => x"0f0b2608",
			535 => x"040bb004",
			536 => x"00d90905",
			537 => x"02900905",
			538 => x"0a02b404",
			539 => x"fea40905",
			540 => x"01510905",
			541 => x"0c04ed04",
			542 => x"01a90905",
			543 => x"0c052e04",
			544 => x"ff7b0905",
			545 => x"008e0905",
			546 => x"0803d020",
			547 => x"0100470c",
			548 => x"040eab08",
			549 => x"01002d04",
			550 => x"ff920905",
			551 => x"01750905",
			552 => x"feb10905",
			553 => x"0c04b304",
			554 => x"fc550905",
			555 => x"0004c104",
			556 => x"fe5d0905",
			557 => x"06016804",
			558 => x"00bf0905",
			559 => x"0100c504",
			560 => x"ff160905",
			561 => x"00000905",
			562 => x"04112a18",
			563 => x"00051508",
			564 => x"0100c204",
			565 => x"fdc90905",
			566 => x"00710905",
			567 => x"0d04f304",
			568 => x"ff010905",
			569 => x"0b04b004",
			570 => x"01a30905",
			571 => x"0704ef04",
			572 => x"fefc0905",
			573 => x"00f00905",
			574 => x"0c043a04",
			575 => x"00000905",
			576 => x"fe8d0905",
			577 => x"040eab9c",
			578 => x"09014f68",
			579 => x"02083338",
			580 => x"0e04f018",
			581 => x"0d058d0c",
			582 => x"0704db08",
			583 => x"06012504",
			584 => x"006d0a99",
			585 => x"fff40a99",
			586 => x"fd750a99",
			587 => x"01007108",
			588 => x"02081d04",
			589 => x"01ba0a99",
			590 => x"ffb80a99",
			591 => x"fee70a99",
			592 => x"0900a810",
			593 => x"03054f08",
			594 => x"09009504",
			595 => x"fe270a99",
			596 => x"01560a99",
			597 => x"05053d04",
			598 => x"00db0a99",
			599 => x"fe3c0a99",
			600 => x"05057408",
			601 => x"0e053404",
			602 => x"02c60a99",
			603 => x"00000a99",
			604 => x"0003f704",
			605 => x"00000a99",
			606 => x"fe610a99",
			607 => x"02083710",
			608 => x"06012d04",
			609 => x"006f0a99",
			610 => x"00040b04",
			611 => x"043e0a99",
			612 => x"0704c304",
			613 => x"025b0a99",
			614 => x"fffe0a99",
			615 => x"0803a310",
			616 => x"01004108",
			617 => x"0504f404",
			618 => x"fd4b0a99",
			619 => x"ff330a99",
			620 => x"08034204",
			621 => x"006b0a99",
			622 => x"001b0a99",
			623 => x"0f06ca08",
			624 => x"0b049d04",
			625 => x"01aa0a99",
			626 => x"fe7b0a99",
			627 => x"06017004",
			628 => x"01a00a99",
			629 => x"00240a99",
			630 => x"0601bb20",
			631 => x"08032604",
			632 => x"fe640a99",
			633 => x"0706440c",
			634 => x"020b3208",
			635 => x"06018804",
			636 => x"ff600a99",
			637 => x"fe3c0a99",
			638 => x"00170a99",
			639 => x"020b3908",
			640 => x"0901d004",
			641 => x"01810a99",
			642 => x"00000a99",
			643 => x"0901c604",
			644 => x"ff980a99",
			645 => x"fe600a99",
			646 => x"0e0b770c",
			647 => x"040c2604",
			648 => x"ff050a99",
			649 => x"07068804",
			650 => x"00c00a99",
			651 => x"02250a99",
			652 => x"07075004",
			653 => x"fe880a99",
			654 => x"00e30a99",
			655 => x"06016714",
			656 => x"040fc604",
			657 => x"fdad0a99",
			658 => x"04100808",
			659 => x"09004204",
			660 => x"00000a99",
			661 => x"00450a99",
			662 => x"01003204",
			663 => x"fe6a0a99",
			664 => x"ffb50a99",
			665 => x"02091108",
			666 => x"01001604",
			667 => x"ffb30a99",
			668 => x"01a80a99",
			669 => x"0803f110",
			670 => x"0803e604",
			671 => x"feab0a99",
			672 => x"020a8604",
			673 => x"ffdb0a99",
			674 => x"0100c304",
			675 => x"020c0a99",
			676 => x"00000a99",
			677 => x"fe860a99",
			678 => x"040a0118",
			679 => x"06013114",
			680 => x"0900a908",
			681 => x"05055704",
			682 => x"fda70c05",
			683 => x"ff340c05",
			684 => x"00033e04",
			685 => x"fe750c05",
			686 => x"0704d604",
			687 => x"00630c05",
			688 => x"018b0c05",
			689 => x"fe3b0c05",
			690 => x"040d5558",
			691 => x"0004b834",
			692 => x"0504e714",
			693 => x"0504e510",
			694 => x"02081108",
			695 => x"06013104",
			696 => x"ff950c05",
			697 => x"01860c05",
			698 => x"03048f04",
			699 => x"fefe0c05",
			700 => x"fd2f0c05",
			701 => x"fcf10c05",
			702 => x"0b048010",
			703 => x"040c3808",
			704 => x"0304cf04",
			705 => x"018d0c05",
			706 => x"ffed0c05",
			707 => x"07047e04",
			708 => x"ff280c05",
			709 => x"01520c05",
			710 => x"0b048108",
			711 => x"0c047804",
			712 => x"fcbe0c05",
			713 => x"00990c05",
			714 => x"09008f04",
			715 => x"ffe90c05",
			716 => x"001e0c05",
			717 => x"0e04b418",
			718 => x"0b047d0c",
			719 => x"0504e708",
			720 => x"0504e204",
			721 => x"01c40c05",
			722 => x"00a00c05",
			723 => x"feec0c05",
			724 => x"0a02ed08",
			725 => x"0704a904",
			726 => x"01d50c05",
			727 => x"010e0c05",
			728 => x"00090c05",
			729 => x"0e04d304",
			730 => x"fd510c05",
			731 => x"01006d04",
			732 => x"01b10c05",
			733 => x"ff920c05",
			734 => x"0f075524",
			735 => x"0e04a520",
			736 => x"07047b10",
			737 => x"0a031b08",
			738 => x"0b047104",
			739 => x"fe7f0c05",
			740 => x"fcf10c05",
			741 => x"0504d704",
			742 => x"ff0e0c05",
			743 => x"00000c05",
			744 => x"0c047708",
			745 => x"040eab04",
			746 => x"01870c05",
			747 => x"ff230c05",
			748 => x"02089804",
			749 => x"fed60c05",
			750 => x"00c70c05",
			751 => x"fcae0c05",
			752 => x"07057314",
			753 => x"02091908",
			754 => x"03056f04",
			755 => x"01d20c05",
			756 => x"fe080c05",
			757 => x"0004b804",
			758 => x"ff6e0c05",
			759 => x"040f0204",
			760 => x"01ce0c05",
			761 => x"ff850c05",
			762 => x"00048e04",
			763 => x"fe6d0c05",
			764 => x"0100e508",
			765 => x"0307c404",
			766 => x"006a0c05",
			767 => x"febe0c05",
			768 => x"012f0c05",
			769 => x"0803a370",
			770 => x"0207a12c",
			771 => x"06013e28",
			772 => x"0a026714",
			773 => x"0207920c",
			774 => x"06012b08",
			775 => x"040ab204",
			776 => x"ffad0d89",
			777 => x"00f00d89",
			778 => x"ff0c0d89",
			779 => x"06012104",
			780 => x"ff5d0d89",
			781 => x"fdd00d89",
			782 => x"0d054110",
			783 => x"06012d08",
			784 => x"0d050d04",
			785 => x"00000d89",
			786 => x"01930d89",
			787 => x"06013504",
			788 => x"fecb0d89",
			789 => x"001f0d89",
			790 => x"01fa0d89",
			791 => x"fe0d0d89",
			792 => x"0207a708",
			793 => x"0f066604",
			794 => x"01a40d89",
			795 => x"00610d89",
			796 => x"040b701c",
			797 => x"0304ef0c",
			798 => x"0f06ac08",
			799 => x"0e044b04",
			800 => x"01150d89",
			801 => x"ff6a0d89",
			802 => x"01f40d89",
			803 => x"0d053508",
			804 => x"06012504",
			805 => x"fe150d89",
			806 => x"ff7e0d89",
			807 => x"03054304",
			808 => x"009a0d89",
			809 => x"000a0d89",
			810 => x"040b8010",
			811 => x"09009908",
			812 => x"06012504",
			813 => x"01740d89",
			814 => x"fe800d89",
			815 => x"0d057504",
			816 => x"01050d89",
			817 => x"ff6f0d89",
			818 => x"040b8308",
			819 => x"0c050c04",
			820 => x"01c20d89",
			821 => x"fe360d89",
			822 => x"0505b104",
			823 => x"00050d89",
			824 => x"ffb40d89",
			825 => x"0a02db10",
			826 => x"06015b08",
			827 => x"01003204",
			828 => x"00000d89",
			829 => x"01910d89",
			830 => x"0208bb04",
			831 => x"ff0a0d89",
			832 => x"00fd0d89",
			833 => x"0c045608",
			834 => x"0a033104",
			835 => x"fdd50d89",
			836 => x"00000d89",
			837 => x"06015120",
			838 => x"07049710",
			839 => x"07047b08",
			840 => x"0e02bd04",
			841 => x"00c90d89",
			842 => x"fe620d89",
			843 => x"01003904",
			844 => x"00000d89",
			845 => x"01a30d89",
			846 => x"02086c08",
			847 => x"08040204",
			848 => x"fe0a0d89",
			849 => x"00000d89",
			850 => x"0c054604",
			851 => x"00320d89",
			852 => x"00000d89",
			853 => x"040d000c",
			854 => x"040ce108",
			855 => x"06016b04",
			856 => x"014e0d89",
			857 => x"ff6c0d89",
			858 => x"fe1b0d89",
			859 => x"040eab08",
			860 => x"0803ac04",
			861 => x"00000d89",
			862 => x"01350d89",
			863 => x"08042b04",
			864 => x"ff520d89",
			865 => x"008a0d89",
			866 => x"07057798",
			867 => x"01003920",
			868 => x"01002504",
			869 => x"fe5b0f3d",
			870 => x"0304350c",
			871 => x"0b046d04",
			872 => x"fef50f3d",
			873 => x"0207da04",
			874 => x"02390f3d",
			875 => x"00000f3d",
			876 => x"0a02bc0c",
			877 => x"08038a08",
			878 => x"0207ca04",
			879 => x"ffb70f3d",
			880 => x"fe260f3d",
			881 => x"00000f3d",
			882 => x"fd560f3d",
			883 => x"0e058740",
			884 => x"0704c120",
			885 => x"03050010",
			886 => x"07047808",
			887 => x"02080704",
			888 => x"00880f3d",
			889 => x"fec00f3d",
			890 => x"03047704",
			891 => x"01790f3d",
			892 => x"00d60f3d",
			893 => x"02085408",
			894 => x"0e04bb04",
			895 => x"00420f3d",
			896 => x"ff840f3d",
			897 => x"0c047204",
			898 => x"ff440f3d",
			899 => x"00c00f3d",
			900 => x"0704c410",
			901 => x"0a02b408",
			902 => x"0d058204",
			903 => x"01aa0f3d",
			904 => x"02b70f3d",
			905 => x"040c6c04",
			906 => x"ffc20f3d",
			907 => x"01700f3d",
			908 => x"0704d508",
			909 => x"0505a004",
			910 => x"000b0f3d",
			911 => x"01c90f3d",
			912 => x"0e04f004",
			913 => x"016e0f3d",
			914 => x"00cc0f3d",
			915 => x"0208981c",
			916 => x"06015610",
			917 => x"0a026d08",
			918 => x"040adc04",
			919 => x"ff3b0f3d",
			920 => x"02e40f3d",
			921 => x"0c04ce04",
			922 => x"fe160f3d",
			923 => x"00000f3d",
			924 => x"02085404",
			925 => x"03250f3d",
			926 => x"0b052204",
			927 => x"ff000f3d",
			928 => x"00f40f3d",
			929 => x"06014a0c",
			930 => x"01006504",
			931 => x"fdf60f3d",
			932 => x"0b053504",
			933 => x"03540f3d",
			934 => x"00110f3d",
			935 => x"0c04f108",
			936 => x"06017704",
			937 => x"00370f3d",
			938 => x"fefe0f3d",
			939 => x"0100c204",
			940 => x"01470f3d",
			941 => x"fe650f3d",
			942 => x"0803260c",
			943 => x"0100c308",
			944 => x"0100bd04",
			945 => x"fe780f3d",
			946 => x"02360f3d",
			947 => x"fe5c0f3d",
			948 => x"040e6328",
			949 => x"08037318",
			950 => x"0e0ab80c",
			951 => x"040d0008",
			952 => x"040b8304",
			953 => x"ff0d0f3d",
			954 => x"01cc0f3d",
			955 => x"fe250f3d",
			956 => x"0601be04",
			957 => x"fe540f3d",
			958 => x"0601c004",
			959 => x"00a30f3d",
			960 => x"fe5c0f3d",
			961 => x"040d8808",
			962 => x"07068804",
			963 => x"01110f3d",
			964 => x"02690f3d",
			965 => x"08039c04",
			966 => x"fe170f3d",
			967 => x"01d10f3d",
			968 => x"0411030c",
			969 => x"08044e04",
			970 => x"fe930f3d",
			971 => x"0a037204",
			972 => x"01980f3d",
			973 => x"fea30f3d",
			974 => x"fe5b0f3d",
			975 => x"0d06119c",
			976 => x"07047840",
			977 => x"07046728",
			978 => x"0c045910",
			979 => x"0b047d0c",
			980 => x"040d0008",
			981 => x"00042104",
			982 => x"fe121119",
			983 => x"01ee1119",
			984 => x"fe651119",
			985 => x"fd651119",
			986 => x"040c7f08",
			987 => x"02081504",
			988 => x"01d21119",
			989 => x"ff101119",
			990 => x"0a02c308",
			991 => x"0504f204",
			992 => x"00b91119",
			993 => x"fd0b1119",
			994 => x"0303f504",
			995 => x"feb41119",
			996 => x"01ae1119",
			997 => x"0a02a910",
			998 => x"06011008",
			999 => x"0f069904",
			1000 => x"01801119",
			1001 => x"ff8c1119",
			1002 => x"01004d04",
			1003 => x"fc781119",
			1004 => x"fe9e1119",
			1005 => x"0803a704",
			1006 => x"01311119",
			1007 => x"fe731119",
			1008 => x"0a027838",
			1009 => x"0208091c",
			1010 => x"0505110c",
			1011 => x"0304ef08",
			1012 => x"07049104",
			1013 => x"fe1f1119",
			1014 => x"00691119",
			1015 => x"fc2a1119",
			1016 => x"03051b08",
			1017 => x"05053104",
			1018 => x"00421119",
			1019 => x"01541119",
			1020 => x"0802fb04",
			1021 => x"005c1119",
			1022 => x"ff3a1119",
			1023 => x"040b3610",
			1024 => x"0a026508",
			1025 => x"040abb04",
			1026 => x"000a1119",
			1027 => x"01b31119",
			1028 => x"040a8804",
			1029 => x"03131119",
			1030 => x"ff5f1119",
			1031 => x"0802fb04",
			1032 => x"fde41119",
			1033 => x"0f06d904",
			1034 => x"001a1119",
			1035 => x"016d1119",
			1036 => x"0003ed04",
			1037 => x"03101119",
			1038 => x"040b8010",
			1039 => x"07049708",
			1040 => x"02083d04",
			1041 => x"002f1119",
			1042 => x"03021119",
			1043 => x"0505df04",
			1044 => x"ff661119",
			1045 => x"01e41119",
			1046 => x"0704be08",
			1047 => x"0704bc04",
			1048 => x"00241119",
			1049 => x"ff481119",
			1050 => x"0704c204",
			1051 => x"00d61119",
			1052 => x"00301119",
			1053 => x"0003a618",
			1054 => x"05061610",
			1055 => x"07051a08",
			1056 => x"0d062b04",
			1057 => x"ff491119",
			1058 => x"00ad1119",
			1059 => x"0001f104",
			1060 => x"ff791119",
			1061 => x"021a1119",
			1062 => x"0802f804",
			1063 => x"fe631119",
			1064 => x"002c1119",
			1065 => x"04110338",
			1066 => x"0b05521c",
			1067 => x"0306a50c",
			1068 => x"01008204",
			1069 => x"fedb1119",
			1070 => x"0f07f204",
			1071 => x"00451119",
			1072 => x"01771119",
			1073 => x"0a029908",
			1074 => x"0f082b04",
			1075 => x"fe2a1119",
			1076 => x"01a21119",
			1077 => x"06017004",
			1078 => x"fcfd1119",
			1079 => x"fe3e1119",
			1080 => x"0306a50c",
			1081 => x"05062608",
			1082 => x"03069604",
			1083 => x"00291119",
			1084 => x"fded1119",
			1085 => x"fd3a1119",
			1086 => x"06018a08",
			1087 => x"07051a04",
			1088 => x"ff621119",
			1089 => x"00ce1119",
			1090 => x"08032604",
			1091 => x"fe701119",
			1092 => x"ffd11119",
			1093 => x"fe6a1119",
			1094 => x"040f02bc",
			1095 => x"0304a750",
			1096 => x"06012b24",
			1097 => x"0207aa10",
			1098 => x"0b047104",
			1099 => x"fd9f12bd",
			1100 => x"040ac904",
			1101 => x"ff6d12bd",
			1102 => x"0c047204",
			1103 => x"004112bd",
			1104 => x"01bd12bd",
			1105 => x"08034f0c",
			1106 => x"0b048008",
			1107 => x"03049704",
			1108 => x"003c12bd",
			1109 => x"fc4a12bd",
			1110 => x"fc8012bd",
			1111 => x"0c044304",
			1112 => x"000012bd",
			1113 => x"01a812bd",
			1114 => x"040c4c18",
			1115 => x"0f065f10",
			1116 => x"06013508",
			1117 => x"0207b704",
			1118 => x"01e312bd",
			1119 => x"008712bd",
			1120 => x"0e03cb04",
			1121 => x"013312bd",
			1122 => x"ff3f12bd",
			1123 => x"08034204",
			1124 => x"00d712bd",
			1125 => x"01f512bd",
			1126 => x"00048208",
			1127 => x"0e03e704",
			1128 => x"000012bd",
			1129 => x"fc3b12bd",
			1130 => x"0f06c508",
			1131 => x"02084b04",
			1132 => x"007c12bd",
			1133 => x"fe5f12bd",
			1134 => x"021512bd",
			1135 => x"0505102c",
			1136 => x"0e03f90c",
			1137 => x"05050208",
			1138 => x"0304b704",
			1139 => x"00cd12bd",
			1140 => x"fdf312bd",
			1141 => x"fa6512bd",
			1142 => x"01004d10",
			1143 => x"01004508",
			1144 => x"0004a704",
			1145 => x"fe7b12bd",
			1146 => x"008f12bd",
			1147 => x"06014604",
			1148 => x"00af12bd",
			1149 => x"fdb212bd",
			1150 => x"0b049108",
			1151 => x"07048004",
			1152 => x"000012bd",
			1153 => x"fc2a12bd",
			1154 => x"0304f704",
			1155 => x"012412bd",
			1156 => x"feda12bd",
			1157 => x"0b049d20",
			1158 => x"0b048e10",
			1159 => x"040bf108",
			1160 => x"06012804",
			1161 => x"010312bd",
			1162 => x"fdd112bd",
			1163 => x"0b048004",
			1164 => x"01e912bd",
			1165 => x"007812bd",
			1166 => x"0c047208",
			1167 => x"0a028d04",
			1168 => x"01e412bd",
			1169 => x"fe1412bd",
			1170 => x"0f071f04",
			1171 => x"00fc12bd",
			1172 => x"025612bd",
			1173 => x"07049010",
			1174 => x"0f074908",
			1175 => x"05051e04",
			1176 => x"009e12bd",
			1177 => x"fe9512bd",
			1178 => x"02089f04",
			1179 => x"036a12bd",
			1180 => x"ff9912bd",
			1181 => x"0304be08",
			1182 => x"0f066604",
			1183 => x"fd3812bd",
			1184 => x"fff712bd",
			1185 => x"0304d804",
			1186 => x"010a12bd",
			1187 => x"001512bd",
			1188 => x"0704bc14",
			1189 => x"0c04780c",
			1190 => x"05050004",
			1191 => x"fe9712bd",
			1192 => x"05050e04",
			1193 => x"00a312bd",
			1194 => x"fe4812bd",
			1195 => x"02082204",
			1196 => x"ff8a12bd",
			1197 => x"013b12bd",
			1198 => x"fe6912bd",
			1199 => x"0c04d190",
			1200 => x"07050464",
			1201 => x"0505b030",
			1202 => x"0c04d014",
			1203 => x"0900d310",
			1204 => x"09008f08",
			1205 => x"03050d04",
			1206 => x"000914d1",
			1207 => x"ff9514d1",
			1208 => x"01005504",
			1209 => x"01a514d1",
			1210 => x"001414d1",
			1211 => x"01e314d1",
			1212 => x"0b04f110",
			1213 => x"0a02a808",
			1214 => x"08033a04",
			1215 => x"ff9c14d1",
			1216 => x"01f714d1",
			1217 => x"040c6004",
			1218 => x"fdbf14d1",
			1219 => x"016314d1",
			1220 => x"08038208",
			1221 => x"0a027f04",
			1222 => x"000914d1",
			1223 => x"023a14d1",
			1224 => x"fffc14d1",
			1225 => x"0900d620",
			1226 => x"0b052010",
			1227 => x"0c04ca08",
			1228 => x"0704da04",
			1229 => x"fe5914d1",
			1230 => x"000014d1",
			1231 => x"0704ed04",
			1232 => x"024714d1",
			1233 => x"fee914d1",
			1234 => x"0f078e08",
			1235 => x"0900c404",
			1236 => x"fee914d1",
			1237 => x"010d14d1",
			1238 => x"0b052404",
			1239 => x"fdb514d1",
			1240 => x"ff4914d1",
			1241 => x"0c04af04",
			1242 => x"025014d1",
			1243 => x"0e061e08",
			1244 => x"0208c004",
			1245 => x"ffee14d1",
			1246 => x"022e14d1",
			1247 => x"02090004",
			1248 => x"fe8114d1",
			1249 => x"00d714d1",
			1250 => x"08037c24",
			1251 => x"0505db0c",
			1252 => x"02085204",
			1253 => x"ff5814d1",
			1254 => x"08036f04",
			1255 => x"023714d1",
			1256 => x"010314d1",
			1257 => x"0d06450c",
			1258 => x"0a02a308",
			1259 => x"0b055404",
			1260 => x"010e14d1",
			1261 => x"fe2114d1",
			1262 => x"fe9514d1",
			1263 => x"09010f08",
			1264 => x"02091904",
			1265 => x"00da14d1",
			1266 => x"022b14d1",
			1267 => x"ffb114d1",
			1268 => x"08038d04",
			1269 => x"fda614d1",
			1270 => x"00ae14d1",
			1271 => x"0c04d220",
			1272 => x"0505df18",
			1273 => x"0d05ab08",
			1274 => x"0f078e04",
			1275 => x"fed714d1",
			1276 => x"00dd14d1",
			1277 => x"0a02b90c",
			1278 => x"01008008",
			1279 => x"02085b04",
			1280 => x"ff1c14d1",
			1281 => x"fd8f14d1",
			1282 => x"ff9714d1",
			1283 => x"ffb914d1",
			1284 => x"0e067104",
			1285 => x"01ef14d1",
			1286 => x"feec14d1",
			1287 => x"0c04ea24",
			1288 => x"0c04e914",
			1289 => x"0705080c",
			1290 => x"0f070904",
			1291 => x"025514d1",
			1292 => x"02087e04",
			1293 => x"fee614d1",
			1294 => x"00ac14d1",
			1295 => x"08036c04",
			1296 => x"fdb014d1",
			1297 => x"009514d1",
			1298 => x"08033a08",
			1299 => x"0a028304",
			1300 => x"01fb14d1",
			1301 => x"fd9314d1",
			1302 => x"02093504",
			1303 => x"022f14d1",
			1304 => x"000014d1",
			1305 => x"01006c18",
			1306 => x"0f07010c",
			1307 => x"0f06e508",
			1308 => x"0f06de04",
			1309 => x"ff5a14d1",
			1310 => x"002914d1",
			1311 => x"fe2a14d1",
			1312 => x"0505ea08",
			1313 => x"0704ef04",
			1314 => x"011a14d1",
			1315 => x"026114d1",
			1316 => x"000014d1",
			1317 => x"01008010",
			1318 => x"0c04f108",
			1319 => x"01007804",
			1320 => x"ff9714d1",
			1321 => x"fe5814d1",
			1322 => x"0e05ac04",
			1323 => x"ff9614d1",
			1324 => x"019114d1",
			1325 => x"0a029308",
			1326 => x"0e06ce04",
			1327 => x"fed914d1",
			1328 => x"000014d1",
			1329 => x"0d061f04",
			1330 => x"013d14d1",
			1331 => x"ffd314d1",
			1332 => x"0004b8b0",
			1333 => x"0a02be54",
			1334 => x"0207a128",
			1335 => x"02076714",
			1336 => x"0003c40c",
			1337 => x"0b049e04",
			1338 => x"fe1216f5",
			1339 => x"0c049804",
			1340 => x"00f916f5",
			1341 => x"fe9716f5",
			1342 => x"0c045c04",
			1343 => x"000016f5",
			1344 => x"01a216f5",
			1345 => x"08037610",
			1346 => x"0a026708",
			1347 => x"02079204",
			1348 => x"ffa616f5",
			1349 => x"fdf416f5",
			1350 => x"0a027504",
			1351 => x"015c16f5",
			1352 => x"ff8f16f5",
			1353 => x"fdb616f5",
			1354 => x"08038a20",
			1355 => x"040cbf10",
			1356 => x"0304e708",
			1357 => x"0b048e04",
			1358 => x"ffe716f5",
			1359 => x"007316f5",
			1360 => x"0d054d04",
			1361 => x"ffbc16f5",
			1362 => x"001616f5",
			1363 => x"0d050f08",
			1364 => x"0004a004",
			1365 => x"000016f5",
			1366 => x"01b716f5",
			1367 => x"06014204",
			1368 => x"fe3f16f5",
			1369 => x"ffef16f5",
			1370 => x"0d050f04",
			1371 => x"ff8216f5",
			1372 => x"0304ef04",
			1373 => x"010216f5",
			1374 => x"020916f5",
			1375 => x"0900a62c",
			1376 => x"03053718",
			1377 => x"09008d10",
			1378 => x"040ca708",
			1379 => x"0004a704",
			1380 => x"fde916f5",
			1381 => x"ffd416f5",
			1382 => x"0c049104",
			1383 => x"010f16f5",
			1384 => x"ff1c16f5",
			1385 => x"09009e04",
			1386 => x"019016f5",
			1387 => x"001616f5",
			1388 => x"0e04ad08",
			1389 => x"0e04a504",
			1390 => x"ff8016f5",
			1391 => x"fcc816f5",
			1392 => x"0e04cc04",
			1393 => x"01a416f5",
			1394 => x"0a02cc04",
			1395 => x"feac16f5",
			1396 => x"00da16f5",
			1397 => x"06016318",
			1398 => x"0305a90c",
			1399 => x"0e052d08",
			1400 => x"0c04af04",
			1401 => x"019b16f5",
			1402 => x"ffcc16f5",
			1403 => x"fe0516f5",
			1404 => x"0f07c704",
			1405 => x"01eb16f5",
			1406 => x"0d05ab04",
			1407 => x"017d16f5",
			1408 => x"ffa416f5",
			1409 => x"0704ec0c",
			1410 => x"0305b004",
			1411 => x"00f816f5",
			1412 => x"0d05b504",
			1413 => x"fe0516f5",
			1414 => x"ff5516f5",
			1415 => x"0d05cf04",
			1416 => x"017516f5",
			1417 => x"040cbf04",
			1418 => x"ff4816f5",
			1419 => x"005316f5",
			1420 => x"0c04762c",
			1421 => x"0304d628",
			1422 => x"0304871c",
			1423 => x"0a02d10c",
			1424 => x"0c043c04",
			1425 => x"000016f5",
			1426 => x"06013504",
			1427 => x"000016f5",
			1428 => x"019716f5",
			1429 => x"0d04e508",
			1430 => x"0c045e04",
			1431 => x"fffd16f5",
			1432 => x"fd6016f5",
			1433 => x"03043704",
			1434 => x"010116f5",
			1435 => x"ff6816f5",
			1436 => x"0004c904",
			1437 => x"000016f5",
			1438 => x"0d04f304",
			1439 => x"007f16f5",
			1440 => x"fda816f5",
			1441 => x"01ad16f5",
			1442 => x"07049710",
			1443 => x"09005d0c",
			1444 => x"0f05fc08",
			1445 => x"09003204",
			1446 => x"000016f5",
			1447 => x"017b16f5",
			1448 => x"fe5616f5",
			1449 => x"019916f5",
			1450 => x"0b04b214",
			1451 => x"0900890c",
			1452 => x"040d5504",
			1453 => x"018916f5",
			1454 => x"06014104",
			1455 => x"010d16f5",
			1456 => x"ff3716f5",
			1457 => x"02089d04",
			1458 => x"fd2316f5",
			1459 => x"000016f5",
			1460 => x"0d056604",
			1461 => x"01a216f5",
			1462 => x"09008908",
			1463 => x"06013e04",
			1464 => x"001216f5",
			1465 => x"fe8e16f5",
			1466 => x"0803a304",
			1467 => x"000016f5",
			1468 => x"011116f5",
			1469 => x"0e053b98",
			1470 => x"0f06d65c",
			1471 => x"06012528",
			1472 => x"0d054118",
			1473 => x"0304ef10",
			1474 => x"00041408",
			1475 => x"0802d204",
			1476 => x"fde41951",
			1477 => x"01691951",
			1478 => x"07049504",
			1479 => x"ff3f1951",
			1480 => x"01931951",
			1481 => x"0e047104",
			1482 => x"fed11951",
			1483 => x"fd6d1951",
			1484 => x"05053a04",
			1485 => x"00191951",
			1486 => x"00032c04",
			1487 => x"00001951",
			1488 => x"08030104",
			1489 => x"01bd1951",
			1490 => x"008c1951",
			1491 => x"03052520",
			1492 => x"0b04bf10",
			1493 => x"05051e08",
			1494 => x"0b049104",
			1495 => x"ffcc1951",
			1496 => x"00c11951",
			1497 => x"05052004",
			1498 => x"fedf1951",
			1499 => x"ffb21951",
			1500 => x"0f06ac08",
			1501 => x"00042d04",
			1502 => x"fef51951",
			1503 => x"005d1951",
			1504 => x"01005804",
			1505 => x"00461951",
			1506 => x"018f1951",
			1507 => x"02082410",
			1508 => x"0207f808",
			1509 => x"0207cf04",
			1510 => x"fecc1951",
			1511 => x"00001951",
			1512 => x"05056b04",
			1513 => x"fd5b1951",
			1514 => x"fe821951",
			1515 => x"00f51951",
			1516 => x"0803a32c",
			1517 => x"040d551c",
			1518 => x"0d050c0c",
			1519 => x"040c0404",
			1520 => x"fceb1951",
			1521 => x"040c7f04",
			1522 => x"01091951",
			1523 => x"feb41951",
			1524 => x"0304fe08",
			1525 => x"0004b004",
			1526 => x"00e01951",
			1527 => x"ff881951",
			1528 => x"00044b04",
			1529 => x"00451951",
			1530 => x"fff21951",
			1531 => x"0f074908",
			1532 => x"07048004",
			1533 => x"00001951",
			1534 => x"fcc81951",
			1535 => x"08037e04",
			1536 => x"00001951",
			1537 => x"015c1951",
			1538 => x"040f0208",
			1539 => x"02090c04",
			1540 => x"01af1951",
			1541 => x"00af1951",
			1542 => x"05057604",
			1543 => x"00001951",
			1544 => x"fe541951",
			1545 => x"0305c848",
			1546 => x"0c04ac20",
			1547 => x"0c049610",
			1548 => x"0f07dc0c",
			1549 => x"040a1504",
			1550 => x"067f1951",
			1551 => x"0f07ce04",
			1552 => x"ff671951",
			1553 => x"fd6f1951",
			1554 => x"01f71951",
			1555 => x"0c049708",
			1556 => x"040b3604",
			1557 => x"ff511951",
			1558 => x"fd8c1951",
			1559 => x"0f079104",
			1560 => x"fe3e1951",
			1561 => x"ffea1951",
			1562 => x"0b04e114",
			1563 => x"08031a04",
			1564 => x"fe681951",
			1565 => x"0e055a08",
			1566 => x"08034f04",
			1567 => x"01231951",
			1568 => x"ff3d1951",
			1569 => x"0c04b104",
			1570 => x"ffdb1951",
			1571 => x"02d11951",
			1572 => x"0207e508",
			1573 => x"0600da04",
			1574 => x"00001951",
			1575 => x"03cb1951",
			1576 => x"0c04af04",
			1577 => x"00e11951",
			1578 => x"0e057f04",
			1579 => x"ff731951",
			1580 => x"fdad1951",
			1581 => x"0305cc14",
			1582 => x"0004640c",
			1583 => x"0d05a804",
			1584 => x"033c1951",
			1585 => x"040b7604",
			1586 => x"ff771951",
			1587 => x"02641951",
			1588 => x"0f07ac04",
			1589 => x"fea01951",
			1590 => x"01e01951",
			1591 => x"06015b20",
			1592 => x"02090510",
			1593 => x"040c2c08",
			1594 => x"06014204",
			1595 => x"006c1951",
			1596 => x"ff991951",
			1597 => x"040c7904",
			1598 => x"013b1951",
			1599 => x"ff2f1951",
			1600 => x"0704d808",
			1601 => x"0d059a04",
			1602 => x"00a31951",
			1603 => x"02871951",
			1604 => x"06015604",
			1605 => x"ffe41951",
			1606 => x"01861951",
			1607 => x"0505a10c",
			1608 => x"02094d08",
			1609 => x"0e05b304",
			1610 => x"fe151951",
			1611 => x"ffb51951",
			1612 => x"00a21951",
			1613 => x"0f080508",
			1614 => x"02090504",
			1615 => x"00191951",
			1616 => x"018a1951",
			1617 => x"0e06ac04",
			1618 => x"ff231951",
			1619 => x"00031951",
			1620 => x"0d0611bc",
			1621 => x"0f06d644",
			1622 => x"0e04c934",
			1623 => x"040eab20",
			1624 => x"03044e10",
			1625 => x"07047d08",
			1626 => x"03041f04",
			1627 => x"01681b55",
			1628 => x"ffba1b55",
			1629 => x"0f05e004",
			1630 => x"00ee1b55",
			1631 => x"01dc1b55",
			1632 => x"0704c108",
			1633 => x"0c049604",
			1634 => x"00011b55",
			1635 => x"ff4f1b55",
			1636 => x"0704c404",
			1637 => x"01931b55",
			1638 => x"00141b55",
			1639 => x"0601560c",
			1640 => x"040fc604",
			1641 => x"fda01b55",
			1642 => x"04112a04",
			1643 => x"005a1b55",
			1644 => x"fe6d1b55",
			1645 => x"0a03bf04",
			1646 => x"014a1b55",
			1647 => x"00001b55",
			1648 => x"06012508",
			1649 => x"02076704",
			1650 => x"fded1b55",
			1651 => x"01811b55",
			1652 => x"0c048f04",
			1653 => x"ffe11b55",
			1654 => x"fdbd1b55",
			1655 => x"0a02853c",
			1656 => x"02085b20",
			1657 => x"03054310",
			1658 => x"09008c08",
			1659 => x"03051b04",
			1660 => x"008a1b55",
			1661 => x"fe621b55",
			1662 => x"0c047404",
			1663 => x"031f1b55",
			1664 => x"01391b55",
			1665 => x"09009508",
			1666 => x"0f071f04",
			1667 => x"fdd41b55",
			1668 => x"ffdc1b55",
			1669 => x"0a026504",
			1670 => x"00a11b55",
			1671 => x"ffcc1b55",
			1672 => x"0208600c",
			1673 => x"03059708",
			1674 => x"040b8504",
			1675 => x"04541b55",
			1676 => x"01991b55",
			1677 => x"006d1b55",
			1678 => x"06013008",
			1679 => x"0e050004",
			1680 => x"00001b55",
			1681 => x"fe6d1b55",
			1682 => x"0c04ea04",
			1683 => x"00fd1b55",
			1684 => x"fedd1b55",
			1685 => x"0e04961c",
			1686 => x"0c047210",
			1687 => x"06014108",
			1688 => x"0f06ea04",
			1689 => x"00a81b55",
			1690 => x"fe561b55",
			1691 => x"0208a404",
			1692 => x"01911b55",
			1693 => x"ff121b55",
			1694 => x"00044204",
			1695 => x"ff371b55",
			1696 => x"0a029504",
			1697 => x"01a31b55",
			1698 => x"00af1b55",
			1699 => x"09009510",
			1700 => x"0f073b08",
			1701 => x"03051b04",
			1702 => x"006e1b55",
			1703 => x"fe7d1b55",
			1704 => x"0a029b04",
			1705 => x"01671b55",
			1706 => x"ff9d1b55",
			1707 => x"0e04bb08",
			1708 => x"06014104",
			1709 => x"02411b55",
			1710 => x"00e01b55",
			1711 => x"040c7f04",
			1712 => x"00011b55",
			1713 => x"00b01b55",
			1714 => x"0003a614",
			1715 => x"0b058710",
			1716 => x"0802be0c",
			1717 => x"07052f04",
			1718 => x"fe6b1b55",
			1719 => x"07053104",
			1720 => x"00ae1b55",
			1721 => x"ff121b55",
			1722 => x"00641b55",
			1723 => x"fe601b55",
			1724 => x"04110330",
			1725 => x"0900dc14",
			1726 => x"0c04f10c",
			1727 => x"0d061d04",
			1728 => x"ff981b55",
			1729 => x"07051804",
			1730 => x"feec1b55",
			1731 => x"fd201b55",
			1732 => x"06015e04",
			1733 => x"ff471b55",
			1734 => x"01c91b55",
			1735 => x"0705180c",
			1736 => x"0e065a04",
			1737 => x"01fc1b55",
			1738 => x"040b5d04",
			1739 => x"fdc91b55",
			1740 => x"ffb61b55",
			1741 => x"0e060008",
			1742 => x"0a02b104",
			1743 => x"fd261b55",
			1744 => x"00001b55",
			1745 => x"0d062a04",
			1746 => x"01d91b55",
			1747 => x"00021b55",
			1748 => x"fe6c1b55",
			1749 => x"0c047988",
			1750 => x"09008a4c",
			1751 => x"03050030",
			1752 => x"0704a720",
			1753 => x"00040210",
			1754 => x"05051408",
			1755 => x"040b2204",
			1756 => x"feb91db1",
			1757 => x"fadf1db1",
			1758 => x"0c047404",
			1759 => x"01a21db1",
			1760 => x"ffe71db1",
			1761 => x"01003f08",
			1762 => x"03042604",
			1763 => x"00f31db1",
			1764 => x"ff051db1",
			1765 => x"0304a704",
			1766 => x"00c41db1",
			1767 => x"fff61db1",
			1768 => x"0c047404",
			1769 => x"01ca1db1",
			1770 => x"06013a08",
			1771 => x"06012d04",
			1772 => x"012e1db1",
			1773 => x"ff121db1",
			1774 => x"01ba1db1",
			1775 => x"08038818",
			1776 => x"0e047f0c",
			1777 => x"0c047408",
			1778 => x"02089304",
			1779 => x"ffc01db1",
			1780 => x"fd511db1",
			1781 => x"fd541db1",
			1782 => x"040c9308",
			1783 => x"00042404",
			1784 => x"fd2d1db1",
			1785 => x"fffa1db1",
			1786 => x"fd181db1",
			1787 => x"01671db1",
			1788 => x"05052d14",
			1789 => x"0b04b010",
			1790 => x"0e04e20c",
			1791 => x"0e046804",
			1792 => x"fff21db1",
			1793 => x"06013d04",
			1794 => x"01021db1",
			1795 => x"02451db1",
			1796 => x"ffb91db1",
			1797 => x"03291db1",
			1798 => x"0c047210",
			1799 => x"0a027004",
			1800 => x"013d1db1",
			1801 => x"0c045b04",
			1802 => x"00351db1",
			1803 => x"03054304",
			1804 => x"fd271db1",
			1805 => x"febc1db1",
			1806 => x"0704c410",
			1807 => x"0e050708",
			1808 => x"0900a204",
			1809 => x"00b31db1",
			1810 => x"02e31db1",
			1811 => x"0305a004",
			1812 => x"ff651db1",
			1813 => x"01101db1",
			1814 => x"05056804",
			1815 => x"fda71db1",
			1816 => x"00001db1",
			1817 => x"0c048f34",
			1818 => x"0a027a14",
			1819 => x"07049304",
			1820 => x"fde61db1",
			1821 => x"01005708",
			1822 => x"06012b04",
			1823 => x"00421db1",
			1824 => x"02971db1",
			1825 => x"0c047e04",
			1826 => x"00051db1",
			1827 => x"fdcc1db1",
			1828 => x"02089818",
			1829 => x"0704900c",
			1830 => x"0b047104",
			1831 => x"01e41db1",
			1832 => x"03045604",
			1833 => x"fe1a1db1",
			1834 => x"00e01db1",
			1835 => x"01004104",
			1836 => x"011d1db1",
			1837 => x"0e049604",
			1838 => x"fe3a1db1",
			1839 => x"fd521db1",
			1840 => x"06014f04",
			1841 => x"010f1db1",
			1842 => x"fe9a1db1",
			1843 => x"03052538",
			1844 => x"0900951c",
			1845 => x"01005910",
			1846 => x"05053108",
			1847 => x"03050d04",
			1848 => x"00201db1",
			1849 => x"fefd1db1",
			1850 => x"0207fa04",
			1851 => x"ffd21db1",
			1852 => x"00f31db1",
			1853 => x"06015108",
			1854 => x"0704bb04",
			1855 => x"00331db1",
			1856 => x"fe961db1",
			1857 => x"01cc1db1",
			1858 => x"08032e0c",
			1859 => x"040b3608",
			1860 => x"0207af04",
			1861 => x"00131db1",
			1862 => x"01f01db1",
			1863 => x"fe491db1",
			1864 => x"040c3208",
			1865 => x"040bb004",
			1866 => x"02eb1db1",
			1867 => x"01c81db1",
			1868 => x"06015204",
			1869 => x"ffe41db1",
			1870 => x"019b1db1",
			1871 => x"09009c1c",
			1872 => x"03057910",
			1873 => x"0208bb08",
			1874 => x"03052704",
			1875 => x"fe4b1db1",
			1876 => x"ffa71db1",
			1877 => x"0a02c604",
			1878 => x"01e01db1",
			1879 => x"ff981db1",
			1880 => x"040ceb08",
			1881 => x"0a02bc04",
			1882 => x"fed11db1",
			1883 => x"fc0b1db1",
			1884 => x"019b1db1",
			1885 => x"01006210",
			1886 => x"03058908",
			1887 => x"02082f04",
			1888 => x"00001db1",
			1889 => x"01701db1",
			1890 => x"0b04c304",
			1891 => x"015f1db1",
			1892 => x"ff181db1",
			1893 => x"0900a708",
			1894 => x"08036c04",
			1895 => x"ff361db1",
			1896 => x"005e1db1",
			1897 => x"0b04ce04",
			1898 => x"011b1db1",
			1899 => x"00141db1",
			1900 => x"0e053ba0",
			1901 => x"0f06d65c",
			1902 => x"06012528",
			1903 => x"0d054118",
			1904 => x"0304f710",
			1905 => x"0504f208",
			1906 => x"0f060a04",
			1907 => x"00052015",
			1908 => x"fce22015",
			1909 => x"0a027d04",
			1910 => x"00f82015",
			1911 => x"feec2015",
			1912 => x"0003cf04",
			1913 => x"fc992015",
			1914 => x"fe1f2015",
			1915 => x"05053104",
			1916 => x"00002015",
			1917 => x"00032c04",
			1918 => x"fff62015",
			1919 => x"0f06bb04",
			1920 => x"01ca2015",
			1921 => x"00e82015",
			1922 => x"03052520",
			1923 => x"0b04bf10",
			1924 => x"05051e08",
			1925 => x"05051404",
			1926 => x"ffde2015",
			1927 => x"01052015",
			1928 => x"0e04a004",
			1929 => x"ff662015",
			1930 => x"01232015",
			1931 => x"0f069908",
			1932 => x"03050004",
			1933 => x"00112015",
			1934 => x"fd7e2015",
			1935 => x"0304fe04",
			1936 => x"01ab2015",
			1937 => x"00712015",
			1938 => x"0d05bd10",
			1939 => x"01006408",
			1940 => x"0d058e04",
			1941 => x"fef92015",
			1942 => x"00a82015",
			1943 => x"01006c04",
			1944 => x"fe5f2015",
			1945 => x"fd4e2015",
			1946 => x"00a82015",
			1947 => x"0900bc2c",
			1948 => x"0b052220",
			1949 => x"0304fe10",
			1950 => x"0d050d08",
			1951 => x"0f071704",
			1952 => x"fee12015",
			1953 => x"01ab2015",
			1954 => x"0004b004",
			1955 => x"010b2015",
			1956 => x"ff802015",
			1957 => x"09007d08",
			1958 => x"0b04b004",
			1959 => x"fdf02015",
			1960 => x"01252015",
			1961 => x"09009804",
			1962 => x"fffb2015",
			1963 => x"00582015",
			1964 => x"07050804",
			1965 => x"fcbd2015",
			1966 => x"0506b604",
			1967 => x"01402015",
			1968 => x"00002015",
			1969 => x"06015208",
			1970 => x"0e052604",
			1971 => x"02d02015",
			1972 => x"010e2015",
			1973 => x"0f077908",
			1974 => x"0305b604",
			1975 => x"01902015",
			1976 => x"00082015",
			1977 => x"020a0004",
			1978 => x"fc352015",
			1979 => x"00002015",
			1980 => x"0003ea38",
			1981 => x"09014330",
			1982 => x"040adc1c",
			1983 => x"0003d10c",
			1984 => x"040abb08",
			1985 => x"06015a04",
			1986 => x"fff72015",
			1987 => x"01bd2015",
			1988 => x"025e2015",
			1989 => x"0a027a08",
			1990 => x"05059504",
			1991 => x"ff722015",
			1992 => x"fe042015",
			1993 => x"06017404",
			1994 => x"01422015",
			1995 => x"ff992015",
			1996 => x"06013504",
			1997 => x"fd942015",
			1998 => x"0208bb08",
			1999 => x"02086204",
			2000 => x"01ac2015",
			2001 => x"03462015",
			2002 => x"0e06ce04",
			2003 => x"fff32015",
			2004 => x"012b2015",
			2005 => x"0a02a004",
			2006 => x"fe702015",
			2007 => x"00592015",
			2008 => x"02088520",
			2009 => x"03058004",
			2010 => x"02ce2015",
			2011 => x"06015210",
			2012 => x"0d05a708",
			2013 => x"0d059004",
			2014 => x"fe3a2015",
			2015 => x"006c2015",
			2016 => x"0a029204",
			2017 => x"fe092015",
			2018 => x"ffc82015",
			2019 => x"0900b104",
			2020 => x"02c92015",
			2021 => x"0900b904",
			2022 => x"fd9e2015",
			2023 => x"006e2015",
			2024 => x"06014a1c",
			2025 => x"0f079d0c",
			2026 => x"0b04df04",
			2027 => x"fe3b2015",
			2028 => x"0f078704",
			2029 => x"017e2015",
			2030 => x"ffc72015",
			2031 => x"0e056808",
			2032 => x"0a029304",
			2033 => x"02a82015",
			2034 => x"004e2015",
			2035 => x"0208dd04",
			2036 => x"ffd12015",
			2037 => x"01e22015",
			2038 => x"0900c610",
			2039 => x"0f078708",
			2040 => x"040be404",
			2041 => x"ff6e2015",
			2042 => x"01572015",
			2043 => x"0505ce04",
			2044 => x"ff3f2015",
			2045 => x"013b2015",
			2046 => x"03061108",
			2047 => x"0208b904",
			2048 => x"007c2015",
			2049 => x"026c2015",
			2050 => x"040b2404",
			2051 => x"fee32015",
			2052 => x"ffdf2015",
			2053 => x"080329b0",
			2054 => x"08031d5c",
			2055 => x"0d053328",
			2056 => x"07049218",
			2057 => x"0304f710",
			2058 => x"00041408",
			2059 => x"0b048d04",
			2060 => x"ff772299",
			2061 => x"01a12299",
			2062 => x"0f06bb04",
			2063 => x"fda92299",
			2064 => x"014d2299",
			2065 => x"00041404",
			2066 => x"fdce2299",
			2067 => x"00d82299",
			2068 => x"0207c50c",
			2069 => x"03049704",
			2070 => x"00002299",
			2071 => x"0d052604",
			2072 => x"fc132299",
			2073 => x"fdf02299",
			2074 => x"008d2299",
			2075 => x"0100731c",
			2076 => x"0b050110",
			2077 => x"07049008",
			2078 => x"01005104",
			2079 => x"00a92299",
			2080 => x"fd4f2299",
			2081 => x"0b04b004",
			2082 => x"01592299",
			2083 => x"000d2299",
			2084 => x"0207da04",
			2085 => x"fef12299",
			2086 => x"040b0f04",
			2087 => x"02952299",
			2088 => x"00c12299",
			2089 => x"0d05a808",
			2090 => x"05058404",
			2091 => x"ffc92299",
			2092 => x"fd642299",
			2093 => x"040b5608",
			2094 => x"0003e504",
			2095 => x"fffe2299",
			2096 => x"fe5b2299",
			2097 => x"0c054304",
			2098 => x"02b02299",
			2099 => x"fecd2299",
			2100 => x"02084530",
			2101 => x"01006420",
			2102 => x"0f06ac10",
			2103 => x"0f068708",
			2104 => x"05052e04",
			2105 => x"01a12299",
			2106 => x"ff422299",
			2107 => x"05051e04",
			2108 => x"00002299",
			2109 => x"fdc32299",
			2110 => x"03051f08",
			2111 => x"06012804",
			2112 => x"001c2299",
			2113 => x"02082299",
			2114 => x"0704c104",
			2115 => x"ffce2299",
			2116 => x"020b2299",
			2117 => x"0900b50c",
			2118 => x"08032004",
			2119 => x"ff682299",
			2120 => x"03056804",
			2121 => x"fce82299",
			2122 => x"fe6a2299",
			2123 => x"01482299",
			2124 => x"01007d14",
			2125 => x"03061110",
			2126 => x"01007108",
			2127 => x"0d058d04",
			2128 => x"00f12299",
			2129 => x"025b2299",
			2130 => x"01007604",
			2131 => x"fe4f2299",
			2132 => x"00322299",
			2133 => x"04392299",
			2134 => x"06015a04",
			2135 => x"fe0f2299",
			2136 => x"0c04cc04",
			2137 => x"02a22299",
			2138 => x"07050804",
			2139 => x"ff582299",
			2140 => x"00a62299",
			2141 => x"02086c48",
			2142 => x"08032e14",
			2143 => x"0f074f10",
			2144 => x"0c045b04",
			2145 => x"fd332299",
			2146 => x"00041d04",
			2147 => x"fe042299",
			2148 => x"08032b04",
			2149 => x"fd942299",
			2150 => x"004e2299",
			2151 => x"00de2299",
			2152 => x"08033114",
			2153 => x"0c04960c",
			2154 => x"02080204",
			2155 => x"005d2299",
			2156 => x"03051f04",
			2157 => x"01782299",
			2158 => x"02bc2299",
			2159 => x"0d057604",
			2160 => x"fd302299",
			2161 => x"014f2299",
			2162 => x"03057910",
			2163 => x"0d058308",
			2164 => x"07049704",
			2165 => x"00022299",
			2166 => x"ffa72299",
			2167 => x"0c04b304",
			2168 => x"ffff2299",
			2169 => x"01a52299",
			2170 => x"0900b908",
			2171 => x"08033604",
			2172 => x"00782299",
			2173 => x"fe9c2299",
			2174 => x"01007604",
			2175 => x"01952299",
			2176 => x"ff662299",
			2177 => x"02086e0c",
			2178 => x"06014f08",
			2179 => x"0b04e304",
			2180 => x"022e2299",
			2181 => x"ffc22299",
			2182 => x"fe802299",
			2183 => x"040c5e20",
			2184 => x"08037410",
			2185 => x"0704da08",
			2186 => x"0704d504",
			2187 => x"00002299",
			2188 => x"00cd2299",
			2189 => x"0505a304",
			2190 => x"ff202299",
			2191 => x"fff52299",
			2192 => x"0900b308",
			2193 => x"09009504",
			2194 => x"01422299",
			2195 => x"fdfc2299",
			2196 => x"0f07b904",
			2197 => x"015d2299",
			2198 => x"ff632299",
			2199 => x"08035310",
			2200 => x"0b04df08",
			2201 => x"00046b04",
			2202 => x"f2602299",
			2203 => x"00002299",
			2204 => x"08034c04",
			2205 => x"fdb42299",
			2206 => x"00002299",
			2207 => x"0c047508",
			2208 => x"0c045b04",
			2209 => x"00092299",
			2210 => x"fee92299",
			2211 => x"08038504",
			2212 => x"00b12299",
			2213 => x"001a2299",
			2214 => x"0208d4b0",
			2215 => x"0c04d064",
			2216 => x"0b04e230",
			2217 => x"0d058214",
			2218 => x"0900b510",
			2219 => x"0d057308",
			2220 => x"0c04b404",
			2221 => x"00042545",
			2222 => x"ff222545",
			2223 => x"0c047404",
			2224 => x"01d92545",
			2225 => x"ff6e2545",
			2226 => x"02272545",
			2227 => x"0505750c",
			2228 => x"09009b04",
			2229 => x"ff6b2545",
			2230 => x"040b6b04",
			2231 => x"00042545",
			2232 => x"01fd2545",
			2233 => x"0b04cf08",
			2234 => x"0d058f04",
			2235 => x"fd5b2545",
			2236 => x"00002545",
			2237 => x"0e051604",
			2238 => x"00ed2545",
			2239 => x"ffe12545",
			2240 => x"0c04ac14",
			2241 => x"06013008",
			2242 => x"040aa904",
			2243 => x"00922545",
			2244 => x"02132545",
			2245 => x"040c7208",
			2246 => x"00046704",
			2247 => x"fede2545",
			2248 => x"008a2545",
			2249 => x"fc9f2545",
			2250 => x"0c04af10",
			2251 => x"02087608",
			2252 => x"0e04f704",
			2253 => x"01ce2545",
			2254 => x"ff132545",
			2255 => x"0a029904",
			2256 => x"02af2545",
			2257 => x"006f2545",
			2258 => x"06016208",
			2259 => x"0c04b104",
			2260 => x"ff132545",
			2261 => x"ffc22545",
			2262 => x"06016404",
			2263 => x"02582545",
			2264 => x"ff732545",
			2265 => x"0c04d120",
			2266 => x"0a02a310",
			2267 => x"0208ab0c",
			2268 => x"06014d08",
			2269 => x"01006a04",
			2270 => x"02052545",
			2271 => x"009b2545",
			2272 => x"03e72545",
			2273 => x"00322545",
			2274 => x"0a02b308",
			2275 => x"0e055204",
			2276 => x"fe712545",
			2277 => x"00042545",
			2278 => x"0704da04",
			2279 => x"001e2545",
			2280 => x"022d2545",
			2281 => x"06014d1c",
			2282 => x"0601420c",
			2283 => x"05058404",
			2284 => x"feab2545",
			2285 => x"0409b304",
			2286 => x"ff162545",
			2287 => x"01042545",
			2288 => x"040c1208",
			2289 => x"0505af04",
			2290 => x"00032545",
			2291 => x"fe982545",
			2292 => x"0208c904",
			2293 => x"fdcb2545",
			2294 => x"fb9a2545",
			2295 => x"06014e04",
			2296 => x"02fe2545",
			2297 => x"05058604",
			2298 => x"feb02545",
			2299 => x"01006e04",
			2300 => x"02822545",
			2301 => x"001f2545",
			2302 => x"0c04cc4c",
			2303 => x"0900b528",
			2304 => x"0b050320",
			2305 => x"06015310",
			2306 => x"0e057808",
			2307 => x"0c048f04",
			2308 => x"ffe82545",
			2309 => x"01572545",
			2310 => x"0c049604",
			2311 => x"00442545",
			2312 => x"fe332545",
			2313 => x"0704bb08",
			2314 => x"03058904",
			2315 => x"00692545",
			2316 => x"fe562545",
			2317 => x"0704d304",
			2318 => x"00c62545",
			2319 => x"ff252545",
			2320 => x"0e056104",
			2321 => x"ff5c2545",
			2322 => x"fdd22545",
			2323 => x"0306ff20",
			2324 => x"0a02a610",
			2325 => x"03061908",
			2326 => x"0900c404",
			2327 => x"01802545",
			2328 => x"032e2545",
			2329 => x"0505bd04",
			2330 => x"ffb22545",
			2331 => x"01822545",
			2332 => x"0704d408",
			2333 => x"0a02bf04",
			2334 => x"febd2545",
			2335 => x"00e62545",
			2336 => x"040c6004",
			2337 => x"00a32545",
			2338 => x"01b22545",
			2339 => x"fdf82545",
			2340 => x"07050324",
			2341 => x"0e057110",
			2342 => x"0a02ac04",
			2343 => x"fea02545",
			2344 => x"00048a04",
			2345 => x"02162545",
			2346 => x"00049c04",
			2347 => x"ff942545",
			2348 => x"01852545",
			2349 => x"0a028b04",
			2350 => x"02352545",
			2351 => x"040be908",
			2352 => x"00043a04",
			2353 => x"fef72545",
			2354 => x"fdd32545",
			2355 => x"040bff04",
			2356 => x"01672545",
			2357 => x"ff442545",
			2358 => x"040b1418",
			2359 => x"09011b0c",
			2360 => x"0c04e904",
			2361 => x"fe1d2545",
			2362 => x"06017304",
			2363 => x"00002545",
			2364 => x"01c62545",
			2365 => x"05068a04",
			2366 => x"fe072545",
			2367 => x"0506f104",
			2368 => x"00082545",
			2369 => x"fe962545",
			2370 => x"00040b10",
			2371 => x"0901f608",
			2372 => x"0003ab04",
			2373 => x"05762545",
			2374 => x"01882545",
			2375 => x"07070c04",
			2376 => x"febb2545",
			2377 => x"00782545",
			2378 => x"0b053308",
			2379 => x"00046404",
			2380 => x"01dd2545",
			2381 => x"00002545",
			2382 => x"0a02a804",
			2383 => x"fef82545",
			2384 => x"00362545",
			2385 => x"0e04bbb8",
			2386 => x"0f070570",
			2387 => x"040c6030",
			2388 => x"01004d18",
			2389 => x"0a02b110",
			2390 => x"06013a08",
			2391 => x"02084504",
			2392 => x"00692831",
			2393 => x"ff2c2831",
			2394 => x"00045204",
			2395 => x"00002831",
			2396 => x"01942831",
			2397 => x"0e03da04",
			2398 => x"fda22831",
			2399 => x"00002831",
			2400 => x"0704a80c",
			2401 => x"00048608",
			2402 => x"0d051904",
			2403 => x"fddf2831",
			2404 => x"ffc52831",
			2405 => x"01c52831",
			2406 => x"040c5808",
			2407 => x"0f06ed04",
			2408 => x"00232831",
			2409 => x"00c92831",
			2410 => x"fec92831",
			2411 => x"08037620",
			2412 => x"06013010",
			2413 => x"03048708",
			2414 => x"03043e04",
			2415 => x"006b2831",
			2416 => x"fd532831",
			2417 => x"01004104",
			2418 => x"00002831",
			2419 => x"01de2831",
			2420 => x"0e043d08",
			2421 => x"0d052504",
			2422 => x"fe992831",
			2423 => x"01ad2831",
			2424 => x"00047904",
			2425 => x"ff492831",
			2426 => x"fd642831",
			2427 => x"0d055a10",
			2428 => x"040cc608",
			2429 => x"01004104",
			2430 => x"ff472831",
			2431 => x"00cc2831",
			2432 => x"0f06f304",
			2433 => x"ffeb2831",
			2434 => x"fe012831",
			2435 => x"0a02bf08",
			2436 => x"0b04cf04",
			2437 => x"fd2b2831",
			2438 => x"ff5a2831",
			2439 => x"040d6e04",
			2440 => x"01262831",
			2441 => x"fe332831",
			2442 => x"0d055924",
			2443 => x"03053918",
			2444 => x"01005a10",
			2445 => x"0e04ad08",
			2446 => x"0208ad04",
			2447 => x"008f2831",
			2448 => x"ff642831",
			2449 => x"00048e04",
			2450 => x"01ba2831",
			2451 => x"00012831",
			2452 => x"0b04b904",
			2453 => x"00b62831",
			2454 => x"fe482831",
			2455 => x"0f076508",
			2456 => x"0e04a904",
			2457 => x"fc362831",
			2458 => x"fec42831",
			2459 => x"00002831",
			2460 => x"05057618",
			2461 => x"05054b0c",
			2462 => x"0b04ce08",
			2463 => x"0704a704",
			2464 => x"ffa92831",
			2465 => x"01d72831",
			2466 => x"fe162831",
			2467 => x"08033704",
			2468 => x"00002831",
			2469 => x"08039304",
			2470 => x"01ac2831",
			2471 => x"00732831",
			2472 => x"01006104",
			2473 => x"fcd82831",
			2474 => x"040cf504",
			2475 => x"01a32831",
			2476 => x"ff402831",
			2477 => x"0d058358",
			2478 => x"05057638",
			2479 => x"01006620",
			2480 => x"0f072b10",
			2481 => x"0b04d108",
			2482 => x"02085904",
			2483 => x"ff4d2831",
			2484 => x"fe112831",
			2485 => x"0d057504",
			2486 => x"01782831",
			2487 => x"ff2a2831",
			2488 => x"01006208",
			2489 => x"03059704",
			2490 => x"005f2831",
			2491 => x"fecd2831",
			2492 => x"05056604",
			2493 => x"ffd52831",
			2494 => x"fd7b2831",
			2495 => x"0e04f70c",
			2496 => x"03056104",
			2497 => x"02cb2831",
			2498 => x"03057704",
			2499 => x"00c12831",
			2500 => x"02162831",
			2501 => x"040c6008",
			2502 => x"06015a04",
			2503 => x"00002831",
			2504 => x"fdcf2831",
			2505 => x"01f72831",
			2506 => x"0305a718",
			2507 => x"0100650c",
			2508 => x"0704c204",
			2509 => x"00df2831",
			2510 => x"0d058104",
			2511 => x"fd962831",
			2512 => x"00002831",
			2513 => x"040c3808",
			2514 => x"03057004",
			2515 => x"ff9f2831",
			2516 => x"fdfe2831",
			2517 => x"fca72831",
			2518 => x"0f07a604",
			2519 => x"01032831",
			2520 => x"ff7d2831",
			2521 => x"0b04e228",
			2522 => x"06013108",
			2523 => x"01006504",
			2524 => x"fdf72831",
			2525 => x"00002831",
			2526 => x"0d05a710",
			2527 => x"0b04e008",
			2528 => x"03057904",
			2529 => x"01d32831",
			2530 => x"00272831",
			2531 => x"03057704",
			2532 => x"ff822831",
			2533 => x"019e2831",
			2534 => x"0a02a808",
			2535 => x"08034c04",
			2536 => x"ff5b2831",
			2537 => x"022f2831",
			2538 => x"040c5204",
			2539 => x"fdc92831",
			2540 => x"00272831",
			2541 => x"0b04f120",
			2542 => x"0a02b110",
			2543 => x"0208bb08",
			2544 => x"01006f04",
			2545 => x"ffca2831",
			2546 => x"fe672831",
			2547 => x"0305f204",
			2548 => x"00d92831",
			2549 => x"02a62831",
			2550 => x"040c9308",
			2551 => x"05058304",
			2552 => x"fcff2831",
			2553 => x"feb02831",
			2554 => x"0305a904",
			2555 => x"fef22831",
			2556 => x"00bf2831",
			2557 => x"05059210",
			2558 => x"0704eb08",
			2559 => x"08036104",
			2560 => x"00902831",
			2561 => x"ff532831",
			2562 => x"0d05a704",
			2563 => x"02f32831",
			2564 => x"01002831",
			2565 => x"0d05a908",
			2566 => x"02090504",
			2567 => x"ff1c2831",
			2568 => x"02062831",
			2569 => x"0305a004",
			2570 => x"01432831",
			2571 => x"fff62831",
			2572 => x"0f0773d4",
			2573 => x"0e046174",
			2574 => x"0b049134",
			2575 => x"01004d1c",
			2576 => x"09007910",
			2577 => x"0c047408",
			2578 => x"07047d04",
			2579 => x"ffe02b07",
			2580 => x"00c22b07",
			2581 => x"0e041604",
			2582 => x"ffc32b07",
			2583 => x"feb72b07",
			2584 => x"0b049008",
			2585 => x"0c047304",
			2586 => x"005e2b07",
			2587 => x"01da2b07",
			2588 => x"ff092b07",
			2589 => x"0c04770c",
			2590 => x"09007d04",
			2591 => x"fec22b07",
			2592 => x"0304c704",
			2593 => x"01e12b07",
			2594 => x"fff42b07",
			2595 => x"0704a808",
			2596 => x"0d053204",
			2597 => x"fd442b07",
			2598 => x"ff1e2b07",
			2599 => x"00ab2b07",
			2600 => x"06014720",
			2601 => x"0e043610",
			2602 => x"09007308",
			2603 => x"01004704",
			2604 => x"00c22b07",
			2605 => x"fcad2b07",
			2606 => x"08032e04",
			2607 => x"003b2b07",
			2608 => x"01602b07",
			2609 => x"09007b08",
			2610 => x"05052004",
			2611 => x"ff8a2b07",
			2612 => x"fd152b07",
			2613 => x"0f069f04",
			2614 => x"ffeb2b07",
			2615 => x"00cc2b07",
			2616 => x"0f06a510",
			2617 => x"0f066608",
			2618 => x"040df504",
			2619 => x"01af2b07",
			2620 => x"fec22b07",
			2621 => x"0704c104",
			2622 => x"fdcd2b07",
			2623 => x"016a2b07",
			2624 => x"0d056608",
			2625 => x"05051e04",
			2626 => x"ff282b07",
			2627 => x"01922b07",
			2628 => x"09008e04",
			2629 => x"fdaa2b07",
			2630 => x"012a2b07",
			2631 => x"0d054f24",
			2632 => x"0c04b420",
			2633 => x"03053310",
			2634 => x"0f06e308",
			2635 => x"0b049004",
			2636 => x"01112b07",
			2637 => x"ff1b2b07",
			2638 => x"0304fe04",
			2639 => x"00d62b07",
			2640 => x"ffe22b07",
			2641 => x"0f074108",
			2642 => x"040b7004",
			2643 => x"ffd62b07",
			2644 => x"fddf2b07",
			2645 => x"08034104",
			2646 => x"02372b07",
			2647 => x"ff522b07",
			2648 => x"fd732b07",
			2649 => x"0e051620",
			2650 => x"0900a810",
			2651 => x"01005c08",
			2652 => x"09009304",
			2653 => x"ffe82b07",
			2654 => x"00f12b07",
			2655 => x"0c04d104",
			2656 => x"ffd52b07",
			2657 => x"fd892b07",
			2658 => x"040ba408",
			2659 => x"03056104",
			2660 => x"01442b07",
			2661 => x"ff4a2b07",
			2662 => x"06015704",
			2663 => x"01882b07",
			2664 => x"001e2b07",
			2665 => x"0900ba10",
			2666 => x"0c049208",
			2667 => x"0c048f04",
			2668 => x"ff8f2b07",
			2669 => x"01612b07",
			2670 => x"0b04d004",
			2671 => x"fe812b07",
			2672 => x"ff672b07",
			2673 => x"08036308",
			2674 => x"01007904",
			2675 => x"00542b07",
			2676 => x"ff492b07",
			2677 => x"021a2b07",
			2678 => x"0704da60",
			2679 => x"0a02b434",
			2680 => x"040bde1c",
			2681 => x"0c04cb10",
			2682 => x"06013508",
			2683 => x"01005904",
			2684 => x"00002b07",
			2685 => x"02202b07",
			2686 => x"040abb04",
			2687 => x"fe3d2b07",
			2688 => x"00002b07",
			2689 => x"0d05de08",
			2690 => x"08034d04",
			2691 => x"02cc2b07",
			2692 => x"00682b07",
			2693 => x"ff052b07",
			2694 => x"0d05330c",
			2695 => x"07047b08",
			2696 => x"0f078e04",
			2697 => x"01352b07",
			2698 => x"00002b07",
			2699 => x"fd972b07",
			2700 => x"0c04d108",
			2701 => x"0d058304",
			2702 => x"009b2b07",
			2703 => x"01692b07",
			2704 => x"ff7d2b07",
			2705 => x"0b050220",
			2706 => x"040c8510",
			2707 => x"05058208",
			2708 => x"0900a704",
			2709 => x"fe7a2b07",
			2710 => x"003d2b07",
			2711 => x"06015b04",
			2712 => x"fd032b07",
			2713 => x"fe712b07",
			2714 => x"0704c008",
			2715 => x"0e04f004",
			2716 => x"01ac2b07",
			2717 => x"ff5e2b07",
			2718 => x"0c049204",
			2719 => x"00002b07",
			2720 => x"01b82b07",
			2721 => x"0c04b104",
			2722 => x"fe7a2b07",
			2723 => x"0e055a04",
			2724 => x"00c32b07",
			2725 => x"02682b07",
			2726 => x"0704ec1c",
			2727 => x"0f078104",
			2728 => x"015e2b07",
			2729 => x"0c04d00c",
			2730 => x"0704ea08",
			2731 => x"0900ba04",
			2732 => x"fe202b07",
			2733 => x"ffcb2b07",
			2734 => x"fdd92b07",
			2735 => x"0c04ec08",
			2736 => x"0505a104",
			2737 => x"01c92b07",
			2738 => x"ffd82b07",
			2739 => x"fd742b07",
			2740 => x"03059904",
			2741 => x"fda92b07",
			2742 => x"0900a708",
			2743 => x"0f079104",
			2744 => x"014b2b07",
			2745 => x"03002b07",
			2746 => x"0c04b408",
			2747 => x"06015604",
			2748 => x"ffdf2b07",
			2749 => x"01232b07",
			2750 => x"0c04b604",
			2751 => x"fec92b07",
			2752 => x"00052b07",
			2753 => x"040f0248",
			2754 => x"04095908",
			2755 => x"07049204",
			2756 => x"00002bd1",
			2757 => x"fe722bd1",
			2758 => x"03041f0c",
			2759 => x"0b045c04",
			2760 => x"ffcf2bd1",
			2761 => x"09006204",
			2762 => x"01e92bd1",
			2763 => x"00ed2bd1",
			2764 => x"09006218",
			2765 => x"03043708",
			2766 => x"0e037004",
			2767 => x"fe722bd1",
			2768 => x"016e2bd1",
			2769 => x"0c043a08",
			2770 => x"0c042104",
			2771 => x"ffae2bd1",
			2772 => x"01872bd1",
			2773 => x"07047e04",
			2774 => x"fdb12bd1",
			2775 => x"ff8d2bd1",
			2776 => x"0e03cb0c",
			2777 => x"02081d08",
			2778 => x"03042e04",
			2779 => x"fe8c2bd1",
			2780 => x"01712bd1",
			2781 => x"fe8f2bd1",
			2782 => x"0f070508",
			2783 => x"0e047804",
			2784 => x"00202bd1",
			2785 => x"ffaa2bd1",
			2786 => x"03055304",
			2787 => x"00772bd1",
			2788 => x"00132bd1",
			2789 => x"0704bc1c",
			2790 => x"0c047814",
			2791 => x"0d04db04",
			2792 => x"fe732bd1",
			2793 => x"0d050c0c",
			2794 => x"02086c08",
			2795 => x"0207d104",
			2796 => x"ff8f2bd1",
			2797 => x"00d92bd1",
			2798 => x"ff8a2bd1",
			2799 => x"fe632bd1",
			2800 => x"02082204",
			2801 => x"ffa72bd1",
			2802 => x"01282bd1",
			2803 => x"fe6b2bd1",
			2804 => x"0900823c",
			2805 => x"0704c034",
			2806 => x"0704bf30",
			2807 => x"0304c71c",
			2808 => x"02086710",
			2809 => x"040c8c08",
			2810 => x"02082204",
			2811 => x"00002ced",
			2812 => x"01192ced",
			2813 => x"0e041604",
			2814 => x"ffc92ced",
			2815 => x"fe712ced",
			2816 => x"09006204",
			2817 => x"feb02ced",
			2818 => x"05050e04",
			2819 => x"01ef2ced",
			2820 => x"00cc2ced",
			2821 => x"05054a10",
			2822 => x"0207d708",
			2823 => x"08031404",
			2824 => x"008c2ced",
			2825 => x"fd3e2ced",
			2826 => x"0c049404",
			2827 => x"ff6a2ced",
			2828 => x"003d2ced",
			2829 => x"01882ced",
			2830 => x"fdbb2ced",
			2831 => x"040e6304",
			2832 => x"01d12ced",
			2833 => x"fee12ced",
			2834 => x"0e042610",
			2835 => x"02074b04",
			2836 => x"ff5d2ced",
			2837 => x"09008408",
			2838 => x"040c1204",
			2839 => x"01ac2ced",
			2840 => x"00002ced",
			2841 => x"01d92ced",
			2842 => x"0c045b14",
			2843 => x"0e04db0c",
			2844 => x"0a028704",
			2845 => x"022a2ced",
			2846 => x"040c5e04",
			2847 => x"00002ced",
			2848 => x"01cb2ced",
			2849 => x"02087c04",
			2850 => x"fe8c2ced",
			2851 => x"01762ced",
			2852 => x"0c047210",
			2853 => x"0208ab0c",
			2854 => x"0d053304",
			2855 => x"fe572ced",
			2856 => x"08035504",
			2857 => x"ffa42ced",
			2858 => x"01492ced",
			2859 => x"fe062ced",
			2860 => x"040c6610",
			2861 => x"00049608",
			2862 => x"08037904",
			2863 => x"fffd2ced",
			2864 => x"ff542ced",
			2865 => x"0e052604",
			2866 => x"01ed2ced",
			2867 => x"00d32ced",
			2868 => x"08036608",
			2869 => x"0704c104",
			2870 => x"00052ced",
			2871 => x"fdf82ced",
			2872 => x"08038504",
			2873 => x"00bd2ced",
			2874 => x"00042ced",
			2875 => x"0c05645c",
			2876 => x"040f7050",
			2877 => x"0409b310",
			2878 => x"0e04f004",
			2879 => x"ff7d2e29",
			2880 => x"0b056904",
			2881 => x"fe112e29",
			2882 => x"0b057404",
			2883 => x"00012e29",
			2884 => x"fe6a2e29",
			2885 => x"0c04b220",
			2886 => x"0e057f10",
			2887 => x"0900b508",
			2888 => x"0e04bb04",
			2889 => x"00662e29",
			2890 => x"00102e29",
			2891 => x"0f075504",
			2892 => x"005d2e29",
			2893 => x"020a2e29",
			2894 => x"0c049608",
			2895 => x"06015f04",
			2896 => x"00b32e29",
			2897 => x"feac2e29",
			2898 => x"0b053304",
			2899 => x"fefa2e29",
			2900 => x"01692e29",
			2901 => x"0c04b410",
			2902 => x"0a028508",
			2903 => x"02086c04",
			2904 => x"01662e29",
			2905 => x"03392e29",
			2906 => x"08033904",
			2907 => x"fe122e29",
			2908 => x"01032e29",
			2909 => x"0c04b508",
			2910 => x"02085204",
			2911 => x"00892e29",
			2912 => x"fda92e29",
			2913 => x"0f07ce04",
			2914 => x"00b62e29",
			2915 => x"00232e29",
			2916 => x"09003d04",
			2917 => x"fe632e29",
			2918 => x"0f062f04",
			2919 => x"011d2e29",
			2920 => x"fe422e29",
			2921 => x"0803260c",
			2922 => x"0e068d08",
			2923 => x"0506a704",
			2924 => x"ffe62e29",
			2925 => x"02162e29",
			2926 => x"fe682e29",
			2927 => x"040eab2c",
			2928 => x"08034710",
			2929 => x"020b1c0c",
			2930 => x"05082108",
			2931 => x"0f0a9204",
			2932 => x"01632e29",
			2933 => x"fe822e29",
			2934 => x"02542e29",
			2935 => x"fe632e29",
			2936 => x"040ce110",
			2937 => x"040c1208",
			2938 => x"0a02b904",
			2939 => x"00782e29",
			2940 => x"feb62e29",
			2941 => x"0e0b9404",
			2942 => x"027e2e29",
			2943 => x"00002e29",
			2944 => x"08037304",
			2945 => x"fe1a2e29",
			2946 => x"0601b304",
			2947 => x"ff052e29",
			2948 => x"01792e29",
			2949 => x"0c057f08",
			2950 => x"04173404",
			2951 => x"01612e29",
			2952 => x"fe842e29",
			2953 => x"fe632e29",
			2954 => x"040f0278",
			2955 => x"0803dc68",
			2956 => x"040d5540",
			2957 => x"0e042620",
			2958 => x"0f065f10",
			2959 => x"0e03cb08",
			2960 => x"0504f204",
			2961 => x"ffd42f45",
			2962 => x"01532f45",
			2963 => x"0704ab04",
			2964 => x"feed2f45",
			2965 => x"01d12f45",
			2966 => x"09007108",
			2967 => x"0e03e704",
			2968 => x"011c2f45",
			2969 => x"ff032f45",
			2970 => x"0704ab04",
			2971 => x"012e2f45",
			2972 => x"ff722f45",
			2973 => x"07047810",
			2974 => x"07046708",
			2975 => x"0c045904",
			2976 => x"fdd62f45",
			2977 => x"01142f45",
			2978 => x"0c045704",
			2979 => x"ffd52f45",
			2980 => x"fd2b2f45",
			2981 => x"0f06d608",
			2982 => x"0b048e04",
			2983 => x"fe902f45",
			2984 => x"ffdd2f45",
			2985 => x"06015304",
			2986 => x"00322f45",
			2987 => x"ffe92f45",
			2988 => x"0f062f08",
			2989 => x"0c047804",
			2990 => x"ff732f45",
			2991 => x"01ed2f45",
			2992 => x"0803a310",
			2993 => x"0a02cb08",
			2994 => x"08038504",
			2995 => x"fdcb2f45",
			2996 => x"00d42f45",
			2997 => x"02096004",
			2998 => x"fb332f45",
			2999 => x"feab2f45",
			3000 => x"0c049508",
			3001 => x"0704a604",
			3002 => x"ff8f2f45",
			3003 => x"fd392f45",
			3004 => x"0a02ed04",
			3005 => x"01b42f45",
			3006 => x"ffa52f45",
			3007 => x"06015304",
			3008 => x"00162f45",
			3009 => x"0a032308",
			3010 => x"0a031504",
			3011 => x"01962f45",
			3012 => x"00002f45",
			3013 => x"024b2f45",
			3014 => x"0704bc14",
			3015 => x"0c04780c",
			3016 => x"05050004",
			3017 => x"fea72f45",
			3018 => x"05050e04",
			3019 => x"00812f45",
			3020 => x"fe802f45",
			3021 => x"04130e04",
			3022 => x"00fe2f45",
			3023 => x"ffea2f45",
			3024 => x"fe6f2f45",
			3025 => x"0e041654",
			3026 => x"040d1b28",
			3027 => x"0208241c",
			3028 => x"0004b014",
			3029 => x"040cc60c",
			3030 => x"08038d08",
			3031 => x"00049204",
			3032 => x"003630f1",
			3033 => x"019430f1",
			3034 => x"fdfe30f1",
			3035 => x"0d051904",
			3036 => x"ffda30f1",
			3037 => x"fc4530f1",
			3038 => x"0a02bf04",
			3039 => x"007230f1",
			3040 => x"019f30f1",
			3041 => x"09005d04",
			3042 => x"fe3130f1",
			3043 => x"00048a04",
			3044 => x"00ea30f1",
			3045 => x"01f030f1",
			3046 => x"09006f24",
			3047 => x"0d051a18",
			3048 => x"05050f10",
			3049 => x"06014108",
			3050 => x"07049104",
			3051 => x"fdae30f1",
			3052 => x"009730f1",
			3053 => x"05050204",
			3054 => x"fff630f1",
			3055 => x"019a30f1",
			3056 => x"09003604",
			3057 => x"000030f1",
			3058 => x"fcb330f1",
			3059 => x"040eab04",
			3060 => x"01b530f1",
			3061 => x"07049404",
			3062 => x"000030f1",
			3063 => x"fea930f1",
			3064 => x"040dca04",
			3065 => x"01cb30f1",
			3066 => x"ffac30f1",
			3067 => x"09007e3c",
			3068 => x"0f069618",
			3069 => x"040bca10",
			3070 => x"040b5608",
			3071 => x"0f065904",
			3072 => x"ff7030f1",
			3073 => x"fd5830f1",
			3074 => x"0e042604",
			3075 => x"020a30f1",
			3076 => x"ff6330f1",
			3077 => x"0a02a604",
			3078 => x"fbbb30f1",
			3079 => x"fdaa30f1",
			3080 => x"0304af04",
			3081 => x"01a530f1",
			3082 => x"0a027710",
			3083 => x"0304d608",
			3084 => x"09007104",
			3085 => x"fe2330f1",
			3086 => x"01f930f1",
			3087 => x"00042804",
			3088 => x"ff3a30f1",
			3089 => x"027e30f1",
			3090 => x"0f06ea08",
			3091 => x"0304df04",
			3092 => x"ff3430f1",
			3093 => x"fd3f30f1",
			3094 => x"02085904",
			3095 => x"017e30f1",
			3096 => x"ffae30f1",
			3097 => x"05051014",
			3098 => x"06013e0c",
			3099 => x"00042004",
			3100 => x"fe5130f1",
			3101 => x"0f06ea04",
			3102 => x"016d30f1",
			3103 => x"ff5f30f1",
			3104 => x"0b049104",
			3105 => x"fda630f1",
			3106 => x"ff2c30f1",
			3107 => x"03052514",
			3108 => x"0d057510",
			3109 => x"0f068708",
			3110 => x"0304df04",
			3111 => x"006730f1",
			3112 => x"fe9530f1",
			3113 => x"07047b04",
			3114 => x"febd30f1",
			3115 => x"006930f1",
			3116 => x"021430f1",
			3117 => x"0f074910",
			3118 => x"09008f08",
			3119 => x"0f073b04",
			3120 => x"fef430f1",
			3121 => x"006530f1",
			3122 => x"0f074104",
			3123 => x"fff630f1",
			3124 => x"ff2630f1",
			3125 => x"03057908",
			3126 => x"00044a04",
			3127 => x"020530f1",
			3128 => x"006c30f1",
			3129 => x"09009e04",
			3130 => x"ff2830f1",
			3131 => x"001430f1",
			3132 => x"0803a36c",
			3133 => x"0a02d14c",
			3134 => x"03044e0c",
			3135 => x"06011904",
			3136 => x"fe553275",
			3137 => x"0b046c04",
			3138 => x"ffe33275",
			3139 => x"01bd3275",
			3140 => x"09007e20",
			3141 => x"0304df10",
			3142 => x"02082408",
			3143 => x"040bb704",
			3144 => x"00483275",
			3145 => x"ff7a3275",
			3146 => x"0c047e04",
			3147 => x"000c3275",
			3148 => x"01733275",
			3149 => x"05051f08",
			3150 => x"06014104",
			3151 => x"ff283275",
			3152 => x"01743275",
			3153 => x"0e046b04",
			3154 => x"ff4b3275",
			3155 => x"fd9d3275",
			3156 => x"01005110",
			3157 => x"05052d08",
			3158 => x"05051104",
			3159 => x"ffde3275",
			3160 => x"00ff3275",
			3161 => x"07048f04",
			3162 => x"fe003275",
			3163 => x"00223275",
			3164 => x"09008b08",
			3165 => x"07049704",
			3166 => x"00333275",
			3167 => x"ff6a3275",
			3168 => x"0e04a904",
			3169 => x"00553275",
			3170 => x"00003275",
			3171 => x"09008a04",
			3172 => x"fcdd3275",
			3173 => x"0b04e208",
			3174 => x"040c9a04",
			3175 => x"fef43275",
			3176 => x"01a43275",
			3177 => x"0900ba08",
			3178 => x"0e051d04",
			3179 => x"00003275",
			3180 => x"fd353275",
			3181 => x"0e05d804",
			3182 => x"016d3275",
			3183 => x"01008404",
			3184 => x"fe123275",
			3185 => x"fff73275",
			3186 => x"040d5514",
			3187 => x"040d0e10",
			3188 => x"0b04a204",
			3189 => x"01943275",
			3190 => x"0b04b904",
			3191 => x"fe2f3275",
			3192 => x"06016c04",
			3193 => x"01a43275",
			3194 => x"ff123275",
			3195 => x"01bf3275",
			3196 => x"0c047518",
			3197 => x"0b048e10",
			3198 => x"07047a04",
			3199 => x"fe893275",
			3200 => x"040eab04",
			3201 => x"01503275",
			3202 => x"0a034104",
			3203 => x"fed73275",
			3204 => x"00003275",
			3205 => x"0303b004",
			3206 => x"00c63275",
			3207 => x"fc8b3275",
			3208 => x"0704a814",
			3209 => x"040e6308",
			3210 => x"05051e04",
			3211 => x"02183275",
			3212 => x"00fe3275",
			3213 => x"06014608",
			3214 => x"0a031004",
			3215 => x"feb03275",
			3216 => x"00003275",
			3217 => x"00f83275",
			3218 => x"0c049408",
			3219 => x"0704bc04",
			3220 => x"fe0e3275",
			3221 => x"00403275",
			3222 => x"00055408",
			3223 => x"09008c04",
			3224 => x"01b13275",
			3225 => x"006b3275",
			3226 => x"0208fe04",
			3227 => x"00003275",
			3228 => x"feb63275",
			3229 => x"07058b64",
			3230 => x"040eab44",
			3231 => x"06010a04",
			3232 => x"fe5e33d9",
			3233 => x"0e048820",
			3234 => x"05054a10",
			3235 => x"03047708",
			3236 => x"09006204",
			3237 => x"00b133d9",
			3238 => x"018433d9",
			3239 => x"09006804",
			3240 => x"fe1033d9",
			3241 => x"00a633d9",
			3242 => x"0b04ce08",
			3243 => x"0f066604",
			3244 => x"004833d9",
			3245 => x"01f633d9",
			3246 => x"0704c104",
			3247 => x"002f33d9",
			3248 => x"01af33d9",
			3249 => x"02087e10",
			3250 => x"06012908",
			3251 => x"05056504",
			3252 => x"003833d9",
			3253 => x"01ee33d9",
			3254 => x"02080904",
			3255 => x"ff3d33d9",
			3256 => x"003d33d9",
			3257 => x"06014a08",
			3258 => x"0d053204",
			3259 => x"ff9b33d9",
			3260 => x"014833d9",
			3261 => x"040c6604",
			3262 => x"004033d9",
			3263 => x"00f333d9",
			3264 => x"020a861c",
			3265 => x"01005614",
			3266 => x"0e03b40c",
			3267 => x"01002504",
			3268 => x"fe5d33d9",
			3269 => x"040fc604",
			3270 => x"fe4833d9",
			3271 => x"00a033d9",
			3272 => x"01002d04",
			3273 => x"fea633d9",
			3274 => x"fcc933d9",
			3275 => x"0e04d304",
			3276 => x"00f533d9",
			3277 => x"fe6733d9",
			3278 => x"000033d9",
			3279 => x"08032614",
			3280 => x"0c054608",
			3281 => x"0c054304",
			3282 => x"fec433d9",
			3283 => x"022033d9",
			3284 => x"0e068d08",
			3285 => x"0506af04",
			3286 => x"fec833d9",
			3287 => x"02f933d9",
			3288 => x"fe5b33d9",
			3289 => x"040e6324",
			3290 => x"0803a020",
			3291 => x"0f0abc10",
			3292 => x"040caf08",
			3293 => x"0c059904",
			3294 => x"000033d9",
			3295 => x"028d33d9",
			3296 => x"09015c04",
			3297 => x"00f233d9",
			3298 => x"fe6833d9",
			3299 => x"0c06a108",
			3300 => x"08036b04",
			3301 => x"fe5d33d9",
			3302 => x"001333d9",
			3303 => x"0f0bae04",
			3304 => x"03af33d9",
			3305 => x"ff8133d9",
			3306 => x"023133d9",
			3307 => x"04110314",
			3308 => x"08044e0c",
			3309 => x"040fc608",
			3310 => x"040f7004",
			3311 => x"fe7733d9",
			3312 => x"003a33d9",
			3313 => x"fe6e33d9",
			3314 => x"08045904",
			3315 => x"012133d9",
			3316 => x"feb933d9",
			3317 => x"fe5d33d9",
			3318 => x"07056180",
			3319 => x"01003210",
			3320 => x"01002504",
			3321 => x"fe3b354d",
			3322 => x"0303bd04",
			3323 => x"0290354d",
			3324 => x"07047e04",
			3325 => x"fe39354d",
			3326 => x"007e354d",
			3327 => x"0e051d3c",
			3328 => x"00048a20",
			3329 => x"0304d810",
			3330 => x"09006208",
			3331 => x"03043e04",
			3332 => x"031c354d",
			3333 => x"fda5354d",
			3334 => x"040c7f04",
			3335 => x"0249354d",
			3336 => x"0078354d",
			3337 => x"09007508",
			3338 => x"0c047804",
			3339 => x"fdf2354d",
			3340 => x"fed1354d",
			3341 => x"02087e04",
			3342 => x"0156354d",
			3343 => x"0251354d",
			3344 => x"040eab10",
			3345 => x"07047d08",
			3346 => x"02081104",
			3347 => x"02b3354d",
			3348 => x"00e2354d",
			3349 => x"0803a304",
			3350 => x"0262354d",
			3351 => x"02dd354d",
			3352 => x"00057a04",
			3353 => x"fe8b354d",
			3354 => x"0f079104",
			3355 => x"024f354d",
			3356 => x"fe85354d",
			3357 => x"040bc418",
			3358 => x"0409b308",
			3359 => x"0c04cf04",
			3360 => x"ff1b354d",
			3361 => x"fe45354d",
			3362 => x"0c04ec08",
			3363 => x"0a024104",
			3364 => x"0222354d",
			3365 => x"fff4354d",
			3366 => x"07050404",
			3367 => x"0082354d",
			3368 => x"0275354d",
			3369 => x"0d061f10",
			3370 => x"0704be08",
			3371 => x"0f07a604",
			3372 => x"fec4354d",
			3373 => x"0147354d",
			3374 => x"07050504",
			3375 => x"01c3354d",
			3376 => x"02c9354d",
			3377 => x"00043104",
			3378 => x"02c0354d",
			3379 => x"01008204",
			3380 => x"0136354d",
			3381 => x"ff1e354d",
			3382 => x"07058b18",
			3383 => x"040d2e0c",
			3384 => x"0a027d04",
			3385 => x"fe4d354d",
			3386 => x"0c054804",
			3387 => x"00e8354d",
			3388 => x"0364354d",
			3389 => x"07057308",
			3390 => x"0e061e04",
			3391 => x"fe90354d",
			3392 => x"0192354d",
			3393 => x"fe46354d",
			3394 => x"08032604",
			3395 => x"fe3b354d",
			3396 => x"040eab1c",
			3397 => x"0803560c",
			3398 => x"09015c04",
			3399 => x"02b3354d",
			3400 => x"0c06de04",
			3401 => x"fe77354d",
			3402 => x"00dc354d",
			3403 => x"020c2a08",
			3404 => x"040c1804",
			3405 => x"fefb354d",
			3406 => x"0293354d",
			3407 => x"05094f04",
			3408 => x"fe83354d",
			3409 => x"01a8354d",
			3410 => x"fe3a354d",
			3411 => x"07057788",
			3412 => x"01003218",
			3413 => x"02074b08",
			3414 => x"0504e404",
			3415 => x"feaf36e9",
			3416 => x"013436e9",
			3417 => x"06014e08",
			3418 => x"02076704",
			3419 => x"ff5736e9",
			3420 => x"fe5736e9",
			3421 => x"0a03ae04",
			3422 => x"006736e9",
			3423 => x"fe8236e9",
			3424 => x"0e057140",
			3425 => x"0704be20",
			3426 => x"03051b10",
			3427 => x"07047808",
			3428 => x"02080704",
			3429 => x"007336e9",
			3430 => x"fe9836e9",
			3431 => x"03049f04",
			3432 => x"015136e9",
			3433 => x"00d536e9",
			3434 => x"02085908",
			3435 => x"09009104",
			3436 => x"fed036e9",
			3437 => x"fff836e9",
			3438 => x"09008604",
			3439 => x"ff5036e9",
			3440 => x"00b136e9",
			3441 => x"0d05ed10",
			3442 => x"0208bb08",
			3443 => x"06012b04",
			3444 => x"020236e9",
			3445 => x"00e136e9",
			3446 => x"08036104",
			3447 => x"02f136e9",
			3448 => x"016836e9",
			3449 => x"06015608",
			3450 => x"02076704",
			3451 => x"fe9b36e9",
			3452 => x"fd1c36e9",
			3453 => x"02093d04",
			3454 => x"01f536e9",
			3455 => x"fe8736e9",
			3456 => x"02089814",
			3457 => x"05061610",
			3458 => x"0704ee08",
			3459 => x"01008204",
			3460 => x"ff2836e9",
			3461 => x"013736e9",
			3462 => x"06015104",
			3463 => x"003f36e9",
			3464 => x"01f636e9",
			3465 => x"fe3036e9",
			3466 => x"06014a0c",
			3467 => x"06013d04",
			3468 => x"ff9136e9",
			3469 => x"08031d04",
			3470 => x"00df36e9",
			3471 => x"03be36e9",
			3472 => x"07050408",
			3473 => x"040c3804",
			3474 => x"ffa536e9",
			3475 => x"00a836e9",
			3476 => x"0d061d04",
			3477 => x"016f36e9",
			3478 => x"004636e9",
			3479 => x"0803260c",
			3480 => x"0100c308",
			3481 => x"0100bd04",
			3482 => x"fe7236e9",
			3483 => x"02b536e9",
			3484 => x"fe5936e9",
			3485 => x"040e632c",
			3486 => x"08037318",
			3487 => x"0e0ab80c",
			3488 => x"040d0008",
			3489 => x"040bb004",
			3490 => x"ff8436e9",
			3491 => x"024936e9",
			3492 => x"fe2336e9",
			3493 => x"0601be04",
			3494 => x"fe5036e9",
			3495 => x"0601c004",
			3496 => x"009236e9",
			3497 => x"fe5236e9",
			3498 => x"040d880c",
			3499 => x"020bbc08",
			3500 => x"020b3204",
			3501 => x"01d736e9",
			3502 => x"00b736e9",
			3503 => x"02bf36e9",
			3504 => x"08039c04",
			3505 => x"fe0c36e9",
			3506 => x"020836e9",
			3507 => x"0411030c",
			3508 => x"08044e04",
			3509 => x"fe8736e9",
			3510 => x"08045904",
			3511 => x"010036e9",
			3512 => x"fe9f36e9",
			3513 => x"fe5836e9",
			3514 => x"00038530",
			3515 => x"06012110",
			3516 => x"0f061a04",
			3517 => x"fe17389d",
			3518 => x"08026404",
			3519 => x"ff33389d",
			3520 => x"01004f04",
			3521 => x"0000389d",
			3522 => x"01aa389d",
			3523 => x"0802cc18",
			3524 => x"06012508",
			3525 => x"08023304",
			3526 => x"0000389d",
			3527 => x"fc5f389d",
			3528 => x"06012d0c",
			3529 => x"06012804",
			3530 => x"fe9e389d",
			3531 => x"06012904",
			3532 => x"000c389d",
			3533 => x"fffa389d",
			3534 => x"fe43389d",
			3535 => x"06016f04",
			3536 => x"014e389d",
			3537 => x"fee3389d",
			3538 => x"0900cd60",
			3539 => x"0704da28",
			3540 => x"0704d91c",
			3541 => x"0704d710",
			3542 => x"0704c408",
			3543 => x"0704c104",
			3544 => x"0005389d",
			3545 => x"00e3389d",
			3546 => x"0b04d004",
			3547 => x"fee9389d",
			3548 => x"ffd9389d",
			3549 => x"0c049304",
			3550 => x"fe89389d",
			3551 => x"0d057604",
			3552 => x"0288389d",
			3553 => x"007c389d",
			3554 => x"0e056808",
			3555 => x"06014904",
			3556 => x"01b3389d",
			3557 => x"027b389d",
			3558 => x"006e389d",
			3559 => x"0704eb1c",
			3560 => x"08034f0c",
			3561 => x"040baa08",
			3562 => x"00042104",
			3563 => x"002f389d",
			3564 => x"fe1c389d",
			3565 => x"01b4389d",
			3566 => x"03058908",
			3567 => x"03057704",
			3568 => x"ff18389d",
			3569 => x"01e0389d",
			3570 => x"01007304",
			3571 => x"fda7389d",
			3572 => x"ff8c389d",
			3573 => x"0f082b10",
			3574 => x"0900a408",
			3575 => x"0b052204",
			3576 => x"ff52389d",
			3577 => x"fc8f389d",
			3578 => x"0900a804",
			3579 => x"0206389d",
			3580 => x"0000389d",
			3581 => x"01007c08",
			3582 => x"07050504",
			3583 => x"fd9d389d",
			3584 => x"ff94389d",
			3585 => x"0000389d",
			3586 => x"0c04af0c",
			3587 => x"0c04ad08",
			3588 => x"0b052204",
			3589 => x"0216389d",
			3590 => x"fe40389d",
			3591 => x"02f4389d",
			3592 => x"0e05e020",
			3593 => x"0208db10",
			3594 => x"0e05bb08",
			3595 => x"08034c04",
			3596 => x"ff73389d",
			3597 => x"01ca389d",
			3598 => x"03062904",
			3599 => x"0310389d",
			3600 => x"016d389d",
			3601 => x"0e05bb08",
			3602 => x"0d062a04",
			3603 => x"01da389d",
			3604 => x"0000389d",
			3605 => x"06016704",
			3606 => x"fd89389d",
			3607 => x"0116389d",
			3608 => x"0f07d510",
			3609 => x"040a9508",
			3610 => x"0802f304",
			3611 => x"ff2a389d",
			3612 => x"0158389d",
			3613 => x"07050304",
			3614 => x"fe4e389d",
			3615 => x"fd1b389d",
			3616 => x"0704ec08",
			3617 => x"02092404",
			3618 => x"fdc8389d",
			3619 => x"0070389d",
			3620 => x"03068304",
			3621 => x"0114389d",
			3622 => x"000b389d",
			3623 => x"0505f978",
			3624 => x"0100361c",
			3625 => x"06013910",
			3626 => x"06013508",
			3627 => x"02071704",
			3628 => x"e5df3a91",
			3629 => x"e4df3a91",
			3630 => x"0504e204",
			3631 => x"e5033a91",
			3632 => x"e6e53a91",
			3633 => x"0303c504",
			3634 => x"ed513a91",
			3635 => x"02080704",
			3636 => x"e9933a91",
			3637 => x"e5033a91",
			3638 => x"03051b28",
			3639 => x"06010a08",
			3640 => x"05050204",
			3641 => x"e4f83a91",
			3642 => x"e5f83a91",
			3643 => x"03050010",
			3644 => x"07047a08",
			3645 => x"0c045404",
			3646 => x"e7b93a91",
			3647 => x"eba43a91",
			3648 => x"03048f04",
			3649 => x"edb43a91",
			3650 => x"ec873a91",
			3651 => x"0d054d08",
			3652 => x"0704a904",
			3653 => x"e8f93a91",
			3654 => x"ebe23a91",
			3655 => x"09008b04",
			3656 => x"ead93a91",
			3657 => x"ed373a91",
			3658 => x"00045418",
			3659 => x"06010e08",
			3660 => x"06010704",
			3661 => x"e4e33a91",
			3662 => x"e5a93a91",
			3663 => x"06013508",
			3664 => x"0704a604",
			3665 => x"e86b3a91",
			3666 => x"eb0f3a91",
			3667 => x"00041d04",
			3668 => x"e7503a91",
			3669 => x"e8ce3a91",
			3670 => x"06017010",
			3671 => x"00048208",
			3672 => x"0704aa04",
			3673 => x"e8f73a91",
			3674 => x"eb583a91",
			3675 => x"09008404",
			3676 => x"e9703a91",
			3677 => x"ecec3a91",
			3678 => x"07051808",
			3679 => x"0305b904",
			3680 => x"ea7d3a91",
			3681 => x"e54a3a91",
			3682 => x"e9ec3a91",
			3683 => x"07055d48",
			3684 => x"03065914",
			3685 => x"0c054510",
			3686 => x"0d062b08",
			3687 => x"03063204",
			3688 => x"e4e93a91",
			3689 => x"e9fe3a91",
			3690 => x"0c052e04",
			3691 => x"e4e83a91",
			3692 => x"e5f83a91",
			3693 => x"e89b3a91",
			3694 => x"06017718",
			3695 => x"00037d08",
			3696 => x"07052f04",
			3697 => x"e5f83a91",
			3698 => x"e4e83a91",
			3699 => x"08039008",
			3700 => x"07050804",
			3701 => x"e6303a91",
			3702 => x"ebbf3a91",
			3703 => x"00052904",
			3704 => x"e5f83a91",
			3705 => x"e5073a91",
			3706 => x"07054510",
			3707 => x"01009d08",
			3708 => x"00042504",
			3709 => x"e89b3a91",
			3710 => x"e5333a91",
			3711 => x"08036804",
			3712 => x"e4e23a91",
			3713 => x"e58b3a91",
			3714 => x"0209f704",
			3715 => x"ee423a91",
			3716 => x"0307c404",
			3717 => x"e4f53a91",
			3718 => x"e8463a91",
			3719 => x"09026b34",
			3720 => x"07057718",
			3721 => x"0f08d410",
			3722 => x"0d066a08",
			3723 => x"0f078e04",
			3724 => x"e4e73a91",
			3725 => x"ea7d3a91",
			3726 => x"03077c04",
			3727 => x"e4ed3a91",
			3728 => x"e5d03a91",
			3729 => x"0c052804",
			3730 => x"e4f73a91",
			3731 => x"ec243a91",
			3732 => x"0803260c",
			3733 => x"0c054608",
			3734 => x"0c054304",
			3735 => x"e4f23a91",
			3736 => x"e6293a91",
			3737 => x"e4df3a91",
			3738 => x"0004dd08",
			3739 => x"0100b404",
			3740 => x"ed993a91",
			3741 => x"e5673a91",
			3742 => x"0a02ed04",
			3743 => x"e5ca3a91",
			3744 => x"e4e03a91",
			3745 => x"00042904",
			3746 => x"e4fc3a91",
			3747 => x"e98c3a91",
			3748 => x"040eaba8",
			3749 => x"0100c374",
			3750 => x"01008040",
			3751 => x"0e057120",
			3752 => x"0900a810",
			3753 => x"03057908",
			3754 => x"09008f04",
			3755 => x"fffd3c15",
			3756 => x"004d3c15",
			3757 => x"0208d404",
			3758 => x"ff153c15",
			3759 => x"009a3c15",
			3760 => x"0207da08",
			3761 => x"0802d804",
			3762 => x"00923c15",
			3763 => x"fe1d3c15",
			3764 => x"0a025e04",
			3765 => x"018f3c15",
			3766 => x"006f3c15",
			3767 => x"0b04c310",
			3768 => x"0704a608",
			3769 => x"0d055904",
			3770 => x"010e3c15",
			3771 => x"fe333c15",
			3772 => x"06014904",
			3773 => x"03b73c15",
			3774 => x"00953c15",
			3775 => x"01006708",
			3776 => x"0f080504",
			3777 => x"fd6c3c15",
			3778 => x"00da3c15",
			3779 => x"0208c704",
			3780 => x"ff8a3c15",
			3781 => x"000d3c15",
			3782 => x"0e05e018",
			3783 => x"0803360c",
			3784 => x"0704f104",
			3785 => x"01c43c15",
			3786 => x"0e057f04",
			3787 => x"00fe3c15",
			3788 => x"fe733c15",
			3789 => x"0b052204",
			3790 => x"00283c15",
			3791 => x"06015b04",
			3792 => x"02993c15",
			3793 => x"01ac3c15",
			3794 => x"07051810",
			3795 => x"01009208",
			3796 => x"0c04ae04",
			3797 => x"01f93c15",
			3798 => x"ffcd3c15",
			3799 => x"040ac904",
			3800 => x"ffda3c15",
			3801 => x"fe1b3c15",
			3802 => x"0802ae04",
			3803 => x"fe803c15",
			3804 => x"0d06b904",
			3805 => x"00853c15",
			3806 => x"01e93c15",
			3807 => x"08034714",
			3808 => x"0c06de10",
			3809 => x"040b8304",
			3810 => x"fe613c15",
			3811 => x"040b8508",
			3812 => x"08030104",
			3813 => x"00003c15",
			3814 => x"00f43c15",
			3815 => x"feb83c15",
			3816 => x"007c3c15",
			3817 => x"0b061b04",
			3818 => x"fe6a3c15",
			3819 => x"0601bb10",
			3820 => x"040cf508",
			3821 => x"0a02bb04",
			3822 => x"016d3c15",
			3823 => x"ffbb3c15",
			3824 => x"0a02e104",
			3825 => x"fe873c15",
			3826 => x"01123c15",
			3827 => x"0e0c7e08",
			3828 => x"040c2604",
			3829 => x"ff703c15",
			3830 => x"014d3c15",
			3831 => x"ffef3c15",
			3832 => x"06016704",
			3833 => x"fe5e3c15",
			3834 => x"02091108",
			3835 => x"01001604",
			3836 => x"ffe73c15",
			3837 => x"017f3c15",
			3838 => x"0a03150c",
			3839 => x"0803e604",
			3840 => x"fec83c15",
			3841 => x"04112a04",
			3842 => x"01c63c15",
			3843 => x"00003c15",
			3844 => x"fe993c15",
			3845 => x"0c057f90",
			3846 => x"040eab78",
			3847 => x"0e04e23c",
			3848 => x"0900951c",
			3849 => x"0b04d210",
			3850 => x"0d054d08",
			3851 => x"03050004",
			3852 => x"004d3d99",
			3853 => x"ff823d99",
			3854 => x"02086804",
			3855 => x"00493d99",
			3856 => x"01623d99",
			3857 => x"0a02bc08",
			3858 => x"02084504",
			3859 => x"ff063d99",
			3860 => x"fce03d99",
			3861 => x"01aa3d99",
			3862 => x"01005c10",
			3863 => x"0e04bb08",
			3864 => x"05053d04",
			3865 => x"00693d99",
			3866 => x"02813d99",
			3867 => x"0f073304",
			3868 => x"fffc3d99",
			3869 => x"02a53d99",
			3870 => x"09009b08",
			3871 => x"0b04c004",
			3872 => x"ff013d99",
			3873 => x"00753d99",
			3874 => x"0f06d604",
			3875 => x"00253d99",
			3876 => x"011f3d99",
			3877 => x"0f07051c",
			3878 => x"0900aa10",
			3879 => x"0b04af08",
			3880 => x"0c047504",
			3881 => x"034b3d99",
			3882 => x"ffd23d99",
			3883 => x"0802e804",
			3884 => x"fec63d99",
			3885 => x"fdaa3d99",
			3886 => x"05057604",
			3887 => x"fdc43d99",
			3888 => x"0e053404",
			3889 => x"00d63d99",
			3890 => x"feb73d99",
			3891 => x"0900af10",
			3892 => x"0208d008",
			3893 => x"0e053b04",
			3894 => x"ffe73d99",
			3895 => x"fee33d99",
			3896 => x"0505af04",
			3897 => x"00c13d99",
			3898 => x"fe0a3d99",
			3899 => x"0e057808",
			3900 => x"0d057404",
			3901 => x"fe4b3d99",
			3902 => x"00d83d99",
			3903 => x"0900cd04",
			3904 => x"ffb73d99",
			3905 => x"00563d99",
			3906 => x"0b05f914",
			3907 => x"01002504",
			3908 => x"fe683d99",
			3909 => x"0f062f04",
			3910 => x"00363d99",
			3911 => x"02088304",
			3912 => x"fd743d99",
			3913 => x"0208f004",
			3914 => x"01153d99",
			3915 => x"fe283d99",
			3916 => x"01b83d99",
			3917 => x"08032608",
			3918 => x"0e068d04",
			3919 => x"01673d99",
			3920 => x"fe633d99",
			3921 => x"040fc628",
			3922 => x"0e0a1b14",
			3923 => x"020aaf0c",
			3924 => x"09016708",
			3925 => x"040d8804",
			3926 => x"01a83d99",
			3927 => x"00003d99",
			3928 => x"feb43d99",
			3929 => x"020b1f04",
			3930 => x"027e3d99",
			3931 => x"00953d99",
			3932 => x"0c06dc0c",
			3933 => x"08034c04",
			3934 => x"fe6d3d99",
			3935 => x"00044304",
			3936 => x"01073d99",
			3937 => x"fef33d99",
			3938 => x"01014b04",
			3939 => x"fea53d99",
			3940 => x"02403d99",
			3941 => x"fe663d99",
			3942 => x"0505f6ac",
			3943 => x"0a027b5c",
			3944 => x"0b048e1c",
			3945 => x"0003e608",
			3946 => x"0e046104",
			3947 => x"fca93f7d",
			3948 => x"fead3f7d",
			3949 => x"040b3c04",
			3950 => x"01573f7d",
			3951 => x"0e042e08",
			3952 => x"0a026204",
			3953 => x"fd1c3f7d",
			3954 => x"00723f7d",
			3955 => x"08031e04",
			3956 => x"fac73f7d",
			3957 => x"fe1a3f7d",
			3958 => x"02085b20",
			3959 => x"040b3610",
			3960 => x"0e045308",
			3961 => x"040b2204",
			3962 => x"01b03f7d",
			3963 => x"ff993f7d",
			3964 => x"09008704",
			3965 => x"fddc3f7d",
			3966 => x"002a3f7d",
			3967 => x"0f06e508",
			3968 => x"02082a04",
			3969 => x"007f3f7d",
			3970 => x"fd703f7d",
			3971 => x"02082404",
			3972 => x"006f3f7d",
			3973 => x"01aa3f7d",
			3974 => x"08031d10",
			3975 => x"0a026d08",
			3976 => x"040acf04",
			3977 => x"ffda3f7d",
			3978 => x"01eb3f7d",
			3979 => x"0208a404",
			3980 => x"fee23f7d",
			3981 => x"02073f7d",
			3982 => x"06013608",
			3983 => x"05054a04",
			3984 => x"02a73f7d",
			3985 => x"ffa63f7d",
			3986 => x"0704c404",
			3987 => x"04133f7d",
			3988 => x"013c3f7d",
			3989 => x"040b9f18",
			3990 => x"00045210",
			3991 => x"0003ed04",
			3992 => x"02ff3f7d",
			3993 => x"01004904",
			3994 => x"01f93f7d",
			3995 => x"0505bd04",
			3996 => x"ff633f7d",
			3997 => x"00613f7d",
			3998 => x"02087604",
			3999 => x"03f53f7d",
			4000 => x"017d3f7d",
			4001 => x"06012b18",
			4002 => x"0704a610",
			4003 => x"07049208",
			4004 => x"08034104",
			4005 => x"018b3f7d",
			4006 => x"fe753f7d",
			4007 => x"0f063b04",
			4008 => x"00013f7d",
			4009 => x"fbcd3f7d",
			4010 => x"05051004",
			4011 => x"fd3b3f7d",
			4012 => x"01cb3f7d",
			4013 => x"0a029e10",
			4014 => x"0900a808",
			4015 => x"0e04bb04",
			4016 => x"00973f7d",
			4017 => x"ffe63f7d",
			4018 => x"0c04ed04",
			4019 => x"01513f7d",
			4020 => x"fef63f7d",
			4021 => x"040c1808",
			4022 => x"0900c604",
			4023 => x"ff3d3f7d",
			4024 => x"00d73f7d",
			4025 => x"0c047204",
			4026 => x"ff9e3f7d",
			4027 => x"00503f7d",
			4028 => x"0802eb18",
			4029 => x"05061614",
			4030 => x"07051a0c",
			4031 => x"06013908",
			4032 => x"0c04ed04",
			4033 => x"00e43f7d",
			4034 => x"00003f7d",
			4035 => x"fe0b3f7d",
			4036 => x"0f05da04",
			4037 => x"ff593f7d",
			4038 => x"02543f7d",
			4039 => x"fe613f7d",
			4040 => x"0411032c",
			4041 => x"0b054310",
			4042 => x"00040204",
			4043 => x"01123f7d",
			4044 => x"0900d304",
			4045 => x"fcbe3f7d",
			4046 => x"02093004",
			4047 => x"ff3b3f7d",
			4048 => x"fdeb3f7d",
			4049 => x"0e0a390c",
			4050 => x"0802ee04",
			4051 => x"038a3f7d",
			4052 => x"0a030804",
			4053 => x"ffe93f7d",
			4054 => x"01f43f7d",
			4055 => x"0601b708",
			4056 => x"0c06e304",
			4057 => x"fe673f7d",
			4058 => x"009d3f7d",
			4059 => x"0f0c3904",
			4060 => x"00cf3f7d",
			4061 => x"ff393f7d",
			4062 => x"fe693f7d",
			4063 => x"09007b88",
			4064 => x"05051d44",
			4065 => x"0505143c",
			4066 => x"02082a1c",
			4067 => x"0304b710",
			4068 => x"040c4c08",
			4069 => x"08031404",
			4070 => x"fe0941a9",
			4071 => x"005d41a9",
			4072 => x"0a02a504",
			4073 => x"fe3941a9",
			4074 => x"ffbc41a9",
			4075 => x"08033708",
			4076 => x"0304d604",
			4077 => x"010941a9",
			4078 => x"fdfb41a9",
			4079 => x"fdd741a9",
			4080 => x"0a02ac10",
			4081 => x"0a02a608",
			4082 => x"0d050204",
			4083 => x"fe4c41a9",
			4084 => x"00b141a9",
			4085 => x"07046604",
			4086 => x"ffdf41a9",
			4087 => x"021741a9",
			4088 => x"06013e08",
			4089 => x"02088904",
			4090 => x"ffae41a9",
			4091 => x"fdbb41a9",
			4092 => x"02088504",
			4093 => x"003441a9",
			4094 => x"01a141a9",
			4095 => x"040d0004",
			4096 => x"01c941a9",
			4097 => x"ffdd41a9",
			4098 => x"06013424",
			4099 => x"0d051b0c",
			4100 => x"0c049308",
			4101 => x"040bfa04",
			4102 => x"fe9941a9",
			4103 => x"018f41a9",
			4104 => x"fd3941a9",
			4105 => x"0004320c",
			4106 => x"0304be04",
			4107 => x"018641a9",
			4108 => x"0207df04",
			4109 => x"fdf041a9",
			4110 => x"000041a9",
			4111 => x"0208b908",
			4112 => x"09005d04",
			4113 => x"000041a9",
			4114 => x"01d441a9",
			4115 => x"ffc741a9",
			4116 => x"0e043614",
			4117 => x"0e041e10",
			4118 => x"0b049108",
			4119 => x"03048f04",
			4120 => x"ffea41a9",
			4121 => x"fd8b41a9",
			4122 => x"06013604",
			4123 => x"017941a9",
			4124 => x"ff6841a9",
			4125 => x"00e841a9",
			4126 => x"0e048508",
			4127 => x"02088304",
			4128 => x"fe7141a9",
			4129 => x"fd1741a9",
			4130 => x"fff741a9",
			4131 => x"0305334c",
			4132 => x"03052f34",
			4133 => x"03052b20",
			4134 => x"03052710",
			4135 => x"03052508",
			4136 => x"0d057504",
			4137 => x"002041a9",
			4138 => x"01e241a9",
			4139 => x"0c047404",
			4140 => x"017841a9",
			4141 => x"fec741a9",
			4142 => x"0a02b308",
			4143 => x"05053d04",
			4144 => x"008e41a9",
			4145 => x"022641a9",
			4146 => x"08038504",
			4147 => x"fdbd41a9",
			4148 => x"018741a9",
			4149 => x"0a027f08",
			4150 => x"0d054e04",
			4151 => x"016b41a9",
			4152 => x"ff1c41a9",
			4153 => x"02088b08",
			4154 => x"0d056604",
			4155 => x"fe0a41a9",
			4156 => x"ff4541a9",
			4157 => x"ffe541a9",
			4158 => x"0b04c20c",
			4159 => x"0704a504",
			4160 => x"00eb41a9",
			4161 => x"0e04a504",
			4162 => x"011a41a9",
			4163 => x"026241a9",
			4164 => x"09009a04",
			4165 => x"ffa841a9",
			4166 => x"0704c404",
			4167 => x"006141a9",
			4168 => x"01c041a9",
			4169 => x"0d05350c",
			4170 => x"0e050008",
			4171 => x"02088904",
			4172 => x"ff5a41a9",
			4173 => x"fd6a41a9",
			4174 => x"00ba41a9",
			4175 => x"03053f1c",
			4176 => x"03053910",
			4177 => x"0a027a08",
			4178 => x"0b04be04",
			4179 => x"fecc41a9",
			4180 => x"01b141a9",
			4181 => x"00045204",
			4182 => x"fe8441a9",
			4183 => x"002441a9",
			4184 => x"0d057408",
			4185 => x"02085904",
			4186 => x"fec741a9",
			4187 => x"fdce41a9",
			4188 => x"00b341a9",
			4189 => x"0305430c",
			4190 => x"0a02bb08",
			4191 => x"02082f04",
			4192 => x"00bf41a9",
			4193 => x"024341a9",
			4194 => x"fe9b41a9",
			4195 => x"0c04b108",
			4196 => x"0c04af04",
			4197 => x"ffea41a9",
			4198 => x"ff5241a9",
			4199 => x"0704c304",
			4200 => x"005f41a9",
			4201 => x"fffb41a9",
			4202 => x"0304d88c",
			4203 => x"040c8c44",
			4204 => x"00048a34",
			4205 => x"0304cf20",
			4206 => x"0304c710",
			4207 => x"06014108",
			4208 => x"0e041e04",
			4209 => x"001b43cd",
			4210 => x"00d943cd",
			4211 => x"09007b04",
			4212 => x"fe5043cd",
			4213 => x"ffec43cd",
			4214 => x"040be908",
			4215 => x"0704a804",
			4216 => x"fd4543cd",
			4217 => x"008543cd",
			4218 => x"0e042604",
			4219 => x"001b43cd",
			4220 => x"01c943cd",
			4221 => x"0b04910c",
			4222 => x"040bd804",
			4223 => x"01ad43cd",
			4224 => x"040c4704",
			4225 => x"fec043cd",
			4226 => x"003843cd",
			4227 => x"09008a04",
			4228 => x"01eb43cd",
			4229 => x"000043cd",
			4230 => x"06014504",
			4231 => x"01c843cd",
			4232 => x"0d051b04",
			4233 => x"fec243cd",
			4234 => x"0d054e04",
			4235 => x"017343cd",
			4236 => x"000043cd",
			4237 => x"040ca718",
			4238 => x"01005114",
			4239 => x"06013904",
			4240 => x"fd6043cd",
			4241 => x"0304b708",
			4242 => x"0b048e04",
			4243 => x"ff2343cd",
			4244 => x"00d043cd",
			4245 => x"06014204",
			4246 => x"ff9943cd",
			4247 => x"fcf943cd",
			4248 => x"017743cd",
			4249 => x"01003f1c",
			4250 => x"0f05ee0c",
			4251 => x"040eab04",
			4252 => x"016843cd",
			4253 => x"06017004",
			4254 => x"ff0d43cd",
			4255 => x"000043cd",
			4256 => x"0b047008",
			4257 => x"0504f204",
			4258 => x"ff4543cd",
			4259 => x"015c43cd",
			4260 => x"0c049304",
			4261 => x"fe0943cd",
			4262 => x"00cb43cd",
			4263 => x"01004308",
			4264 => x"0004f704",
			4265 => x"01c243cd",
			4266 => x"ff5843cd",
			4267 => x"0b047d04",
			4268 => x"fdfa43cd",
			4269 => x"0f06d004",
			4270 => x"ffe843cd",
			4271 => x"017a43cd",
			4272 => x"0900771c",
			4273 => x"06012b0c",
			4274 => x"0e045308",
			4275 => x"040d8804",
			4276 => x"01d043cd",
			4277 => x"000043cd",
			4278 => x"000043cd",
			4279 => x"06013904",
			4280 => x"fd8743cd",
			4281 => x"0e045a08",
			4282 => x"0f06ed04",
			4283 => x"023843cd",
			4284 => x"ffb243cd",
			4285 => x"fe9143cd",
			4286 => x"0f06c130",
			4287 => x"09008814",
			4288 => x"01005310",
			4289 => x"0e045308",
			4290 => x"07049704",
			4291 => x"001343cd",
			4292 => x"01cf43cd",
			4293 => x"05053c04",
			4294 => x"fe7543cd",
			4295 => x"009c43cd",
			4296 => x"fd6043cd",
			4297 => x"0d056710",
			4298 => x"0f06bb08",
			4299 => x"08031e04",
			4300 => x"016243cd",
			4301 => x"000443cd",
			4302 => x"03050d04",
			4303 => x"fe3043cd",
			4304 => x"ffaf43cd",
			4305 => x"0e045304",
			4306 => x"fda843cd",
			4307 => x"040bde04",
			4308 => x"ff1f43cd",
			4309 => x"012743cd",
			4310 => x"08034220",
			4311 => x"040ba410",
			4312 => x"0e047808",
			4313 => x"0d054104",
			4314 => x"fdfa43cd",
			4315 => x"00bb43cd",
			4316 => x"05057604",
			4317 => x"004343cd",
			4318 => x"ffdf43cd",
			4319 => x"0f074908",
			4320 => x"08032604",
			4321 => x"021543cd",
			4322 => x"000c43cd",
			4323 => x"0d058e04",
			4324 => x"020c43cd",
			4325 => x"009443cd",
			4326 => x"07047c0c",
			4327 => x"05052d08",
			4328 => x"05051d04",
			4329 => x"007243cd",
			4330 => x"025e43cd",
			4331 => x"ff2043cd",
			4332 => x"00048608",
			4333 => x"08036904",
			4334 => x"ffee43cd",
			4335 => x"ff9543cd",
			4336 => x"040c3804",
			4337 => x"01d643cd",
			4338 => x"000c43cd",
			4339 => x"0207a170",
			4340 => x"02076724",
			4341 => x"0003c410",
			4342 => x"0b049e04",
			4343 => x"fddb4621",
			4344 => x"0c049808",
			4345 => x"00034b04",
			4346 => x"ffd74621",
			4347 => x"01484621",
			4348 => x"fe714621",
			4349 => x"0c045c10",
			4350 => x"07047908",
			4351 => x"07046304",
			4352 => x"001e4621",
			4353 => x"fecc4621",
			4354 => x"01001f04",
			4355 => x"00004621",
			4356 => x"010e4621",
			4357 => x"01b64621",
			4358 => x"0b048e28",
			4359 => x"07047a1c",
			4360 => x"0704670c",
			4361 => x"06012b04",
			4362 => x"00004621",
			4363 => x"0a030d04",
			4364 => x"01554621",
			4365 => x"00004621",
			4366 => x"0c045908",
			4367 => x"02079804",
			4368 => x"00004621",
			4369 => x"00224621",
			4370 => x"06012904",
			4371 => x"00004621",
			4372 => x"fd334621",
			4373 => x"0f064208",
			4374 => x"01002d04",
			4375 => x"00004621",
			4376 => x"01a74621",
			4377 => x"ffd94621",
			4378 => x"05052c10",
			4379 => x"02077704",
			4380 => x"001f4621",
			4381 => x"0c049308",
			4382 => x"00046c04",
			4383 => x"fdeb4621",
			4384 => x"fc704621",
			4385 => x"ff064621",
			4386 => x"00043d10",
			4387 => x"06012108",
			4388 => x"0f068104",
			4389 => x"01794621",
			4390 => x"ffa64621",
			4391 => x"09008c04",
			4392 => x"fd374621",
			4393 => x"ff4e4621",
			4394 => x"01a14621",
			4395 => x"00040758",
			4396 => x"040b4634",
			4397 => x"0a028a20",
			4398 => x"0a026f10",
			4399 => x"08031808",
			4400 => x"040b3c04",
			4401 => x"00354621",
			4402 => x"fe2d4621",
			4403 => x"0b04c004",
			4404 => x"02774621",
			4405 => x"006f4621",
			4406 => x"040af508",
			4407 => x"01006f04",
			4408 => x"02a14621",
			4409 => x"00084621",
			4410 => x"0c04ce04",
			4411 => x"fe6e4621",
			4412 => x"00004621",
			4413 => x"0505f908",
			4414 => x"01008204",
			4415 => x"00be4621",
			4416 => x"026e4621",
			4417 => x"07051a04",
			4418 => x"fe784621",
			4419 => x"08032e04",
			4420 => x"fee94621",
			4421 => x"016e4621",
			4422 => x"01004904",
			4423 => x"fd6b4621",
			4424 => x"0003f110",
			4425 => x"08032608",
			4426 => x"0003ee04",
			4427 => x"ffc44621",
			4428 => x"fbdd4621",
			4429 => x"0c063a04",
			4430 => x"00004621",
			4431 => x"01894621",
			4432 => x"0c04cc08",
			4433 => x"0b04e004",
			4434 => x"00f34621",
			4435 => x"02a24621",
			4436 => x"08032304",
			4437 => x"013c4621",
			4438 => x"fed84621",
			4439 => x"0304b738",
			4440 => x"040c3218",
			4441 => x"0b049d10",
			4442 => x"07049208",
			4443 => x"06012b04",
			4444 => x"ff8d4621",
			4445 => x"01594621",
			4446 => x"040bbf04",
			4447 => x"01c64621",
			4448 => x"ff284621",
			4449 => x"0b04ae04",
			4450 => x"01de4621",
			4451 => x"004f4621",
			4452 => x"00048510",
			4453 => x"0c045b08",
			4454 => x"0b047f04",
			4455 => x"fe854621",
			4456 => x"01be4621",
			4457 => x"06012d04",
			4458 => x"fffc4621",
			4459 => x"fe2c4621",
			4460 => x"0c047608",
			4461 => x"0c047404",
			4462 => x"00754621",
			4463 => x"fe8e4621",
			4464 => x"0c047904",
			4465 => x"01854621",
			4466 => x"002f4621",
			4467 => x"08031d18",
			4468 => x"03056f0c",
			4469 => x"0c04ad08",
			4470 => x"0b04a004",
			4471 => x"00b14621",
			4472 => x"fee44621",
			4473 => x"01fa4621",
			4474 => x"0305f908",
			4475 => x"00040b04",
			4476 => x"fe9a4621",
			4477 => x"fd754621",
			4478 => x"00a74621",
			4479 => x"08031e04",
			4480 => x"01ad4621",
			4481 => x"0c047308",
			4482 => x"0c045c04",
			4483 => x"ffed4621",
			4484 => x"ff1d4621",
			4485 => x"0c047404",
			4486 => x"009c4621",
			4487 => x"ffff4621",
			4488 => x"07049090",
			4489 => x"0304af38",
			4490 => x"08031410",
			4491 => x"0207aa08",
			4492 => x"0c047304",
			4493 => x"fe0148ad",
			4494 => x"017d48ad",
			4495 => x"0e03da04",
			4496 => x"000048ad",
			4497 => x"fb6b48ad",
			4498 => x"040c3810",
			4499 => x"0601390c",
			4500 => x"0c045704",
			4501 => x"00a748ad",
			4502 => x"01003f04",
			4503 => x"00e648ad",
			4504 => x"01d648ad",
			4505 => x"006648ad",
			4506 => x"00046c08",
			4507 => x"03046704",
			4508 => x"000048ad",
			4509 => x"fcd948ad",
			4510 => x"09007108",
			4511 => x"0207cf04",
			4512 => x"013a48ad",
			4513 => x"ff9a48ad",
			4514 => x"0e03da04",
			4515 => x"ff2748ad",
			4516 => x"01a248ad",
			4517 => x"0c047628",
			4518 => x"0c045610",
			4519 => x"040c850c",
			4520 => x"03051708",
			4521 => x"07047904",
			4522 => x"00cf48ad",
			4523 => x"029548ad",
			4524 => x"fe5e48ad",
			4525 => x"fdaa48ad",
			4526 => x"0207df08",
			4527 => x"08032904",
			4528 => x"ff2548ad",
			4529 => x"fc5f48ad",
			4530 => x"0a028d08",
			4531 => x"00040b04",
			4532 => x"fdec48ad",
			4533 => x"001748ad",
			4534 => x"08036104",
			4535 => x"fdaa48ad",
			4536 => x"ff2948ad",
			4537 => x"07047d18",
			4538 => x"0304c708",
			4539 => x"02082a04",
			4540 => x"01df48ad",
			4541 => x"ffd948ad",
			4542 => x"0f073b08",
			4543 => x"0c049004",
			4544 => x"fcbe48ad",
			4545 => x"feff48ad",
			4546 => x"0208b404",
			4547 => x"024348ad",
			4548 => x"ffa248ad",
			4549 => x"0e04680c",
			4550 => x"0f06b504",
			4551 => x"002548ad",
			4552 => x"0304d804",
			4553 => x"013c48ad",
			4554 => x"026548ad",
			4555 => x"07048004",
			4556 => x"017c48ad",
			4557 => x"0d056604",
			4558 => x"ff0048ad",
			4559 => x"00dd48ad",
			4560 => x"0704ad4c",
			4561 => x"0704ac38",
			4562 => x"0f065f1c",
			4563 => x"0a025c0c",
			4564 => x"06011004",
			4565 => x"fe1448ad",
			4566 => x"0c049604",
			4567 => x"01ed48ad",
			4568 => x"000048ad",
			4569 => x"0e03f108",
			4570 => x"0d052804",
			4571 => x"ff5a48ad",
			4572 => x"013348ad",
			4573 => x"0f064a04",
			4574 => x"fbe548ad",
			4575 => x"fe9e48ad",
			4576 => x"0c04b410",
			4577 => x"0704a808",
			4578 => x"07049704",
			4579 => x"006b48ad",
			4580 => x"ffa848ad",
			4581 => x"0a02c904",
			4582 => x"00a448ad",
			4583 => x"fe9b48ad",
			4584 => x"01005c04",
			4585 => x"000148ad",
			4586 => x"0900a204",
			4587 => x"fd5348ad",
			4588 => x"ff0548ad",
			4589 => x"09009d10",
			4590 => x"0d055b08",
			4591 => x"0c049904",
			4592 => x"022c48ad",
			4593 => x"005048ad",
			4594 => x"03052704",
			4595 => x"ffb148ad",
			4596 => x"012248ad",
			4597 => x"02d248ad",
			4598 => x"0704be30",
			4599 => x"0a02bc1c",
			4600 => x"00046b10",
			4601 => x"09008f08",
			4602 => x"01005504",
			4603 => x"ff9848ad",
			4604 => x"fd1548ad",
			4605 => x"0a029e04",
			4606 => x"ffbc48ad",
			4607 => x"fe9448ad",
			4608 => x"0d057408",
			4609 => x"0d054c04",
			4610 => x"ff8248ad",
			4611 => x"018448ad",
			4612 => x"ff2648ad",
			4613 => x"0a02c308",
			4614 => x"08038804",
			4615 => x"fc0848ad",
			4616 => x"fe9648ad",
			4617 => x"0c049708",
			4618 => x"0c049104",
			4619 => x"002448ad",
			4620 => x"fd8248ad",
			4621 => x"00c948ad",
			4622 => x"0704c420",
			4623 => x"0704c110",
			4624 => x"0208ab08",
			4625 => x"0704bf04",
			4626 => x"00d048ad",
			4627 => x"ff8f48ad",
			4628 => x"06015204",
			4629 => x"020648ad",
			4630 => x"003f48ad",
			4631 => x"040b3c08",
			4632 => x"08031a04",
			4633 => x"018248ad",
			4634 => x"040f48ad",
			4635 => x"00042804",
			4636 => x"ffe248ad",
			4637 => x"011548ad",
			4638 => x"0704d40c",
			4639 => x"040cbf08",
			4640 => x"0a02c404",
			4641 => x"ff2b48ad",
			4642 => x"fc6648ad",
			4643 => x"018148ad",
			4644 => x"0900b708",
			4645 => x"0e055a04",
			4646 => x"fff848ad",
			4647 => x"ff0348ad",
			4648 => x"0704da04",
			4649 => x"010c48ad",
			4650 => x"001548ad",
			4651 => x"04095904",
			4652 => x"fe314a11",
			4653 => x"0704aa58",
			4654 => x"07049730",
			4655 => x"07049310",
			4656 => x"0100620c",
			4657 => x"09009e08",
			4658 => x"05055904",
			4659 => x"ffe44a11",
			4660 => x"02aa4a11",
			4661 => x"02674a11",
			4662 => x"fe294a11",
			4663 => x"0b049110",
			4664 => x"0f05e008",
			4665 => x"0c047804",
			4666 => x"00004a11",
			4667 => x"fce64a11",
			4668 => x"0b048e04",
			4669 => x"00a04a11",
			4670 => x"01df4a11",
			4671 => x"0b049e08",
			4672 => x"0c047904",
			4673 => x"fd724a11",
			4674 => x"ff8e4a11",
			4675 => x"0f072b04",
			4676 => x"00374a11",
			4677 => x"01a94a11",
			4678 => x"05051414",
			4679 => x"040c0408",
			4680 => x"0704a704",
			4681 => x"fe844a11",
			4682 => x"01ad4a11",
			4683 => x"02084408",
			4684 => x"0304a704",
			4685 => x"fe474a11",
			4686 => x"fbed4a11",
			4687 => x"00454a11",
			4688 => x"02090c10",
			4689 => x"040c9308",
			4690 => x"01006b04",
			4691 => x"ffa34a11",
			4692 => x"01364a11",
			4693 => x"0d053f04",
			4694 => x"fffc4a11",
			4695 => x"01364a11",
			4696 => x"fd184a11",
			4697 => x"0704ab18",
			4698 => x"06012404",
			4699 => x"fe844a11",
			4700 => x"05056610",
			4701 => x"05054808",
			4702 => x"0c049704",
			4703 => x"01434a11",
			4704 => x"ff494a11",
			4705 => x"06013504",
			4706 => x"00c44a11",
			4707 => x"02624a11",
			4708 => x"00174a11",
			4709 => x"0a024720",
			4710 => x"0c04d410",
			4711 => x"0305b008",
			4712 => x"03058704",
			4713 => x"010c4a11",
			4714 => x"feb84a11",
			4715 => x"06013604",
			4716 => x"01e44a11",
			4717 => x"00004a11",
			4718 => x"040a6908",
			4719 => x"040a0104",
			4720 => x"ff454a11",
			4721 => x"fe314a11",
			4722 => x"02094304",
			4723 => x"01954a11",
			4724 => x"ffab4a11",
			4725 => x"040c6610",
			4726 => x"0c047308",
			4727 => x"040b8304",
			4728 => x"005f4a11",
			4729 => x"02484a11",
			4730 => x"0900b904",
			4731 => x"ffd84a11",
			4732 => x"00194a11",
			4733 => x"08035b08",
			4734 => x"040c9a04",
			4735 => x"fbe14a11",
			4736 => x"ff184a11",
			4737 => x"08038504",
			4738 => x"00de4a11",
			4739 => x"fff04a11",
			4740 => x"09008fb0",
			4741 => x"03050d4c",
			4742 => x"0f06ed24",
			4743 => x"03050720",
			4744 => x"0e042610",
			4745 => x"0c049508",
			4746 => x"0c045904",
			4747 => x"00964ca5",
			4748 => x"ffd84ca5",
			4749 => x"03049704",
			4750 => x"00454ca5",
			4751 => x"017c4ca5",
			4752 => x"06013e08",
			4753 => x"09008204",
			4754 => x"ff7a4ca5",
			4755 => x"003f4ca5",
			4756 => x"06014504",
			4757 => x"fe974ca5",
			4758 => x"ffc54ca5",
			4759 => x"014b4ca5",
			4760 => x"09008018",
			4761 => x"0704930c",
			4762 => x"05052008",
			4763 => x"0304fe04",
			4764 => x"00884ca5",
			4765 => x"ff164ca5",
			4766 => x"fe814ca5",
			4767 => x"08034f04",
			4768 => x"ff704ca5",
			4769 => x"00067104",
			4770 => x"01dc4ca5",
			4771 => x"00004ca5",
			4772 => x"040bde04",
			4773 => x"ffce4ca5",
			4774 => x"09008d08",
			4775 => x"0704bd04",
			4776 => x"01fd4ca5",
			4777 => x"00984ca5",
			4778 => x"007d4ca5",
			4779 => x"02085228",
			4780 => x"05053b10",
			4781 => x"0d052604",
			4782 => x"00a44ca5",
			4783 => x"0207c504",
			4784 => x"02164ca5",
			4785 => x"09007f04",
			4786 => x"002c4ca5",
			4787 => x"fdf14ca5",
			4788 => x"05053c08",
			4789 => x"0f06de04",
			4790 => x"01ba4ca5",
			4791 => x"00604ca5",
			4792 => x"00043f08",
			4793 => x"040b2204",
			4794 => x"fe234ca5",
			4795 => x"003d4ca5",
			4796 => x"0c049204",
			4797 => x"ff914ca5",
			4798 => x"fdd94ca5",
			4799 => x"040c0c1c",
			4800 => x"0305390c",
			4801 => x"05053b08",
			4802 => x"00045b04",
			4803 => x"00184ca5",
			4804 => x"02144ca5",
			4805 => x"02714ca5",
			4806 => x"0f076b08",
			4807 => x"040bc404",
			4808 => x"ff7a4ca5",
			4809 => x"fdc64ca5",
			4810 => x"0e053b04",
			4811 => x"01f24ca5",
			4812 => x"00004ca5",
			4813 => x"0c049010",
			4814 => x"0d054c08",
			4815 => x"05052d04",
			4816 => x"00264ca5",
			4817 => x"fe994ca5",
			4818 => x"0b04c004",
			4819 => x"02064ca5",
			4820 => x"00004ca5",
			4821 => x"0b04af08",
			4822 => x"07049504",
			4823 => x"feef4ca5",
			4824 => x"01064ca5",
			4825 => x"06013e04",
			4826 => x"011a4ca5",
			4827 => x"fe214ca5",
			4828 => x"03053960",
			4829 => x"0b04c024",
			4830 => x"06013110",
			4831 => x"040ab204",
			4832 => x"fef04ca5",
			4833 => x"03052708",
			4834 => x"0f06bb04",
			4835 => x"01e44ca5",
			4836 => x"ffcf4ca5",
			4837 => x"023f4ca5",
			4838 => x"08031b04",
			4839 => x"fdf44ca5",
			4840 => x"00045f08",
			4841 => x"00045704",
			4842 => x"000c4ca5",
			4843 => x"fd7b4ca5",
			4844 => x"0c04af04",
			4845 => x"00ea4ca5",
			4846 => x"ff584ca5",
			4847 => x"0f06e320",
			4848 => x"03051b10",
			4849 => x"0e044408",
			4850 => x"06014e04",
			4851 => x"00ce4ca5",
			4852 => x"feca4ca5",
			4853 => x"0e047804",
			4854 => x"01d74ca5",
			4855 => x"00974ca5",
			4856 => x"09009b08",
			4857 => x"0c049404",
			4858 => x"fdd34ca5",
			4859 => x"ffa74ca5",
			4860 => x"040be904",
			4861 => x"00374ca5",
			4862 => x"01d94ca5",
			4863 => x"0f06f90c",
			4864 => x"0b04c304",
			4865 => x"017b4ca5",
			4866 => x"0e04a504",
			4867 => x"01a24ca5",
			4868 => x"03294ca5",
			4869 => x"0f071708",
			4870 => x"0f070f04",
			4871 => x"00d74ca5",
			4872 => x"feaf4ca5",
			4873 => x"06015204",
			4874 => x"02054ca5",
			4875 => x"00d74ca5",
			4876 => x"03053f10",
			4877 => x"02085908",
			4878 => x"0d056504",
			4879 => x"01d34ca5",
			4880 => x"fec74ca5",
			4881 => x"08036b04",
			4882 => x"fd244ca5",
			4883 => x"ff974ca5",
			4884 => x"0305430c",
			4885 => x"08036308",
			4886 => x"05055804",
			4887 => x"01034ca5",
			4888 => x"02704ca5",
			4889 => x"00004ca5",
			4890 => x"02084d10",
			4891 => x"08034508",
			4892 => x"0e04a504",
			4893 => x"02084ca5",
			4894 => x"ffd64ca5",
			4895 => x"03056104",
			4896 => x"fdcf4ca5",
			4897 => x"fff14ca5",
			4898 => x"0704bc08",
			4899 => x"03058004",
			4900 => x"00cc4ca5",
			4901 => x"00084ca5",
			4902 => x"0b04bf04",
			4903 => x"febd4ca5",
			4904 => x"000a4ca5",
			4905 => x"09007194",
			4906 => x"0e03e75c",
			4907 => x"0a02d42c",
			4908 => x"08036c14",
			4909 => x"01004510",
			4910 => x"0c045c08",
			4911 => x"06012b04",
			4912 => x"fd244f59",
			4913 => x"ffa54f59",
			4914 => x"07047804",
			4915 => x"fed84f59",
			4916 => x"01b54f59",
			4917 => x"fd604f59",
			4918 => x"0900550c",
			4919 => x"0e033e08",
			4920 => x"02082204",
			4921 => x"01d74f59",
			4922 => x"00004f59",
			4923 => x"fdeb4f59",
			4924 => x"02082408",
			4925 => x"01003c04",
			4926 => x"009a4f59",
			4927 => x"01b54f59",
			4928 => x"00374f59",
			4929 => x"05050e1c",
			4930 => x"07047a0c",
			4931 => x"02074b04",
			4932 => x"01714f59",
			4933 => x"0f069004",
			4934 => x"fdc84f59",
			4935 => x"00d84f59",
			4936 => x"06013d08",
			4937 => x"06013104",
			4938 => x"fec64f59",
			4939 => x"fc174f59",
			4940 => x"0c047a04",
			4941 => x"016c4f59",
			4942 => x"00004f59",
			4943 => x"0d051908",
			4944 => x"0d050c04",
			4945 => x"fe464f59",
			4946 => x"fb3c4f59",
			4947 => x"0c049204",
			4948 => x"01494f59",
			4949 => x"0207da04",
			4950 => x"007d4f59",
			4951 => x"fe154f59",
			4952 => x"08035620",
			4953 => x"08033010",
			4954 => x"0704950c",
			4955 => x"0a025904",
			4956 => x"ff604f59",
			4957 => x"0504f304",
			4958 => x"00004f59",
			4959 => x"fc4d4f59",
			4960 => x"01064f59",
			4961 => x"01003c04",
			4962 => x"fd5b4f59",
			4963 => x"0b047d04",
			4964 => x"ffee4f59",
			4965 => x"0f069904",
			4966 => x"00874f59",
			4967 => x"01fb4f59",
			4968 => x"0e03f104",
			4969 => x"fd234f59",
			4970 => x"09006f10",
			4971 => x"08038508",
			4972 => x"0a02a104",
			4973 => x"00324f59",
			4974 => x"fd844f59",
			4975 => x"040d6e04",
			4976 => x"00474f59",
			4977 => x"fdbc4f59",
			4978 => x"00344f59",
			4979 => x"0c047968",
			4980 => x"0704a83c",
			4981 => x"0601311c",
			4982 => x"0505110c",
			4983 => x"0c047808",
			4984 => x"08034804",
			4985 => x"feed4f59",
			4986 => x"01af4f59",
			4987 => x"fbfb4f59",
			4988 => x"0e048808",
			4989 => x"05053a04",
			4990 => x"00e64f59",
			4991 => x"fefc4f59",
			4992 => x"06012b04",
			4993 => x"fff84f59",
			4994 => x"fe5b4f59",
			4995 => x"0c047310",
			4996 => x"0a027d08",
			4997 => x"01005704",
			4998 => x"02d54f59",
			4999 => x"00004f59",
			5000 => x"0c045c04",
			5001 => x"00124f59",
			5002 => x"febc4f59",
			5003 => x"06013508",
			5004 => x"07049104",
			5005 => x"027b4f59",
			5006 => x"00a34f59",
			5007 => x"06013604",
			5008 => x"ff5a4f59",
			5009 => x"00ab4f59",
			5010 => x"0704c420",
			5011 => x"06014910",
			5012 => x"0c047408",
			5013 => x"01005304",
			5014 => x"010d4f59",
			5015 => x"028c4f59",
			5016 => x"0c047604",
			5017 => x"fff14f59",
			5018 => x"01424f59",
			5019 => x"0a02a808",
			5020 => x"05055704",
			5021 => x"fd474f59",
			5022 => x"ff9c4f59",
			5023 => x"02083d04",
			5024 => x"fe244f59",
			5025 => x"015f4f59",
			5026 => x"0a027204",
			5027 => x"002d4f59",
			5028 => x"040ba404",
			5029 => x"fd514f59",
			5030 => x"ff7d4f59",
			5031 => x"0c04902c",
			5032 => x"0505681c",
			5033 => x"09009310",
			5034 => x"05054808",
			5035 => x"05052004",
			5036 => x"000b4f59",
			5037 => x"fed24f59",
			5038 => x"02083804",
			5039 => x"02f14f59",
			5040 => x"00004f59",
			5041 => x"040afc04",
			5042 => x"00c64f59",
			5043 => x"0b04af04",
			5044 => x"ff254f59",
			5045 => x"fd764f59",
			5046 => x"0b04e208",
			5047 => x"0b04d304",
			5048 => x"ff494f59",
			5049 => x"03ac4f59",
			5050 => x"08033a04",
			5051 => x"ff454f59",
			5052 => x"fe294f59",
			5053 => x"0c049114",
			5054 => x"0d053404",
			5055 => x"02194f59",
			5056 => x"0b04b208",
			5057 => x"0b04af04",
			5058 => x"007d4f59",
			5059 => x"fda14f59",
			5060 => x"01006304",
			5061 => x"020c4f59",
			5062 => x"00204f59",
			5063 => x"09009710",
			5064 => x"0e04b408",
			5065 => x"09008f04",
			5066 => x"ffd04f59",
			5067 => x"008f4f59",
			5068 => x"0b049f04",
			5069 => x"01a54f59",
			5070 => x"ff1e4f59",
			5071 => x"0e04a008",
			5072 => x"0704bb04",
			5073 => x"023e4f59",
			5074 => x"00ad4f59",
			5075 => x"0c049204",
			5076 => x"01194f59",
			5077 => x"000b4f59",
			5078 => x"0e04bbbc",
			5079 => x"0f070568",
			5080 => x"040c4c38",
			5081 => x"03049718",
			5082 => x"08030808",
			5083 => x"0b049104",
			5084 => x"fdf0523d",
			5085 => x"015a523d",
			5086 => x"08036f08",
			5087 => x"07049304",
			5088 => x"0186523d",
			5089 => x"0069523d",
			5090 => x"0b048d04",
			5091 => x"0114523d",
			5092 => x"fdd4523d",
			5093 => x"0d056910",
			5094 => x"03051b08",
			5095 => x"0207da04",
			5096 => x"ffbe523d",
			5097 => x"0042523d",
			5098 => x"09008c04",
			5099 => x"fde0523d",
			5100 => x"ffc8523d",
			5101 => x"06014508",
			5102 => x"040a3a04",
			5103 => x"fe48523d",
			5104 => x"016b523d",
			5105 => x"0704bf04",
			5106 => x"fe35523d",
			5107 => x"0057523d",
			5108 => x"0004a31c",
			5109 => x"0d055c10",
			5110 => x"09008808",
			5111 => x"0304ef04",
			5112 => x"ff92523d",
			5113 => x"fe07523d",
			5114 => x"0c048f04",
			5115 => x"ffd3523d",
			5116 => x"018a523d",
			5117 => x"00048104",
			5118 => x"0063523d",
			5119 => x"0e047804",
			5120 => x"fcb1523d",
			5121 => x"ff18523d",
			5122 => x"040cbf08",
			5123 => x"0f06e504",
			5124 => x"01c4523d",
			5125 => x"0082523d",
			5126 => x"0e047108",
			5127 => x"07047a04",
			5128 => x"fe90523d",
			5129 => x"002a523d",
			5130 => x"fddd523d",
			5131 => x"0e04ad38",
			5132 => x"0e04a520",
			5133 => x"0704a610",
			5134 => x"01005208",
			5135 => x"09007704",
			5136 => x"ff66523d",
			5137 => x"00b6523d",
			5138 => x"03050d04",
			5139 => x"0158523d",
			5140 => x"feb4523d",
			5141 => x"0b04d108",
			5142 => x"0e049d04",
			5143 => x"017a523d",
			5144 => x"000c523d",
			5145 => x"06014a04",
			5146 => x"0118523d",
			5147 => x"fdbc523d",
			5148 => x"0601410c",
			5149 => x"08033904",
			5150 => x"feba523d",
			5151 => x"03052f04",
			5152 => x"00bd523d",
			5153 => x"0255523d",
			5154 => x"0b04e008",
			5155 => x"040ca004",
			5156 => x"fde5523d",
			5157 => x"0040523d",
			5158 => x"00a8523d",
			5159 => x"01004b04",
			5160 => x"fde9523d",
			5161 => x"0305330c",
			5162 => x"0b04bf08",
			5163 => x"00049204",
			5164 => x"024e523d",
			5165 => x"00dc523d",
			5166 => x"0000523d",
			5167 => x"0d054e04",
			5168 => x"feea523d",
			5169 => x"0f071104",
			5170 => x"ffa3523d",
			5171 => x"0191523d",
			5172 => x"09009e58",
			5173 => x"0f072d20",
			5174 => x"0208681c",
			5175 => x"0f06ea0c",
			5176 => x"09008a08",
			5177 => x"0002ee04",
			5178 => x"0000523d",
			5179 => x"00b2523d",
			5180 => x"fe0c523d",
			5181 => x"08031a08",
			5182 => x"0f070504",
			5183 => x"fefc523d",
			5184 => x"0137523d",
			5185 => x"03053304",
			5186 => x"0024523d",
			5187 => x"fec8523d",
			5188 => x"fd3f523d",
			5189 => x"06014f1c",
			5190 => x"0601300c",
			5191 => x"00041408",
			5192 => x"03056f04",
			5193 => x"008e523d",
			5194 => x"fe5d523d",
			5195 => x"fa3b523d",
			5196 => x"08033c08",
			5197 => x"03058904",
			5198 => x"0172523d",
			5199 => x"fec2523d",
			5200 => x"040bcc04",
			5201 => x"ff19523d",
			5202 => x"0033523d",
			5203 => x"0004960c",
			5204 => x"03055304",
			5205 => x"0025523d",
			5206 => x"040c4c04",
			5207 => x"fea0523d",
			5208 => x"fd13523d",
			5209 => x"09009808",
			5210 => x"0b04b004",
			5211 => x"01c2523d",
			5212 => x"fde5523d",
			5213 => x"0c04b304",
			5214 => x"019a523d",
			5215 => x"0035523d",
			5216 => x"0305612c",
			5217 => x"0900a91c",
			5218 => x"0b04c10c",
			5219 => x"06013d04",
			5220 => x"02d1523d",
			5221 => x"0f071f04",
			5222 => x"ff53523d",
			5223 => x"0240523d",
			5224 => x"01006208",
			5225 => x"0b04cf04",
			5226 => x"fffe523d",
			5227 => x"01ff523d",
			5228 => x"06014104",
			5229 => x"fe2a523d",
			5230 => x"0082523d",
			5231 => x"0d057604",
			5232 => x"03ae523d",
			5233 => x"0e04f708",
			5234 => x"0003ee04",
			5235 => x"0092523d",
			5236 => x"021a523d",
			5237 => x"0000523d",
			5238 => x"01006218",
			5239 => x"040bde0c",
			5240 => x"0d058308",
			5241 => x"0f074f04",
			5242 => x"ff4c523d",
			5243 => x"014f523d",
			5244 => x"fe19523d",
			5245 => x"0f07a308",
			5246 => x"0704bc04",
			5247 => x"0305523d",
			5248 => x"01d7523d",
			5249 => x"ff01523d",
			5250 => x"0900a80c",
			5251 => x"01006304",
			5252 => x"fd64523d",
			5253 => x"02090504",
			5254 => x"ff65523d",
			5255 => x"0211523d",
			5256 => x"0b04c008",
			5257 => x"0704bc04",
			5258 => x"fdae523d",
			5259 => x"ffa4523d",
			5260 => x"0b04e104",
			5261 => x"0077523d",
			5262 => x"fff9523d",
			5263 => x"0f0773d8",
			5264 => x"03050074",
			5265 => x"0900823c",
			5266 => x"0b04af1c",
			5267 => x"0304ef10",
			5268 => x"0b049108",
			5269 => x"0f06ed04",
			5270 => x"ffc5551b",
			5271 => x"00d7551b",
			5272 => x"0f06b504",
			5273 => x"0023551b",
			5274 => x"011f551b",
			5275 => x"0c045704",
			5276 => x"01f7551b",
			5277 => x"06013e04",
			5278 => x"fe0a551b",
			5279 => x"0034551b",
			5280 => x"0d054110",
			5281 => x"0a02bc08",
			5282 => x"0e046104",
			5283 => x"0001551b",
			5284 => x"fe46551b",
			5285 => x"09007d04",
			5286 => x"0000551b",
			5287 => x"fd02551b",
			5288 => x"0f069f08",
			5289 => x"0a031504",
			5290 => x"01a4551b",
			5291 => x"ff09551b",
			5292 => x"0304be04",
			5293 => x"00d1551b",
			5294 => x"fdd9551b",
			5295 => x"0c047818",
			5296 => x"0004350c",
			5297 => x"0704aa08",
			5298 => x"0a027404",
			5299 => x"00a8551b",
			5300 => x"fe62551b",
			5301 => x"0219551b",
			5302 => x"0d052604",
			5303 => x"0013551b",
			5304 => x"0f06b204",
			5305 => x"0116551b",
			5306 => x"020a551b",
			5307 => x"09008610",
			5308 => x"040c1208",
			5309 => x"06012004",
			5310 => x"0000551b",
			5311 => x"01fd551b",
			5312 => x"07049504",
			5313 => x"fe9a551b",
			5314 => x"00ec551b",
			5315 => x"05054908",
			5316 => x"00047104",
			5317 => x"ff2c551b",
			5318 => x"0082551b",
			5319 => x"0704bb04",
			5320 => x"01e5551b",
			5321 => x"0019551b",
			5322 => x"07049028",
			5323 => x"0f073b18",
			5324 => x"0a027b0c",
			5325 => x"00040708",
			5326 => x"0e04e204",
			5327 => x"fe3c551b",
			5328 => x"0000551b",
			5329 => x"013e551b",
			5330 => x"0e048f04",
			5331 => x"fd94551b",
			5332 => x"03051b04",
			5333 => x"ffeb551b",
			5334 => x"fe25551b",
			5335 => x"040b9104",
			5336 => x"0262551b",
			5337 => x"03051b04",
			5338 => x"0180551b",
			5339 => x"0b049e04",
			5340 => x"fff3551b",
			5341 => x"fd91551b",
			5342 => x"09009520",
			5343 => x"0b049f10",
			5344 => x"0c049308",
			5345 => x"0a028704",
			5346 => x"01ec551b",
			5347 => x"ffa6551b",
			5348 => x"00045804",
			5349 => x"00dc551b",
			5350 => x"0252551b",
			5351 => x"0704a808",
			5352 => x"0f072504",
			5353 => x"feda551b",
			5354 => x"ffdc551b",
			5355 => x"0b04d204",
			5356 => x"fffa551b",
			5357 => x"fe77551b",
			5358 => x"0704ad0c",
			5359 => x"0c04b408",
			5360 => x"0003f204",
			5361 => x"ff90551b",
			5362 => x"00bd551b",
			5363 => x"fe5e551b",
			5364 => x"0704bb08",
			5365 => x"0e051004",
			5366 => x"fd38551b",
			5367 => x"0000551b",
			5368 => x"0704ed04",
			5369 => x"ffd4551b",
			5370 => x"0061551b",
			5371 => x"0e059d54",
			5372 => x"00043e24",
			5373 => x"0c04d220",
			5374 => x"0e057810",
			5375 => x"05058408",
			5376 => x"06014504",
			5377 => x"0017551b",
			5378 => x"0307551b",
			5379 => x"0704bf04",
			5380 => x"fe5c551b",
			5381 => x"00d8551b",
			5382 => x"0a027208",
			5383 => x"0d05a904",
			5384 => x"0254551b",
			5385 => x"ff92551b",
			5386 => x"0f07b204",
			5387 => x"fe5d551b",
			5388 => x"009d551b",
			5389 => x"02bb551b",
			5390 => x"040bca10",
			5391 => x"0803610c",
			5392 => x"0305a908",
			5393 => x"0f078e04",
			5394 => x"fe2c551b",
			5395 => x"00d2551b",
			5396 => x"fdd3551b",
			5397 => x"0019551b",
			5398 => x"0900b510",
			5399 => x"0c04d108",
			5400 => x"0f07ce04",
			5401 => x"005b551b",
			5402 => x"ff2e551b",
			5403 => x"040c6c04",
			5404 => x"fdc4551b",
			5405 => x"00b6551b",
			5406 => x"0505b108",
			5407 => x"0b051204",
			5408 => x"00aa551b",
			5409 => x"021e551b",
			5410 => x"0305d904",
			5411 => x"fc2a551b",
			5412 => x"0047551b",
			5413 => x"0e05ac20",
			5414 => x"0c04cf14",
			5415 => x"0505af10",
			5416 => x"0305e908",
			5417 => x"0305d104",
			5418 => x"ff0d551b",
			5419 => x"0196551b",
			5420 => x"08036104",
			5421 => x"ff39551b",
			5422 => x"fdf2551b",
			5423 => x"01cf551b",
			5424 => x"0900cb04",
			5425 => x"fd86551b",
			5426 => x"0b058704",
			5427 => x"00c8551b",
			5428 => x"0000551b",
			5429 => x"0704aa04",
			5430 => x"fe3c551b",
			5431 => x"05059310",
			5432 => x"040b9d08",
			5433 => x"040af504",
			5434 => x"01a0551b",
			5435 => x"fefb551b",
			5436 => x"0305f904",
			5437 => x"0000551b",
			5438 => x"02aa551b",
			5439 => x"0d05ca08",
			5440 => x"0f081604",
			5441 => x"feb6551b",
			5442 => x"0144551b",
			5443 => x"0b052004",
			5444 => x"0099551b",
			5445 => x"fff9551b",
			5446 => x"07056158",
			5447 => x"040eab3c",
			5448 => x"03040e08",
			5449 => x"0d04db04",
			5450 => x"00db564d",
			5451 => x"021c564d",
			5452 => x"09006214",
			5453 => x"03043708",
			5454 => x"07047b04",
			5455 => x"ff9d564d",
			5456 => x"01f4564d",
			5457 => x"0f064a04",
			5458 => x"fc83564d",
			5459 => x"040c0404",
			5460 => x"0006564d",
			5461 => x"fe18564d",
			5462 => x"03048f10",
			5463 => x"0f065208",
			5464 => x"01004504",
			5465 => x"00f9564d",
			5466 => x"ff9f564d",
			5467 => x"0803ac04",
			5468 => x"018d564d",
			5469 => x"ffa3564d",
			5470 => x"09007508",
			5471 => x"0304c004",
			5472 => x"ffd9564d",
			5473 => x"fe60564d",
			5474 => x"03050004",
			5475 => x"0074564d",
			5476 => x"0024564d",
			5477 => x"06014a08",
			5478 => x"0d054c04",
			5479 => x"fe56564d",
			5480 => x"fff9564d",
			5481 => x"07049504",
			5482 => x"0146564d",
			5483 => x"0e044b04",
			5484 => x"fd51564d",
			5485 => x"06016808",
			5486 => x"0803d004",
			5487 => x"ff55564d",
			5488 => x"011e564d",
			5489 => x"fe66564d",
			5490 => x"08032610",
			5491 => x"0901430c",
			5492 => x"09012704",
			5493 => x"fe6b564d",
			5494 => x"0f07c004",
			5495 => x"feec564d",
			5496 => x"01dc564d",
			5497 => x"fe64564d",
			5498 => x"040fc628",
			5499 => x"0a02e818",
			5500 => x"040d4210",
			5501 => x"0e0a1b08",
			5502 => x"0b067d04",
			5503 => x"0011564d",
			5504 => x"018a564d",
			5505 => x"0b079504",
			5506 => x"fe67564d",
			5507 => x"00de564d",
			5508 => x"0a02dd04",
			5509 => x"fe3b564d",
			5510 => x"ffe1564d",
			5511 => x"0f0c3908",
			5512 => x"0004a004",
			5513 => x"012c564d",
			5514 => x"0245564d",
			5515 => x"07075204",
			5516 => x"fe75564d",
			5517 => x"025c564d",
			5518 => x"04110308",
			5519 => x"0005b004",
			5520 => x"fe93564d",
			5521 => x"01c7564d",
			5522 => x"fe67564d",
			5523 => x"07057760",
			5524 => x"01003920",
			5525 => x"01002504",
			5526 => x"fe555789",
			5527 => x"0304350c",
			5528 => x"0b046d04",
			5529 => x"fec65789",
			5530 => x"01002a04",
			5531 => x"000c5789",
			5532 => x"023b5789",
			5533 => x"0a02bc0c",
			5534 => x"08038a08",
			5535 => x"07049204",
			5536 => x"fe485789",
			5537 => x"ffd15789",
			5538 => x"00005789",
			5539 => x"fd4f5789",
			5540 => x"00049624",
			5541 => x"00034b04",
			5542 => x"fe655789",
			5543 => x"06013510",
			5544 => x"0d059b08",
			5545 => x"03055304",
			5546 => x"01145789",
			5547 => x"fff75789",
			5548 => x"0b053104",
			5549 => x"02715789",
			5550 => x"00d75789",
			5551 => x"040b4a08",
			5552 => x"0c050504",
			5553 => x"ffae5789",
			5554 => x"01d85789",
			5555 => x"0704be04",
			5556 => x"00735789",
			5557 => x"00e65789",
			5558 => x"0410bb18",
			5559 => x"040c790c",
			5560 => x"0900be08",
			5561 => x"0f075d04",
			5562 => x"02525789",
			5563 => x"00c65789",
			5564 => x"02f95789",
			5565 => x"07047804",
			5566 => x"00005789",
			5567 => x"040df504",
			5568 => x"01715789",
			5569 => x"00875789",
			5570 => x"fe6f5789",
			5571 => x"0803260c",
			5572 => x"0100c308",
			5573 => x"0100bd04",
			5574 => x"fe6c5789",
			5575 => x"03645789",
			5576 => x"fe565789",
			5577 => x"040e6328",
			5578 => x"08034c14",
			5579 => x"01011908",
			5580 => x"040c2604",
			5581 => x"03cc5789",
			5582 => x"fe745789",
			5583 => x"0c06c708",
			5584 => x"08032804",
			5585 => x"00ee5789",
			5586 => x"fe565789",
			5587 => x"02345789",
			5588 => x"0f0c9c10",
			5589 => x"0c061408",
			5590 => x"09015804",
			5591 => x"02cb5789",
			5592 => x"ff905789",
			5593 => x"040cb604",
			5594 => x"048d5789",
			5595 => x"00f65789",
			5596 => x"feba5789",
			5597 => x"04110308",
			5598 => x"0410e104",
			5599 => x"fe7e5789",
			5600 => x"ff455789",
			5601 => x"fe555789",
			5602 => x"07057760",
			5603 => x"040eab44",
			5604 => x"06010a08",
			5605 => x"06010604",
			5606 => x"fe5858bd",
			5607 => x"ffb558bd",
			5608 => x"0e054b20",
			5609 => x"0900b510",
			5610 => x"040c2608",
			5611 => x"06013e04",
			5612 => x"010c58bd",
			5613 => x"003358bd",
			5614 => x"09008f04",
			5615 => x"010758bd",
			5616 => x"01a158bd",
			5617 => x"05058308",
			5618 => x"040bb204",
			5619 => x"050d58bd",
			5620 => x"02f458bd",
			5621 => x"040b5b04",
			5622 => x"010358bd",
			5623 => x"025158bd",
			5624 => x"0c04e710",
			5625 => x"06016c08",
			5626 => x"0704d604",
			5627 => x"ffc058bd",
			5628 => x"00a458bd",
			5629 => x"07051804",
			5630 => x"fea658bd",
			5631 => x"005258bd",
			5632 => x"09014208",
			5633 => x"06015604",
			5634 => x"006f58bd",
			5635 => x"016a58bd",
			5636 => x"fe4758bd",
			5637 => x"06014a08",
			5638 => x"0b04c004",
			5639 => x"fe5058bd",
			5640 => x"fef658bd",
			5641 => x"07049504",
			5642 => x"01b458bd",
			5643 => x"040f0204",
			5644 => x"009358bd",
			5645 => x"09007508",
			5646 => x"09003004",
			5647 => x"fe7b58bd",
			5648 => x"ffcd58bd",
			5649 => x"fe3a58bd",
			5650 => x"0803260c",
			5651 => x"0c054608",
			5652 => x"0705a104",
			5653 => x"fe8f58bd",
			5654 => x"018958bd",
			5655 => x"fe5158bd",
			5656 => x"040e632c",
			5657 => x"08035218",
			5658 => x"0f0ad90c",
			5659 => x"040c6008",
			5660 => x"0901db04",
			5661 => x"031b58bd",
			5662 => x"ff6a58bd",
			5663 => x"fe6458bd",
			5664 => x"08032804",
			5665 => x"000058bd",
			5666 => x"07073804",
			5667 => x"fe5058bd",
			5668 => x"000058bd",
			5669 => x"0c054c04",
			5670 => x"feb958bd",
			5671 => x"0f0c3908",
			5672 => x"0d093404",
			5673 => x"015b58bd",
			5674 => x"03ab58bd",
			5675 => x"0601d004",
			5676 => x"fe1d58bd",
			5677 => x"017658bd",
			5678 => x"fe5658bd",
			5679 => x"040d5574",
			5680 => x"0004b84c",
			5681 => x"040a011c",
			5682 => x"0802c318",
			5683 => x"0409b30c",
			5684 => x"0305e108",
			5685 => x"01006304",
			5686 => x"fe645a61",
			5687 => x"012f5a61",
			5688 => x"fe505a61",
			5689 => x"01008a08",
			5690 => x"0704bf04",
			5691 => x"000c5a61",
			5692 => x"02105a61",
			5693 => x"fe985a61",
			5694 => x"fdc75a61",
			5695 => x"0802d510",
			5696 => x"0b05a80c",
			5697 => x"0d05a708",
			5698 => x"03058904",
			5699 => x"01685a61",
			5700 => x"febf5a61",
			5701 => x"025a5a61",
			5702 => x"fe7d5a61",
			5703 => x"0207da10",
			5704 => x"040c7208",
			5705 => x"01006804",
			5706 => x"ffe95a61",
			5707 => x"fdfd5a61",
			5708 => x"03043704",
			5709 => x"01855a61",
			5710 => x"fd5e5a61",
			5711 => x"01004108",
			5712 => x"03049f04",
			5713 => x"ffab5a61",
			5714 => x"fe375a61",
			5715 => x"0304b704",
			5716 => x"00ea5a61",
			5717 => x"00155a61",
			5718 => x"0e04b41c",
			5719 => x"0b047d0c",
			5720 => x"0504e708",
			5721 => x"0504e204",
			5722 => x"01d25a61",
			5723 => x"00a85a61",
			5724 => x"fec45a61",
			5725 => x"0803c70c",
			5726 => x"0704a904",
			5727 => x"01e05a61",
			5728 => x"0e043604",
			5729 => x"ffbd5a61",
			5730 => x"01b15a61",
			5731 => x"00005a61",
			5732 => x"0e04d304",
			5733 => x"fcaf5a61",
			5734 => x"01006d04",
			5735 => x"01bd5a61",
			5736 => x"ff8a5a61",
			5737 => x"0f075530",
			5738 => x"01005524",
			5739 => x"07047b10",
			5740 => x"0e036108",
			5741 => x"07047904",
			5742 => x"fe775a61",
			5743 => x"00005a61",
			5744 => x"0b047104",
			5745 => x"fedb5a61",
			5746 => x"fc245a61",
			5747 => x"040d8804",
			5748 => x"01175a61",
			5749 => x"02082f08",
			5750 => x"0e033e04",
			5751 => x"fe6d5a61",
			5752 => x"00cf5a61",
			5753 => x"02083704",
			5754 => x"fc665a61",
			5755 => x"ff085a61",
			5756 => x"0c04af04",
			5757 => x"faa35a61",
			5758 => x"03055804",
			5759 => x"014f5a61",
			5760 => x"00005a61",
			5761 => x"07057318",
			5762 => x"02091908",
			5763 => x"03056f04",
			5764 => x"02045a61",
			5765 => x"fde55a61",
			5766 => x"0004b804",
			5767 => x"ff425a61",
			5768 => x"040f0208",
			5769 => x"07050604",
			5770 => x"01665a61",
			5771 => x"027f5a61",
			5772 => x"ff695a61",
			5773 => x"08039c04",
			5774 => x"fe5f5a61",
			5775 => x"0c06320c",
			5776 => x"0506f108",
			5777 => x"0e05ac04",
			5778 => x"00005a61",
			5779 => x"feec5a61",
			5780 => x"018a5a61",
			5781 => x"0e09c104",
			5782 => x"00005a61",
			5783 => x"fea75a61",
			5784 => x"07057760",
			5785 => x"040eab48",
			5786 => x"06010a08",
			5787 => x"06010604",
			5788 => x"fe545b9d",
			5789 => x"ff9e5b9d",
			5790 => x"0e04e220",
			5791 => x"0704a710",
			5792 => x"0304c008",
			5793 => x"0c045504",
			5794 => x"ffdc5b9d",
			5795 => x"01865b9d",
			5796 => x"09007504",
			5797 => x"fe7e5b9d",
			5798 => x"00e35b9d",
			5799 => x"02086f08",
			5800 => x"06012d04",
			5801 => x"01e35b9d",
			5802 => x"01265b9d",
			5803 => x"00044604",
			5804 => x"03785b9d",
			5805 => x"01f05b9d",
			5806 => x"040bb210",
			5807 => x"0c04e908",
			5808 => x"0a028504",
			5809 => x"00715b9d",
			5810 => x"ff435b9d",
			5811 => x"09013d04",
			5812 => x"01935b9d",
			5813 => x"fe4b5b9d",
			5814 => x"06017108",
			5815 => x"0900b304",
			5816 => x"00c35b9d",
			5817 => x"01735b9d",
			5818 => x"0c04f104",
			5819 => x"feff5b9d",
			5820 => x"015b5b9d",
			5821 => x"06014a04",
			5822 => x"fe4e5b9d",
			5823 => x"07049504",
			5824 => x"01e35b9d",
			5825 => x"040f0204",
			5826 => x"00b25b9d",
			5827 => x"09007508",
			5828 => x"09003004",
			5829 => x"fe715b9d",
			5830 => x"ffc25b9d",
			5831 => x"fe3a5b9d",
			5832 => x"0803260c",
			5833 => x"0c054608",
			5834 => x"0705a104",
			5835 => x"fe815b9d",
			5836 => x"01d85b9d",
			5837 => x"fe4c5b9d",
			5838 => x"040e6330",
			5839 => x"08035218",
			5840 => x"0f0ad90c",
			5841 => x"040c6008",
			5842 => x"040ba404",
			5843 => x"ffba5b9d",
			5844 => x"03c85b9d",
			5845 => x"fe5e5b9d",
			5846 => x"08032804",
			5847 => x"00005b9d",
			5848 => x"07073804",
			5849 => x"fe4b5b9d",
			5850 => x"00005b9d",
			5851 => x"08039c10",
			5852 => x"040d5508",
			5853 => x"040c1204",
			5854 => x"ff5c5b9d",
			5855 => x"01ca5b9d",
			5856 => x"00045404",
			5857 => x"00005b9d",
			5858 => x"fdff5b9d",
			5859 => x"0100ef04",
			5860 => x"01685b9d",
			5861 => x"03475b9d",
			5862 => x"fe515b9d",
			5863 => x"0b05856c",
			5864 => x"01003218",
			5865 => x"0601390c",
			5866 => x"040cf508",
			5867 => x"040c8504",
			5868 => x"fe895d19",
			5869 => x"00145d19",
			5870 => x"fe445d19",
			5871 => x"0d050f08",
			5872 => x"0303bd04",
			5873 => x"02105d19",
			5874 => x"ff1b5d19",
			5875 => x"fe425d19",
			5876 => x"0e04bb24",
			5877 => x"06010a04",
			5878 => x"fe485d19",
			5879 => x"0d054d10",
			5880 => x"0304fe08",
			5881 => x"0b047d04",
			5882 => x"01065d19",
			5883 => x"01e35d19",
			5884 => x"0004a004",
			5885 => x"00aa5d19",
			5886 => x"023f5d19",
			5887 => x"06012808",
			5888 => x"0e047f04",
			5889 => x"02c55d19",
			5890 => x"034f5d19",
			5891 => x"0f06ac04",
			5892 => x"00eb5d19",
			5893 => x"02295d19",
			5894 => x"040bd814",
			5895 => x"06010e04",
			5896 => x"fe4e5d19",
			5897 => x"06013a08",
			5898 => x"0f06ed04",
			5899 => x"ffd95d19",
			5900 => x"01aa5d19",
			5901 => x"00046004",
			5902 => x"00225d19",
			5903 => x"03385d19",
			5904 => x"06017110",
			5905 => x"0b04c008",
			5906 => x"05051d04",
			5907 => x"fe885d19",
			5908 => x"00c25d19",
			5909 => x"040c6004",
			5910 => x"01755d19",
			5911 => x"023e5d19",
			5912 => x"0f090508",
			5913 => x"0f07eb04",
			5914 => x"ffe35d19",
			5915 => x"fe915d19",
			5916 => x"01035d19",
			5917 => x"0c05602c",
			5918 => x"0f084f10",
			5919 => x"05061504",
			5920 => x"00195d19",
			5921 => x"0f080e04",
			5922 => x"fe4a5d19",
			5923 => x"0b059604",
			5924 => x"01235d19",
			5925 => x"fe485d19",
			5926 => x"09014714",
			5927 => x"040f0210",
			5928 => x"0f090d08",
			5929 => x"0d069f04",
			5930 => x"02e55d19",
			5931 => x"ff8e5d19",
			5932 => x"00043f04",
			5933 => x"044c5d19",
			5934 => x"01bd5d19",
			5935 => x"fe815d19",
			5936 => x"00047d04",
			5937 => x"fe315d19",
			5938 => x"006d5d19",
			5939 => x"08032604",
			5940 => x"fe425d19",
			5941 => x"040eab20",
			5942 => x"0e0a2a10",
			5943 => x"040cce08",
			5944 => x"0901d004",
			5945 => x"03445d19",
			5946 => x"00775d19",
			5947 => x"0a02cc04",
			5948 => x"feb95d19",
			5949 => x"035e5d19",
			5950 => x"0601c008",
			5951 => x"0c06de04",
			5952 => x"fe545d19",
			5953 => x"018f5d19",
			5954 => x"08037304",
			5955 => x"ff685d19",
			5956 => x"02865d19",
			5957 => x"fe425d19",
			5958 => x"07056180",
			5959 => x"040eab60",
			5960 => x"03048f20",
			5961 => x"0c045510",
			5962 => x"0207b504",
			5963 => x"006d5ead",
			5964 => x"0f06a508",
			5965 => x"0504e204",
			5966 => x"01545ead",
			5967 => x"fd1a5ead",
			5968 => x"015e5ead",
			5969 => x"0a024504",
			5970 => x"fe195ead",
			5971 => x"0f069908",
			5972 => x"02082a04",
			5973 => x"00e55ead",
			5974 => x"feb25ead",
			5975 => x"021c5ead",
			5976 => x"09007520",
			5977 => x"0304c010",
			5978 => x"0b047108",
			5979 => x"03049f04",
			5980 => x"013b5ead",
			5981 => x"fd405ead",
			5982 => x"02081d04",
			5983 => x"ff195ead",
			5984 => x"00e65ead",
			5985 => x"0f06d008",
			5986 => x"05050f04",
			5987 => x"fbce5ead",
			5988 => x"fdfa5ead",
			5989 => x"09007104",
			5990 => x"fd555ead",
			5991 => x"ff9f5ead",
			5992 => x"03050010",
			5993 => x"0f06d608",
			5994 => x"0a027d04",
			5995 => x"00de5ead",
			5996 => x"00015ead",
			5997 => x"09008204",
			5998 => x"00ab5ead",
			5999 => x"01895ead",
			6000 => x"0d054d08",
			6001 => x"09009504",
			6002 => x"ff825ead",
			6003 => x"00d15ead",
			6004 => x"0c045b04",
			6005 => x"02d45ead",
			6006 => x"00395ead",
			6007 => x"06014a08",
			6008 => x"0d054c04",
			6009 => x"fe565ead",
			6010 => x"ffc35ead",
			6011 => x"07049504",
			6012 => x"015f5ead",
			6013 => x"0a02f708",
			6014 => x"0c050c04",
			6015 => x"008b5ead",
			6016 => x"ff455ead",
			6017 => x"0c04b604",
			6018 => x"fd045ead",
			6019 => x"03055f04",
			6020 => x"00065ead",
			6021 => x"fe815ead",
			6022 => x"08032610",
			6023 => x"0100c30c",
			6024 => x"09012704",
			6025 => x"fe595ead",
			6026 => x"0207fa04",
			6027 => x"fece5ead",
			6028 => x"02155ead",
			6029 => x"fe635ead",
			6030 => x"040fc62c",
			6031 => x"0c054c10",
			6032 => x"040df508",
			6033 => x"0a028e04",
			6034 => x"00005ead",
			6035 => x"fe0d5ead",
			6036 => x"0100df04",
			6037 => x"fefe5ead",
			6038 => x"00f65ead",
			6039 => x"0100c30c",
			6040 => x"05075608",
			6041 => x"0b05e704",
			6042 => x"01b05ead",
			6043 => x"03865ead",
			6044 => x"fee25ead",
			6045 => x"0c06c208",
			6046 => x"0901db04",
			6047 => x"00845ead",
			6048 => x"ff205ead",
			6049 => x"01014704",
			6050 => x"ff8d5ead",
			6051 => x"01e75ead",
			6052 => x"0411030c",
			6053 => x"0c057f08",
			6054 => x"0803d004",
			6055 => x"ffc75ead",
			6056 => x"02b85ead",
			6057 => x"fe865ead",
			6058 => x"fe655ead",
			6059 => x"03044e48",
			6060 => x"0e03793c",
			6061 => x"03041d24",
			6062 => x"02078008",
			6063 => x"0f053704",
			6064 => x"00006061",
			6065 => x"01af6061",
			6066 => x"0f05e00c",
			6067 => x"06014e08",
			6068 => x"0f05da04",
			6069 => x"fe656061",
			6070 => x"00006061",
			6071 => x"00006061",
			6072 => x"0c047308",
			6073 => x"0004d204",
			6074 => x"00f26061",
			6075 => x"ff156061",
			6076 => x"04108904",
			6077 => x"01846061",
			6078 => x"00006061",
			6079 => x"0d04e508",
			6080 => x"0b046004",
			6081 => x"febf6061",
			6082 => x"fa9b6061",
			6083 => x"0b048e08",
			6084 => x"07046304",
			6085 => x"00006061",
			6086 => x"fef06061",
			6087 => x"0410e104",
			6088 => x"011b6061",
			6089 => x"00006061",
			6090 => x"06011904",
			6091 => x"fea16061",
			6092 => x"02083104",
			6093 => x"01c86061",
			6094 => x"ffed6061",
			6095 => x"0f064a38",
			6096 => x"06012d18",
			6097 => x"0d052608",
			6098 => x"03047704",
			6099 => x"006c6061",
			6100 => x"fe126061",
			6101 => x"0704a508",
			6102 => x"09008004",
			6103 => x"014d6061",
			6104 => x"feb86061",
			6105 => x"00034b04",
			6106 => x"ffbf6061",
			6107 => x"01b06061",
			6108 => x"0b047e04",
			6109 => x"00c06061",
			6110 => x"0004a00c",
			6111 => x"040c3808",
			6112 => x"02079204",
			6113 => x"fdc96061",
			6114 => x"00006061",
			6115 => x"fc6d6061",
			6116 => x"0f064208",
			6117 => x"00053e04",
			6118 => x"01826061",
			6119 => x"00006061",
			6120 => x"06014604",
			6121 => x"00006061",
			6122 => x"fd396061",
			6123 => x"03049f20",
			6124 => x"08031d08",
			6125 => x"03048f04",
			6126 => x"fc1b6061",
			6127 => x"00006061",
			6128 => x"040c4708",
			6129 => x"0c049404",
			6130 => x"01c96061",
			6131 => x"ff226061",
			6132 => x"00048608",
			6133 => x"0f069004",
			6134 => x"fe4c6061",
			6135 => x"00d96061",
			6136 => x"07047c04",
			6137 => x"ff996061",
			6138 => x"00ff6061",
			6139 => x"0900791c",
			6140 => x"0208110c",
			6141 => x"0e03f904",
			6142 => x"00fa6061",
			6143 => x"040bbf04",
			6144 => x"ffb16061",
			6145 => x"fdcc6061",
			6146 => x"0304be08",
			6147 => x"02084404",
			6148 => x"019a6061",
			6149 => x"ffc16061",
			6150 => x"0f06d004",
			6151 => x"fe256061",
			6152 => x"ffb56061",
			6153 => x"0e057810",
			6154 => x"0f07a608",
			6155 => x"0c045504",
			6156 => x"fea66061",
			6157 => x"000f6061",
			6158 => x"0a028e04",
			6159 => x"02556061",
			6160 => x"00536061",
			6161 => x"0704ec08",
			6162 => x"0704da04",
			6163 => x"ffd66061",
			6164 => x"ff186061",
			6165 => x"0f074104",
			6166 => x"02276061",
			6167 => x"fff56061",
			6168 => x"05061588",
			6169 => x"01003614",
			6170 => x"06013508",
			6171 => x"02071704",
			6172 => x"ff4d622d",
			6173 => x"fe2a622d",
			6174 => x"01002504",
			6175 => x"fe30622d",
			6176 => x"07047a04",
			6177 => x"ff81622d",
			6178 => x"03f1622d",
			6179 => x"0e051d34",
			6180 => x"00045f1c",
			6181 => x"0e04780c",
			6182 => x"06010604",
			6183 => x"fe4b622d",
			6184 => x"0a029d04",
			6185 => x"0336622d",
			6186 => x"ff9b622d",
			6187 => x"0704a708",
			6188 => x"06014104",
			6189 => x"012c622d",
			6190 => x"ff5d622d",
			6191 => x"02084d04",
			6192 => x"01b9622d",
			6193 => x"02ef622d",
			6194 => x"0c045408",
			6195 => x"02080704",
			6196 => x"021f622d",
			6197 => x"fed6622d",
			6198 => x"05054b08",
			6199 => x"0e049604",
			6200 => x"0316622d",
			6201 => x"020d622d",
			6202 => x"0b053104",
			6203 => x"038d622d",
			6204 => x"fe6b622d",
			6205 => x"00044a20",
			6206 => x"02087e10",
			6207 => x"0704d708",
			6208 => x"0e058e04",
			6209 => x"ff90622d",
			6210 => x"fe1e622d",
			6211 => x"02079b04",
			6212 => x"fe46622d",
			6213 => x"00ec622d",
			6214 => x"06014208",
			6215 => x"05057504",
			6216 => x"008f622d",
			6217 => x"0574622d",
			6218 => x"0c04d404",
			6219 => x"0036622d",
			6220 => x"023b622d",
			6221 => x"06017310",
			6222 => x"0c04d208",
			6223 => x"00048204",
			6224 => x"0191622d",
			6225 => x"02db622d",
			6226 => x"01008004",
			6227 => x"033c622d",
			6228 => x"045a622d",
			6229 => x"07051808",
			6230 => x"02099504",
			6231 => x"fe20622d",
			6232 => x"ff99622d",
			6233 => x"06018004",
			6234 => x"0486622d",
			6235 => x"ff42622d",
			6236 => x"07057738",
			6237 => x"0e065a14",
			6238 => x"05061608",
			6239 => x"0305e904",
			6240 => x"fe7f622d",
			6241 => x"01c7622d",
			6242 => x"0208c004",
			6243 => x"fe3e622d",
			6244 => x"0004dd04",
			6245 => x"02df622d",
			6246 => x"fe58622d",
			6247 => x"09013118",
			6248 => x"07051f0c",
			6249 => x"06017004",
			6250 => x"01dd622d",
			6251 => x"01009904",
			6252 => x"010c622d",
			6253 => x"fe53622d",
			6254 => x"00039504",
			6255 => x"fe3d622d",
			6256 => x"08039004",
			6257 => x"038d622d",
			6258 => x"ff8b622d",
			6259 => x"00047d08",
			6260 => x"0c056004",
			6261 => x"fe23622d",
			6262 => x"013e622d",
			6263 => x"0202622d",
			6264 => x"09026b20",
			6265 => x"0803260c",
			6266 => x"0c054608",
			6267 => x"0c054304",
			6268 => x"fe4c622d",
			6269 => x"00c7622d",
			6270 => x"fe27622d",
			6271 => x"0004dd10",
			6272 => x"08035608",
			6273 => x"09015a04",
			6274 => x"03bf622d",
			6275 => x"fe6a622d",
			6276 => x"020c2a04",
			6277 => x"0208622d",
			6278 => x"ff53622d",
			6279 => x"fe28622d",
			6280 => x"07072204",
			6281 => x"fe31622d",
			6282 => x"021f622d",
			6283 => x"0506158c",
			6284 => x"0100391c",
			6285 => x"01002504",
			6286 => x"fe3263f9",
			6287 => x"0f06200c",
			6288 => x"07047804",
			6289 => x"ffd063f9",
			6290 => x"0207d104",
			6291 => x"03d063f9",
			6292 => x"016863f9",
			6293 => x"02083108",
			6294 => x"00047d04",
			6295 => x"fe0763f9",
			6296 => x"004e63f9",
			6297 => x"fe2b63f9",
			6298 => x"040c0c3c",
			6299 => x"0305391c",
			6300 => x"0304d80c",
			6301 => x"0802d404",
			6302 => x"ff9963f9",
			6303 => x"0a029e04",
			6304 => x"02c963f9",
			6305 => x"006963f9",
			6306 => x"0b04bf08",
			6307 => x"0f073904",
			6308 => x"014063f9",
			6309 => x"03dc63f9",
			6310 => x"0802e904",
			6311 => x"040263f9",
			6312 => x"022a63f9",
			6313 => x"0704d510",
			6314 => x"03057908",
			6315 => x"0d058e04",
			6316 => x"00df63f9",
			6317 => x"030b63f9",
			6318 => x"0a029e04",
			6319 => x"000d63f9",
			6320 => x"fec363f9",
			6321 => x"01009708",
			6322 => x"0409b304",
			6323 => x"fe6f63f9",
			6324 => x"019763f9",
			6325 => x"02093d04",
			6326 => x"fe4463f9",
			6327 => x"001e63f9",
			6328 => x"03065920",
			6329 => x"0704be10",
			6330 => x"00048a08",
			6331 => x"0304df04",
			6332 => x"029863f9",
			6333 => x"017063f9",
			6334 => x"040da904",
			6335 => x"02c263f9",
			6336 => x"017d63f9",
			6337 => x"040eab08",
			6338 => x"040c6604",
			6339 => x"029363f9",
			6340 => x"031363f9",
			6341 => x"0305c804",
			6342 => x"000063f9",
			6343 => x"fe6463f9",
			6344 => x"0c050510",
			6345 => x"0a02c108",
			6346 => x"040c5e04",
			6347 => x"ffeb63f9",
			6348 => x"033a63f9",
			6349 => x"0f089c04",
			6350 => x"fe3b63f9",
			6351 => x"016163f9",
			6352 => x"02fc63f9",
			6353 => x"07057730",
			6354 => x"0f07c708",
			6355 => x"0d061d04",
			6356 => x"ff7a63f9",
			6357 => x"fe4363f9",
			6358 => x"0100bc1c",
			6359 => x"0a02db10",
			6360 => x"0c04ed08",
			6361 => x"09010f04",
			6362 => x"009b63f9",
			6363 => x"fe7863f9",
			6364 => x"07051c04",
			6365 => x"000163f9",
			6366 => x"029563f9",
			6367 => x"0d06c708",
			6368 => x"0c054804",
			6369 => x"fe5163f9",
			6370 => x"005b63f9",
			6371 => x"00fc63f9",
			6372 => x"0c052804",
			6373 => x"fe3163f9",
			6374 => x"0f08bf04",
			6375 => x"fe7163f9",
			6376 => x"014063f9",
			6377 => x"0803260c",
			6378 => x"07058b08",
			6379 => x"0c054604",
			6380 => x"000063f9",
			6381 => x"fe9163f9",
			6382 => x"fe3263f9",
			6383 => x"040e6318",
			6384 => x"0803560c",
			6385 => x"09015a04",
			6386 => x"032963f9",
			6387 => x"0c06de04",
			6388 => x"fe6763f9",
			6389 => x"00f963f9",
			6390 => x"0803a008",
			6391 => x"040d6e04",
			6392 => x"01b963f9",
			6393 => x"fe2563f9",
			6394 => x"049063f9",
			6395 => x"0100e304",
			6396 => x"fe3163f9",
			6397 => x"000763f9",
			6398 => x"05060888",
			6399 => x"0100361c",
			6400 => x"06013910",
			6401 => x"09005508",
			6402 => x"02071704",
			6403 => x"ff3065e5",
			6404 => x"fe1d65e5",
			6405 => x"02087c04",
			6406 => x"00aa65e5",
			6407 => x"fe6265e5",
			6408 => x"0d050d08",
			6409 => x"07047a04",
			6410 => x"ff9a65e5",
			6411 => x"051965e5",
			6412 => x"fe2e65e5",
			6413 => x"0e04f034",
			6414 => x"0e047814",
			6415 => x"06010604",
			6416 => x"fe3b65e5",
			6417 => x"0704a708",
			6418 => x"0304af04",
			6419 => x"043d65e5",
			6420 => x"034265e5",
			6421 => x"06012d04",
			6422 => x"050c65e5",
			6423 => x"044865e5",
			6424 => x"02086210",
			6425 => x"0d058308",
			6426 => x"0a027204",
			6427 => x"02f965e5",
			6428 => x"018865e5",
			6429 => x"0f069004",
			6430 => x"01db65e5",
			6431 => x"04ac65e5",
			6432 => x"0704a708",
			6433 => x"0a02bf04",
			6434 => x"023865e5",
			6435 => x"048465e5",
			6436 => x"0d05b604",
			6437 => x"04cd65e5",
			6438 => x"fe3565e5",
			6439 => x"02086c1c",
			6440 => x"0a02a110",
			6441 => x"06013608",
			6442 => x"06011504",
			6443 => x"fe3965e5",
			6444 => x"01e565e5",
			6445 => x"06015604",
			6446 => x"ff7b65e5",
			6447 => x"025c65e5",
			6448 => x"0900aa04",
			6449 => x"004b65e5",
			6450 => x"02085904",
			6451 => x"059965e5",
			6452 => x"03a065e5",
			6453 => x"06017310",
			6454 => x"0c04d408",
			6455 => x"0e054404",
			6456 => x"035365e5",
			6457 => x"016f65e5",
			6458 => x"0a028b04",
			6459 => x"01d265e5",
			6460 => x"04a865e5",
			6461 => x"07051b08",
			6462 => x"03062104",
			6463 => x"000065e5",
			6464 => x"fe4f65e5",
			6465 => x"032265e5",
			6466 => x"07057744",
			6467 => x"0f07960c",
			6468 => x"0f071104",
			6469 => x"fe3a65e5",
			6470 => x"0f076d04",
			6471 => x"ff9465e5",
			6472 => x"fe6065e5",
			6473 => x"06016f18",
			6474 => x"0d06870c",
			6475 => x"0803b408",
			6476 => x"07053204",
			6477 => x"02ec65e5",
			6478 => x"052b65e5",
			6479 => x"fe8065e5",
			6480 => x"0f08b108",
			6481 => x"06016b04",
			6482 => x"fe3565e5",
			6483 => x"000065e5",
			6484 => x"01a165e5",
			6485 => x"07052f10",
			6486 => x"01009508",
			6487 => x"0e064304",
			6488 => x"fe9c65e5",
			6489 => x"035265e5",
			6490 => x"0100a604",
			6491 => x"ff0365e5",
			6492 => x"fe1865e5",
			6493 => x"0209b708",
			6494 => x"0100ad04",
			6495 => x"050265e5",
			6496 => x"014565e5",
			6497 => x"0f08e604",
			6498 => x"fe5265e5",
			6499 => x"007f65e5",
			6500 => x"09026b24",
			6501 => x"0803260c",
			6502 => x"0c054608",
			6503 => x"02098104",
			6504 => x"fe4865e5",
			6505 => x"00cb65e5",
			6506 => x"fe1a65e5",
			6507 => x"0803dc10",
			6508 => x"08035608",
			6509 => x"09015a04",
			6510 => x"04d365e5",
			6511 => x"fe5965e5",
			6512 => x"0100e804",
			6513 => x"ff7765e5",
			6514 => x"028765e5",
			6515 => x"0a031504",
			6516 => x"ff0265e5",
			6517 => x"fe1965e5",
			6518 => x"07072204",
			6519 => x"fe2165e5",
			6520 => x"029065e5",
			6521 => x"040a0120",
			6522 => x"0802c31c",
			6523 => x"0409b314",
			6524 => x"0f06a50c",
			6525 => x"0f063b04",
			6526 => x"fe266751",
			6527 => x"06010304",
			6528 => x"00006751",
			6529 => x"01b36751",
			6530 => x"06011804",
			6531 => x"ff926751",
			6532 => x"fe4a6751",
			6533 => x"06013104",
			6534 => x"01eb6751",
			6535 => x"fe756751",
			6536 => x"fdd66751",
			6537 => x"0802d518",
			6538 => x"0b05a814",
			6539 => x"0d05a710",
			6540 => x"0305890c",
			6541 => x"0d054208",
			6542 => x"0f069604",
			6543 => x"00be6751",
			6544 => x"fd1f6751",
			6545 => x"01ea6751",
			6546 => x"fed66751",
			6547 => x"023f6751",
			6548 => x"fe846751",
			6549 => x"02086c40",
			6550 => x"02086720",
			6551 => x"02086210",
			6552 => x"06013508",
			6553 => x"0c048f04",
			6554 => x"ffe86751",
			6555 => x"006e6751",
			6556 => x"0c047804",
			6557 => x"00426751",
			6558 => x"ffc46751",
			6559 => x"0f06ed08",
			6560 => x"05054a04",
			6561 => x"00006751",
			6562 => x"fc9c6751",
			6563 => x"06014e04",
			6564 => x"01c26751",
			6565 => x"00456751",
			6566 => x"01005a10",
			6567 => x"07049308",
			6568 => x"040c8c04",
			6569 => x"fdf96751",
			6570 => x"01316751",
			6571 => x"0b04bf04",
			6572 => x"029a6751",
			6573 => x"00006751",
			6574 => x"0900a208",
			6575 => x"06014204",
			6576 => x"fc756751",
			6577 => x"fe946751",
			6578 => x"08034804",
			6579 => x"fe6e6751",
			6580 => x"ffd16751",
			6581 => x"06014a20",
			6582 => x"05058210",
			6583 => x"03050008",
			6584 => x"01004304",
			6585 => x"fe716751",
			6586 => x"01606751",
			6587 => x"05051404",
			6588 => x"fdea6751",
			6589 => x"003a6751",
			6590 => x"07050108",
			6591 => x"08031d04",
			6592 => x"00186751",
			6593 => x"01796751",
			6594 => x"0305cc04",
			6595 => x"fd066751",
			6596 => x"00906751",
			6597 => x"0900b510",
			6598 => x"040c9308",
			6599 => x"08038804",
			6600 => x"ffaf6751",
			6601 => x"fde26751",
			6602 => x"09009704",
			6603 => x"ffe66751",
			6604 => x"00e36751",
			6605 => x"0505af08",
			6606 => x"040b9704",
			6607 => x"ff9c6751",
			6608 => x"00f36751",
			6609 => x"01007804",
			6610 => x"ff586751",
			6611 => x"00256751",
			6612 => x"0e061e98",
			6613 => x"0900cd58",
			6614 => x"0b05353c",
			6615 => x"0e059620",
			6616 => x"0900c210",
			6617 => x"0b053108",
			6618 => x"0900a804",
			6619 => x"fffa695d",
			6620 => x"003b695d",
			6621 => x"06014a04",
			6622 => x"018a695d",
			6623 => x"fd57695d",
			6624 => x"040b5d08",
			6625 => x"01007704",
			6626 => x"0072695d",
			6627 => x"fe17695d",
			6628 => x"0f07c704",
			6629 => x"0216695d",
			6630 => x"fe48695d",
			6631 => x"0f07c710",
			6632 => x"0704ee08",
			6633 => x"0003f104",
			6634 => x"ff8c695d",
			6635 => x"fe47695d",
			6636 => x"0b052204",
			6637 => x"ffea695d",
			6638 => x"019e695d",
			6639 => x"0e059d04",
			6640 => x"01dc695d",
			6641 => x"00044604",
			6642 => x"00b9695d",
			6643 => x"ffa4695d",
			6644 => x"040c600c",
			6645 => x"06014e08",
			6646 => x"0d05f704",
			6647 => x"00d0695d",
			6648 => x"ff43695d",
			6649 => x"fcf3695d",
			6650 => x"040cce04",
			6651 => x"0145695d",
			6652 => x"0c04f104",
			6653 => x"fdfd695d",
			6654 => x"01006604",
			6655 => x"ff28695d",
			6656 => x"011b695d",
			6657 => x"00045330",
			6658 => x"0704f114",
			6659 => x"0b051408",
			6660 => x"03062104",
			6661 => x"00eb695d",
			6662 => x"fed6695d",
			6663 => x"01008004",
			6664 => x"0301695d",
			6665 => x"01008604",
			6666 => x"0000695d",
			6667 => x"0273695d",
			6668 => x"08033610",
			6669 => x"02083008",
			6670 => x"0e05f704",
			6671 => x"0191695d",
			6672 => x"0000695d",
			6673 => x"0d060304",
			6674 => x"fdcd695d",
			6675 => x"ff3a695d",
			6676 => x"040bd808",
			6677 => x"06015f04",
			6678 => x"019d695d",
			6679 => x"ff96695d",
			6680 => x"fe39695d",
			6681 => x"0d063f0c",
			6682 => x"06017404",
			6683 => x"01c7695d",
			6684 => x"06017c04",
			6685 => x"000a695d",
			6686 => x"ff69695d",
			6687 => x"fe71695d",
			6688 => x"0f08f93c",
			6689 => x"0c04e720",
			6690 => x"0b04f404",
			6691 => x"014b695d",
			6692 => x"0208ad0c",
			6693 => x"06015a08",
			6694 => x"0f07ce04",
			6695 => x"ff9b695d",
			6696 => x"fe0c695d",
			6697 => x"01a3695d",
			6698 => x"07050508",
			6699 => x"0c04b004",
			6700 => x"ff53695d",
			6701 => x"fdfd695d",
			6702 => x"0900e704",
			6703 => x"007b695d",
			6704 => x"fea1695d",
			6705 => x"03067804",
			6706 => x"020a695d",
			6707 => x"0c04ea08",
			6708 => x"0d064704",
			6709 => x"0180695d",
			6710 => x"feec695d",
			6711 => x"0c04ec08",
			6712 => x"0f088e04",
			6713 => x"fdb0695d",
			6714 => x"0000695d",
			6715 => x"01008404",
			6716 => x"0102695d",
			6717 => x"ff8e695d",
			6718 => x"0308a914",
			6719 => x"09014f0c",
			6720 => x"06019104",
			6721 => x"01f3695d",
			6722 => x"09011b04",
			6723 => x"0000695d",
			6724 => x"0150695d",
			6725 => x"07060004",
			6726 => x"fec2695d",
			6727 => x"00aa695d",
			6728 => x"040ba404",
			6729 => x"fe79695d",
			6730 => x"0100f80c",
			6731 => x"0803c704",
			6732 => x"fe64695d",
			6733 => x"0004f704",
			6734 => x"0000695d",
			6735 => x"ff90695d",
			6736 => x"08037308",
			6737 => x"0f0abc04",
			6738 => x"019b695d",
			6739 => x"ff52695d",
			6740 => x"020bbc04",
			6741 => x"0000695d",
			6742 => x"0183695d",
			6743 => x"040df5b8",
			6744 => x"0505f964",
			6745 => x"0900d33c",
			6746 => x"03061120",
			6747 => x"0900af10",
			6748 => x"0e054b08",
			6749 => x"0900a904",
			6750 => x"00076b41",
			6751 => x"00a96b41",
			6752 => x"0208f204",
			6753 => x"fec46b41",
			6754 => x"00486b41",
			6755 => x"0e057108",
			6756 => x"0b050004",
			6757 => x"003d6b41",
			6758 => x"00f36b41",
			6759 => x"06014204",
			6760 => x"01076b41",
			6761 => x"ffe56b41",
			6762 => x"06015710",
			6763 => x"0505a108",
			6764 => x"0b050004",
			6765 => x"012a6b41",
			6766 => x"03836b41",
			6767 => x"0704ed04",
			6768 => x"fec66b41",
			6769 => x"00416b41",
			6770 => x"01006e04",
			6771 => x"01456b41",
			6772 => x"0c04ec04",
			6773 => x"feac6b41",
			6774 => x"00786b41",
			6775 => x"0e05f714",
			6776 => x"0c04b904",
			6777 => x"04266b41",
			6778 => x"08032508",
			6779 => x"0b053504",
			6780 => x"fe746b41",
			6781 => x"02816b41",
			6782 => x"0c04f104",
			6783 => x"024e6b41",
			6784 => x"007a6b41",
			6785 => x"0c04b004",
			6786 => x"02b06b41",
			6787 => x"0c04e908",
			6788 => x"040c1804",
			6789 => x"fedb6b41",
			6790 => x"010d6b41",
			6791 => x"07050104",
			6792 => x"ff426b41",
			6793 => x"01a86b41",
			6794 => x"08032618",
			6795 => x"09014314",
			6796 => x"0b055204",
			6797 => x"fdb56b41",
			6798 => x"0e065a08",
			6799 => x"040a9504",
			6800 => x"00396b41",
			6801 => x"fdfb6b41",
			6802 => x"0a028704",
			6803 => x"007e6b41",
			6804 => x"fe4b6b41",
			6805 => x"fe676b41",
			6806 => x"0c052820",
			6807 => x"040b8a10",
			6808 => x"0b056308",
			6809 => x"02093a04",
			6810 => x"fe616b41",
			6811 => x"00a66b41",
			6812 => x"0100b004",
			6813 => x"01466b41",
			6814 => x"ff2e6b41",
			6815 => x"0e062e08",
			6816 => x"0b056304",
			6817 => x"ffdb6b41",
			6818 => x"fcd56b41",
			6819 => x"0f085c04",
			6820 => x"015b6b41",
			6821 => x"ff016b41",
			6822 => x"040c2c10",
			6823 => x"0601a708",
			6824 => x"040bc404",
			6825 => x"014f6b41",
			6826 => x"031a6b41",
			6827 => x"0b07b104",
			6828 => x"fea86b41",
			6829 => x"01c66b41",
			6830 => x"08035204",
			6831 => x"fe7c6b41",
			6832 => x"0c054c04",
			6833 => x"ff616b41",
			6834 => x"00d96b41",
			6835 => x"0803d01c",
			6836 => x"0100470c",
			6837 => x"040eab08",
			6838 => x"09004f04",
			6839 => x"ff746b41",
			6840 => x"01886b41",
			6841 => x"fea36b41",
			6842 => x"0f075504",
			6843 => x"fbac6b41",
			6844 => x"06016808",
			6845 => x"0a02dd04",
			6846 => x"ff586b41",
			6847 => x"00e86b41",
			6848 => x"fe5f6b41",
			6849 => x"04112a1c",
			6850 => x"0c047b08",
			6851 => x"0c047404",
			6852 => x"013a6b41",
			6853 => x"fe5e6b41",
			6854 => x"0b04b004",
			6855 => x"019c6b41",
			6856 => x"020a8608",
			6857 => x"02092004",
			6858 => x"00006b41",
			6859 => x"fe466b41",
			6860 => x"040fc604",
			6861 => x"01ac6b41",
			6862 => x"ff4b6b41",
			6863 => x"fe8f6b41",
			6864 => x"08033488",
			6865 => x"00042954",
			6866 => x"06015638",
			6867 => x"0100791c",
			6868 => x"06014610",
			6869 => x"0b051408",
			6870 => x"01006c04",
			6871 => x"00166d7d",
			6872 => x"ff8d6d7d",
			6873 => x"01007504",
			6874 => x"01d26d7d",
			6875 => x"ffca6d7d",
			6876 => x"0003dd04",
			6877 => x"03d06d7d",
			6878 => x"00041d04",
			6879 => x"009c6d7d",
			6880 => x"fe136d7d",
			6881 => x"06014210",
			6882 => x"01007e08",
			6883 => x"0505b104",
			6884 => x"fdd86d7d",
			6885 => x"ffe66d7d",
			6886 => x"0b053504",
			6887 => x"02466d7d",
			6888 => x"ffab6d7d",
			6889 => x"040b5d08",
			6890 => x"07051b04",
			6891 => x"fe6c6d7d",
			6892 => x"00186d7d",
			6893 => x"00336d7d",
			6894 => x"0802eb04",
			6895 => x"fe626d7d",
			6896 => x"0f07c008",
			6897 => x"040ad504",
			6898 => x"00fe6d7d",
			6899 => x"028a6d7d",
			6900 => x"0802ee08",
			6901 => x"0003aa04",
			6902 => x"00006d7d",
			6903 => x"07c36d7d",
			6904 => x"0e061e04",
			6905 => x"fef26d7d",
			6906 => x"008d6d7d",
			6907 => x"07047b14",
			6908 => x"0304be08",
			6909 => x"08032b04",
			6910 => x"00006d7d",
			6911 => x"01326d7d",
			6912 => x"05050108",
			6913 => x"0c044004",
			6914 => x"00006d7d",
			6915 => x"00e16d7d",
			6916 => x"fd4c6d7d",
			6917 => x"02082410",
			6918 => x"08032c08",
			6919 => x"05052004",
			6920 => x"01936d7d",
			6921 => x"ff376d7d",
			6922 => x"0f06c104",
			6923 => x"01e66d7d",
			6924 => x"02db6d7d",
			6925 => x"0100630c",
			6926 => x"08032904",
			6927 => x"021b6d7d",
			6928 => x"0704bf04",
			6929 => x"ff756d7d",
			6930 => x"00c36d7d",
			6931 => x"fdf96d7d",
			6932 => x"03049f4c",
			6933 => x"040c7220",
			6934 => x"0a02b014",
			6935 => x"0f060a08",
			6936 => x"0e039704",
			6937 => x"01786d7d",
			6938 => x"fe786d7d",
			6939 => x"0504e704",
			6940 => x"00076d7d",
			6941 => x"0a028304",
			6942 => x"00006d7d",
			6943 => x"01796d7d",
			6944 => x"0e03e708",
			6945 => x"05050004",
			6946 => x"01426d7d",
			6947 => x"fd776d7d",
			6948 => x"019d6d7d",
			6949 => x"0004920c",
			6950 => x"0b049008",
			6951 => x"03046f04",
			6952 => x"00796d7d",
			6953 => x"fcd26d7d",
			6954 => x"002f6d7d",
			6955 => x"01003f10",
			6956 => x"0f05e608",
			6957 => x"040eab04",
			6958 => x"01986d7d",
			6959 => x"ff176d7d",
			6960 => x"0f06bb04",
			6961 => x"fe936d7d",
			6962 => x"01956d7d",
			6963 => x"040da908",
			6964 => x"05050304",
			6965 => x"01c76d7d",
			6966 => x"00486d7d",
			6967 => x"0803d004",
			6968 => x"fe9a6d7d",
			6969 => x"007b6d7d",
			6970 => x"0f066d0c",
			6971 => x"0c049c08",
			6972 => x"0c047704",
			6973 => x"feef6d7d",
			6974 => x"fd896d7d",
			6975 => x"00ad6d7d",
			6976 => x"0304b720",
			6977 => x"01004110",
			6978 => x"05050f08",
			6979 => x"0504e204",
			6980 => x"00846d7d",
			6981 => x"fe396d7d",
			6982 => x"0b060b04",
			6983 => x"01096d7d",
			6984 => x"00006d7d",
			6985 => x"0207f808",
			6986 => x"0c047304",
			6987 => x"002c6d7d",
			6988 => x"01e56d7d",
			6989 => x"01004904",
			6990 => x"01466d7d",
			6991 => x"ff236d7d",
			6992 => x"0f06ed10",
			6993 => x"0e047808",
			6994 => x"00043204",
			6995 => x"fdfb6d7d",
			6996 => x"ffe66d7d",
			6997 => x"0c04b304",
			6998 => x"fedc6d7d",
			6999 => x"00cb6d7d",
			7000 => x"0e04bb08",
			7001 => x"0704a704",
			7002 => x"ffeb6d7d",
			7003 => x"00a16d7d",
			7004 => x"0f073304",
			7005 => x"ff446d7d",
			7006 => x"ffea6d7d",
			7007 => x"0505b1ac",
			7008 => x"0c04ac4c",
			7009 => x"0c049830",
			7010 => x"0900be20",
			7011 => x"0704d310",
			7012 => x"0704c108",
			7013 => x"0704ad04",
			7014 => x"00136fb1",
			7015 => x"ffae6fb1",
			7016 => x"0c049504",
			7017 => x"00416fb1",
			7018 => x"01ab6fb1",
			7019 => x"0505a008",
			7020 => x"06014204",
			7021 => x"ffeb6fb1",
			7022 => x"fee36fb1",
			7023 => x"00045804",
			7024 => x"02206fb1",
			7025 => x"00006fb1",
			7026 => x"06014504",
			7027 => x"fe916fb1",
			7028 => x"0e05b304",
			7029 => x"02a96fb1",
			7030 => x"0d05b504",
			7031 => x"ff416fb1",
			7032 => x"01e36fb1",
			7033 => x"0704ac0c",
			7034 => x"0207fa04",
			7035 => x"00006fb1",
			7036 => x"040c0c04",
			7037 => x"fe386fb1",
			7038 => x"fd1d6fb1",
			7039 => x"0e05520c",
			7040 => x"0f074908",
			7041 => x"01006604",
			7042 => x"00056fb1",
			7043 => x"fdef6fb1",
			7044 => x"01ec6fb1",
			7045 => x"fe0d6fb1",
			7046 => x"0c04b428",
			7047 => x"07049208",
			7048 => x"040bf104",
			7049 => x"fdba6fb1",
			7050 => x"ff9e6fb1",
			7051 => x"0b04ce10",
			7052 => x"0b04c008",
			7053 => x"0704a604",
			7054 => x"01b26fb1",
			7055 => x"005a6fb1",
			7056 => x"02089304",
			7057 => x"01f56fb1",
			7058 => x"00476fb1",
			7059 => x"0a028008",
			7060 => x"040ae804",
			7061 => x"00156fb1",
			7062 => x"01066fb1",
			7063 => x"02088504",
			7064 => x"ff926fb1",
			7065 => x"00766fb1",
			7066 => x"0c04b618",
			7067 => x"0b04c208",
			7068 => x"05055704",
			7069 => x"ff216fb1",
			7070 => x"02b86fb1",
			7071 => x"05059108",
			7072 => x"00047504",
			7073 => x"fd9f6fb1",
			7074 => x"ff0d6fb1",
			7075 => x"0704da04",
			7076 => x"011f6fb1",
			7077 => x"fe436fb1",
			7078 => x"0c04cd10",
			7079 => x"0704d608",
			7080 => x"040b4204",
			7081 => x"fe076fb1",
			7082 => x"00296fb1",
			7083 => x"0900bc04",
			7084 => x"02096fb1",
			7085 => x"00006fb1",
			7086 => x"06014d08",
			7087 => x"0f070504",
			7088 => x"007d6fb1",
			7089 => x"ff266fb1",
			7090 => x"0a028e04",
			7091 => x"01da6fb1",
			7092 => x"000c6fb1",
			7093 => x"0704eb20",
			7094 => x"0c04e71c",
			7095 => x"040b1508",
			7096 => x"00039e04",
			7097 => x"ff706fb1",
			7098 => x"fdbd6fb1",
			7099 => x"0b052008",
			7100 => x"0900c804",
			7101 => x"018e6fb1",
			7102 => x"ff636fb1",
			7103 => x"0900d908",
			7104 => x"0900c004",
			7105 => x"fd1d6fb1",
			7106 => x"fe356fb1",
			7107 => x"00346fb1",
			7108 => x"00ac6fb1",
			7109 => x"0f080520",
			7110 => x"0d05c304",
			7111 => x"fe406fb1",
			7112 => x"040c930c",
			7113 => x"0f07fe08",
			7114 => x"040c1804",
			7115 => x"00216fb1",
			7116 => x"011d6fb1",
			7117 => x"021b6fb1",
			7118 => x"0900c208",
			7119 => x"06015e04",
			7120 => x"fe006fb1",
			7121 => x"01356fb1",
			7122 => x"06016704",
			7123 => x"f9566fb1",
			7124 => x"ff2c6fb1",
			7125 => x"0e05f714",
			7126 => x"06016c0c",
			7127 => x"0900d908",
			7128 => x"0b054304",
			7129 => x"fd286fb1",
			7130 => x"ff9d6fb1",
			7131 => x"010d6fb1",
			7132 => x"06017304",
			7133 => x"01796fb1",
			7134 => x"00006fb1",
			7135 => x"0208d60c",
			7136 => x"0d061104",
			7137 => x"ffdd6fb1",
			7138 => x"06016704",
			7139 => x"fe2a6fb1",
			7140 => x"ffef6fb1",
			7141 => x"06015b08",
			7142 => x"0c04ea04",
			7143 => x"01d56fb1",
			7144 => x"00196fb1",
			7145 => x"07050404",
			7146 => x"feb96fb1",
			7147 => x"00076fb1",
			7148 => x"0c04d1a0",
			7149 => x"07050470",
			7150 => x"0505b03c",
			7151 => x"0c04d020",
			7152 => x"03060910",
			7153 => x"0305f208",
			7154 => x"0d05cf04",
			7155 => x"000671e5",
			7156 => x"01de71e5",
			7157 => x"0b050304",
			7158 => x"fffd71e5",
			7159 => x"feac71e5",
			7160 => x"0c04ac08",
			7161 => x"08036804",
			7162 => x"feb671e5",
			7163 => x"00e071e5",
			7164 => x"0704c004",
			7165 => x"fee271e5",
			7166 => x"013971e5",
			7167 => x"0704d60c",
			7168 => x"0704d208",
			7169 => x"0900a204",
			7170 => x"ff9671e5",
			7171 => x"01bb71e5",
			7172 => x"fe5a71e5",
			7173 => x"0a02bb08",
			7174 => x"0704ee04",
			7175 => x"023671e5",
			7176 => x"008f71e5",
			7177 => x"0208f204",
			7178 => x"016071e5",
			7179 => x"ff8d71e5",
			7180 => x"0900d620",
			7181 => x"0b052010",
			7182 => x"0c04ca08",
			7183 => x"0704da04",
			7184 => x"fe7371e5",
			7185 => x"000071e5",
			7186 => x"0704ed04",
			7187 => x"021771e5",
			7188 => x"ff0071e5",
			7189 => x"06014608",
			7190 => x"040ad504",
			7191 => x"ff2a71e5",
			7192 => x"00f171e5",
			7193 => x"040c5804",
			7194 => x"fe5371e5",
			7195 => x"fffa71e5",
			7196 => x"0c04af04",
			7197 => x"020f71e5",
			7198 => x"0e061e08",
			7199 => x"0208c004",
			7200 => x"fff071e5",
			7201 => x"020371e5",
			7202 => x"02090004",
			7203 => x"fe9671e5",
			7204 => x"00be71e5",
			7205 => x"08037c28",
			7206 => x"0505db0c",
			7207 => x"02085204",
			7208 => x"ff6671e5",
			7209 => x"08036f04",
			7210 => x"021e71e5",
			7211 => x"00f071e5",
			7212 => x"0d064510",
			7213 => x"06016308",
			7214 => x"0208ab04",
			7215 => x"ff3771e5",
			7216 => x"01e571e5",
			7217 => x"040b1604",
			7218 => x"00ac71e5",
			7219 => x"fe2271e5",
			7220 => x"09010f08",
			7221 => x"02091904",
			7222 => x"00c671e5",
			7223 => x"020c71e5",
			7224 => x"ffcc71e5",
			7225 => x"08038d04",
			7226 => x"fdc471e5",
			7227 => x"009f71e5",
			7228 => x"0c04d21c",
			7229 => x"0505df14",
			7230 => x"0b04f004",
			7231 => x"003371e5",
			7232 => x"0a02bb0c",
			7233 => x"01008008",
			7234 => x"02085b04",
			7235 => x"ff2b71e5",
			7236 => x"fdba71e5",
			7237 => x"ff9f71e5",
			7238 => x"ff9671e5",
			7239 => x"0e067104",
			7240 => x"01cf71e5",
			7241 => x"fef971e5",
			7242 => x"0c04ea28",
			7243 => x"0c04e918",
			7244 => x"07050810",
			7245 => x"0e051608",
			7246 => x"01006b04",
			7247 => x"003071e5",
			7248 => x"021671e5",
			7249 => x"0e055204",
			7250 => x"fdc971e5",
			7251 => x"004a71e5",
			7252 => x"08036c04",
			7253 => x"fdc571e5",
			7254 => x"008b71e5",
			7255 => x"01007904",
			7256 => x"022971e5",
			7257 => x"0e062e04",
			7258 => x"ffe771e5",
			7259 => x"0a029904",
			7260 => x"01ee71e5",
			7261 => x"000071e5",
			7262 => x"0601561c",
			7263 => x"040c440c",
			7264 => x"08035a08",
			7265 => x"0d05ed04",
			7266 => x"000071e5",
			7267 => x"fe6571e5",
			7268 => x"fdaa71e5",
			7269 => x"0d061108",
			7270 => x"01005904",
			7271 => x"000071e5",
			7272 => x"01b071e5",
			7273 => x"06015204",
			7274 => x"ff6071e5",
			7275 => x"000071e5",
			7276 => x"02085b0c",
			7277 => x"0d062a08",
			7278 => x"0b058304",
			7279 => x"01d571e5",
			7280 => x"000071e5",
			7281 => x"000071e5",
			7282 => x"0900b108",
			7283 => x"0416b604",
			7284 => x"019571e5",
			7285 => x"000071e5",
			7286 => x"0d05dc04",
			7287 => x"ff0371e5",
			7288 => x"fffb71e5",
			7289 => x"09007b78",
			7290 => x"0c04913c",
			7291 => x"0c048f38",
			7292 => x"040d6e1c",
			7293 => x"0e03e70c",
			7294 => x"0b049108",
			7295 => x"0f069f04",
			7296 => x"fffb7441",
			7297 => x"01df7441",
			7298 => x"01a47441",
			7299 => x"0f06b208",
			7300 => x"00047004",
			7301 => x"ffa07441",
			7302 => x"fea27441",
			7303 => x"0c047a04",
			7304 => x"001d7441",
			7305 => x"fdb87441",
			7306 => x"0a02ed10",
			7307 => x"03040508",
			7308 => x"0303f504",
			7309 => x"00007441",
			7310 => x"f6b17441",
			7311 => x"0004b804",
			7312 => x"00007441",
			7313 => x"fe197441",
			7314 => x"0a02f304",
			7315 => x"01a07441",
			7316 => x"0e033e04",
			7317 => x"fec07441",
			7318 => x"00007441",
			7319 => x"01b97441",
			7320 => x"0304d82c",
			7321 => x"01004514",
			7322 => x"0f06ca0c",
			7323 => x"01003908",
			7324 => x"0e038e04",
			7325 => x"ffa27441",
			7326 => x"00047441",
			7327 => x"01be7441",
			7328 => x"0f06de04",
			7329 => x"fedc7441",
			7330 => x"00877441",
			7331 => x"0d052610",
			7332 => x"09007508",
			7333 => x"0d051904",
			7334 => x"febb7441",
			7335 => x"fcc87441",
			7336 => x"0b049004",
			7337 => x"feca7441",
			7338 => x"01737441",
			7339 => x"05052d04",
			7340 => x"01cc7441",
			7341 => x"fe207441",
			7342 => x"0c049504",
			7343 => x"fccc7441",
			7344 => x"0e047108",
			7345 => x"0f06ed04",
			7346 => x"00007441",
			7347 => x"01237441",
			7348 => x"fe277441",
			7349 => x"03053348",
			7350 => x"03052f34",
			7351 => x"03052b20",
			7352 => x"09009b10",
			7353 => x"01005c08",
			7354 => x"07047b04",
			7355 => x"ff677441",
			7356 => x"00387441",
			7357 => x"0704ac04",
			7358 => x"00ac7441",
			7359 => x"fefe7441",
			7360 => x"01006408",
			7361 => x"05057504",
			7362 => x"01c77441",
			7363 => x"ff617441",
			7364 => x"0900a204",
			7365 => x"ff3e7441",
			7366 => x"01db7441",
			7367 => x"0601410c",
			7368 => x"0c049608",
			7369 => x"0c048f04",
			7370 => x"ff9b7441",
			7371 => x"01957441",
			7372 => x"fe847441",
			7373 => x"0f073304",
			7374 => x"fdd87441",
			7375 => x"fee17441",
			7376 => x"0b04c20c",
			7377 => x"0704a504",
			7378 => x"010a7441",
			7379 => x"0e04a504",
			7380 => x"01307441",
			7381 => x"027f7441",
			7382 => x"0d056904",
			7383 => x"ffdc7441",
			7384 => x"017d7441",
			7385 => x"09009330",
			7386 => x"0f071f14",
			7387 => x"0f06e308",
			7388 => x"040b0904",
			7389 => x"fea67441",
			7390 => x"007c7441",
			7391 => x"0704bf08",
			7392 => x"0a029d04",
			7393 => x"fe497441",
			7394 => x"ff507441",
			7395 => x"fd4f7441",
			7396 => x"05055710",
			7397 => x"0c047608",
			7398 => x"03054f04",
			7399 => x"fd907441",
			7400 => x"ff8f7441",
			7401 => x"0c049804",
			7402 => x"00417441",
			7403 => x"fea07441",
			7404 => x"09008d04",
			7405 => x"ffe47441",
			7406 => x"0e04f904",
			7407 => x"02687441",
			7408 => x"00b17441",
			7409 => x"0c04b120",
			7410 => x"0c04af10",
			7411 => x"0c04ae08",
			7412 => x"0900cf04",
			7413 => x"ffcc7441",
			7414 => x"01a17441",
			7415 => x"0704db04",
			7416 => x"010c7441",
			7417 => x"ffe87441",
			7418 => x"0d05a908",
			7419 => x"0704d304",
			7420 => x"ff1a7441",
			7421 => x"00787441",
			7422 => x"0704ec04",
			7423 => x"fdf97441",
			7424 => x"ff7b7441",
			7425 => x"0704c310",
			7426 => x"0704be08",
			7427 => x"0b04be04",
			7428 => x"023b7441",
			7429 => x"ffd37441",
			7430 => x"0c04b404",
			7431 => x"015a7441",
			7432 => x"00617441",
			7433 => x"0900ad08",
			7434 => x"01006204",
			7435 => x"00607441",
			7436 => x"ff467441",
			7437 => x"01006804",
			7438 => x"02727441",
			7439 => x"000c7441",
			7440 => x"0c0479c0",
			7441 => x"09008c6c",
			7442 => x"0305003c",
			7443 => x"09007e20",
			7444 => x"01004b10",
			7445 => x"06011c08",
			7446 => x"0b048d04",
			7447 => x"fe0376c5",
			7448 => x"00f376c5",
			7449 => x"01003f04",
			7450 => x"ffa476c5",
			7451 => x"005e76c5",
			7452 => x"0b049108",
			7453 => x"05051104",
			7454 => x"fd9c76c5",
			7455 => x"ffd976c5",
			7456 => x"07049204",
			7457 => x"01e876c5",
			7458 => x"ffae76c5",
			7459 => x"040b690c",
			7460 => x"0e045308",
			7461 => x"0304c704",
			7462 => x"01cb76c5",
			7463 => x"ffb076c5",
			7464 => x"fe5876c5",
			7465 => x"0a029608",
			7466 => x"0b048e04",
			7467 => x"ffa376c5",
			7468 => x"01d876c5",
			7469 => x"00048604",
			7470 => x"ff5976c5",
			7471 => x"019576c5",
			7472 => x"02085214",
			7473 => x"0601350c",
			7474 => x"01005004",
			7475 => x"fd6e76c5",
			7476 => x"02081b04",
			7477 => x"feff76c5",
			7478 => x"014b76c5",
			7479 => x"07049204",
			7480 => x"fea576c5",
			7481 => x"fdb676c5",
			7482 => x"0a029e10",
			7483 => x"03053908",
			7484 => x"05051f04",
			7485 => x"ff9e76c5",
			7486 => x"020476c5",
			7487 => x"040c0a04",
			7488 => x"fdff76c5",
			7489 => x"01c876c5",
			7490 => x"0a02be08",
			7491 => x"0c047504",
			7492 => x"fe1376c5",
			7493 => x"ff7c76c5",
			7494 => x"015876c5",
			7495 => x"05052d18",
			7496 => x"0b04ae10",
			7497 => x"0c04780c",
			7498 => x"0e04b408",
			7499 => x"02084404",
			7500 => x"027376c5",
			7501 => x"016a76c5",
			7502 => x"001176c5",
			7503 => x"ff1476c5",
			7504 => x"09009504",
			7505 => x"017b76c5",
			7506 => x"037276c5",
			7507 => x"0a027820",
			7508 => x"040ae810",
			7509 => x"0a025308",
			7510 => x"040a8804",
			7511 => x"ffd076c5",
			7512 => x"01eb76c5",
			7513 => x"0c047604",
			7514 => x"ff7276c5",
			7515 => x"fe2976c5",
			7516 => x"01005e08",
			7517 => x"03054804",
			7518 => x"019876c5",
			7519 => x"ff0276c5",
			7520 => x"05056604",
			7521 => x"035776c5",
			7522 => x"00c776c5",
			7523 => x"0c04730c",
			7524 => x"05055508",
			7525 => x"08034f04",
			7526 => x"fff776c5",
			7527 => x"fdc776c5",
			7528 => x"013276c5",
			7529 => x"01005e08",
			7530 => x"0a028204",
			7531 => x"ff3876c5",
			7532 => x"014176c5",
			7533 => x"0e04a904",
			7534 => x"fd5976c5",
			7535 => x"001e76c5",
			7536 => x"0c048f3c",
			7537 => x"040b9114",
			7538 => x"01005c0c",
			7539 => x"07049304",
			7540 => x"fea076c5",
			7541 => x"0704aa04",
			7542 => x"00aa76c5",
			7543 => x"027176c5",
			7544 => x"0c047b04",
			7545 => x"004476c5",
			7546 => x"fde976c5",
			7547 => x"0004a018",
			7548 => x"0e04960c",
			7549 => x"0207bc04",
			7550 => x"fd1676c5",
			7551 => x"08036f04",
			7552 => x"007676c5",
			7553 => x"fe0976c5",
			7554 => x"02089804",
			7555 => x"fd7e76c5",
			7556 => x"0e050704",
			7557 => x"00ca76c5",
			7558 => x"fea176c5",
			7559 => x"08039904",
			7560 => x"01b276c5",
			7561 => x"0207eb08",
			7562 => x"09002d04",
			7563 => x"000076c5",
			7564 => x"019c76c5",
			7565 => x"fe7f76c5",
			7566 => x"05050008",
			7567 => x"00053e04",
			7568 => x"01b876c5",
			7569 => x"000076c5",
			7570 => x"0704ed20",
			7571 => x"0704da10",
			7572 => x"0704d708",
			7573 => x"0704c404",
			7574 => x"001176c5",
			7575 => x"ff9476c5",
			7576 => x"0704d904",
			7577 => x"00b776c5",
			7578 => x"023276c5",
			7579 => x"0b051208",
			7580 => x"00042104",
			7581 => x"ffe276c5",
			7582 => x"fea376c5",
			7583 => x"040c1804",
			7584 => x"000376c5",
			7585 => x"021076c5",
			7586 => x"03066910",
			7587 => x"06015108",
			7588 => x"0900a404",
			7589 => x"fe5376c5",
			7590 => x"001976c5",
			7591 => x"05061604",
			7592 => x"00ca76c5",
			7593 => x"fd4976c5",
			7594 => x"07051808",
			7595 => x"01008c04",
			7596 => x"ffce76c5",
			7597 => x"fe7376c5",
			7598 => x"0e05e904",
			7599 => x"fdf176c5",
			7600 => x"002676c5",
			7601 => x"0a02a090",
			7602 => x"0803616c",
			7603 => x"0208f938",
			7604 => x"0b047f18",
			7605 => x"0b04700c",
			7606 => x"0b046f08",
			7607 => x"0a027704",
			7608 => x"fd607951",
			7609 => x"00eb7951",
			7610 => x"fd907951",
			7611 => x"0802fc04",
			7612 => x"fee27951",
			7613 => x"02084504",
			7614 => x"01d27951",
			7615 => x"005f7951",
			7616 => x"0a028010",
			7617 => x"08032e08",
			7618 => x"01004704",
			7619 => x"febc7951",
			7620 => x"00097951",
			7621 => x"0900af04",
			7622 => x"00567951",
			7623 => x"030a7951",
			7624 => x"02086c08",
			7625 => x"00040b04",
			7626 => x"01ac7951",
			7627 => x"ffa97951",
			7628 => x"08035804",
			7629 => x"ffea7951",
			7630 => x"00ee7951",
			7631 => x"08032014",
			7632 => x"08031e10",
			7633 => x"0b059908",
			7634 => x"01006c04",
			7635 => x"00007951",
			7636 => x"01ac7951",
			7637 => x"040b3604",
			7638 => x"fed27951",
			7639 => x"00567951",
			7640 => x"fdfd7951",
			7641 => x"0a028e10",
			7642 => x"0a027f08",
			7643 => x"08032c04",
			7644 => x"ff617951",
			7645 => x"00007951",
			7646 => x"09012004",
			7647 => x"02847951",
			7648 => x"00007951",
			7649 => x"0a029508",
			7650 => x"040b8504",
			7651 => x"00367951",
			7652 => x"feb17951",
			7653 => x"02093004",
			7654 => x"009e7951",
			7655 => x"01b37951",
			7656 => x"040c4710",
			7657 => x"0a029e08",
			7658 => x"0c047504",
			7659 => x"00467951",
			7660 => x"02507951",
			7661 => x"0304df04",
			7662 => x"02097951",
			7663 => x"ffa77951",
			7664 => x"00047104",
			7665 => x"feac7951",
			7666 => x"0900820c",
			7667 => x"07049108",
			7668 => x"09005d04",
			7669 => x"ffa17951",
			7670 => x"01d97951",
			7671 => x"fee87951",
			7672 => x"01f27951",
			7673 => x"040c4450",
			7674 => x"0004823c",
			7675 => x"08036920",
			7676 => x"08036810",
			7677 => x"040c0a08",
			7678 => x"040be404",
			7679 => x"ffcc7951",
			7680 => x"ff287951",
			7681 => x"0704bf04",
			7682 => x"ff837951",
			7683 => x"00c37951",
			7684 => x"0208ab08",
			7685 => x"0704a604",
			7686 => x"028a7951",
			7687 => x"ffab7951",
			7688 => x"040bde04",
			7689 => x"fef67951",
			7690 => x"02727951",
			7691 => x"040bd80c",
			7692 => x"0c04b104",
			7693 => x"fee57951",
			7694 => x"00045204",
			7695 => x"00007951",
			7696 => x"02247951",
			7697 => x"05053b08",
			7698 => x"08036e04",
			7699 => x"02107951",
			7700 => x"ff2b7951",
			7701 => x"0900c204",
			7702 => x"feb37951",
			7703 => x"ffa87951",
			7704 => x"01005004",
			7705 => x"ff287951",
			7706 => x"040c380c",
			7707 => x"0e056808",
			7708 => x"0a02bc04",
			7709 => x"02737951",
			7710 => x"01737951",
			7711 => x"00007951",
			7712 => x"00167951",
			7713 => x"09009830",
			7714 => x"01005a20",
			7715 => x"01005610",
			7716 => x"00049a08",
			7717 => x"040c9304",
			7718 => x"fff47951",
			7719 => x"fed37951",
			7720 => x"040cc604",
			7721 => x"00b37951",
			7722 => x"ffd17951",
			7723 => x"05052e08",
			7724 => x"05052c04",
			7725 => x"01887951",
			7726 => x"feaa7951",
			7727 => x"0e04b404",
			7728 => x"01a27951",
			7729 => x"00387951",
			7730 => x"0b04df0c",
			7731 => x"0e04f908",
			7732 => x"0f075704",
			7733 => x"fe9d7951",
			7734 => x"01007951",
			7735 => x"fd3a7951",
			7736 => x"01507951",
			7737 => x"0f07871c",
			7738 => x"0f076310",
			7739 => x"040cf508",
			7740 => x"0f075d04",
			7741 => x"00997951",
			7742 => x"fe577951",
			7743 => x"0f074604",
			7744 => x"fdb47951",
			7745 => x"00af7951",
			7746 => x"0a02a904",
			7747 => x"00877951",
			7748 => x"0a02d404",
			7749 => x"02167951",
			7750 => x"00687951",
			7751 => x"00046b0c",
			7752 => x"0b051104",
			7753 => x"02347951",
			7754 => x"0c04ec04",
			7755 => x"fe7b7951",
			7756 => x"007c7951",
			7757 => x"040c6008",
			7758 => x"0704d704",
			7759 => x"fdee7951",
			7760 => x"ff687951",
			7761 => x"0a02c104",
			7762 => x"00d67951",
			7763 => x"ffb97951",
			7764 => x"09008fc4",
			7765 => x"03050d6c",
			7766 => x"0f06ed40",
			7767 => x"0e041620",
			7768 => x"0304af10",
			7769 => x"01005108",
			7770 => x"09007104",
			7771 => x"ffeb7bd5",
			7772 => x"009d7bd5",
			7773 => x"06012504",
			7774 => x"005a7bd5",
			7775 => x"fce97bd5",
			7776 => x"0f06c508",
			7777 => x"0a02b404",
			7778 => x"01df7bd5",
			7779 => x"00267bd5",
			7780 => x"06013e04",
			7781 => x"fe247bd5",
			7782 => x"01717bd5",
			7783 => x"09007710",
			7784 => x"0304af08",
			7785 => x"08038104",
			7786 => x"019e7bd5",
			7787 => x"feed7bd5",
			7788 => x"0f06d004",
			7789 => x"fd787bd5",
			7790 => x"ffa07bd5",
			7791 => x"0f067a08",
			7792 => x"06012104",
			7793 => x"00e87bd5",
			7794 => x"fe647bd5",
			7795 => x"07047b04",
			7796 => x"fe8e7bd5",
			7797 => x"001b7bd5",
			7798 => x"09007b18",
			7799 => x"0304ef0c",
			7800 => x"05052008",
			7801 => x"01004104",
			7802 => x"ff417bd5",
			7803 => x"01367bd5",
			7804 => x"fd3c7bd5",
			7805 => x"0e045304",
			7806 => x"fbce7bd5",
			7807 => x"0f072b04",
			7808 => x"fe1c7bd5",
			7809 => x"00ea7bd5",
			7810 => x"05050304",
			7811 => x"fef27bd5",
			7812 => x"06013e08",
			7813 => x"09007f04",
			7814 => x"00f67bd5",
			7815 => x"02067bd5",
			7816 => x"0e048804",
			7817 => x"01217bd5",
			7818 => x"ff597bd5",
			7819 => x"02088330",
			7820 => x"0b049f14",
			7821 => x"03051708",
			7822 => x"00045204",
			7823 => x"fdb97bd5",
			7824 => x"ffa47bd5",
			7825 => x"07049408",
			7826 => x"0e04a004",
			7827 => x"01cc7bd5",
			7828 => x"fe7e7bd5",
			7829 => x"02ca7bd5",
			7830 => x"05055510",
			7831 => x"0704a608",
			7832 => x"05052b04",
			7833 => x"fcd77bd5",
			7834 => x"fe777bd5",
			7835 => x"0704ab04",
			7836 => x"ffaf7bd5",
			7837 => x"fe6a7bd5",
			7838 => x"09008e08",
			7839 => x"0e04a504",
			7840 => x"00077bd5",
			7841 => x"02b57bd5",
			7842 => x"fe2b7bd5",
			7843 => x"0c047610",
			7844 => x"02089d04",
			7845 => x"00867bd5",
			7846 => x"0208bb04",
			7847 => x"fccf7bd5",
			7848 => x"0e04bb04",
			7849 => x"01ba7bd5",
			7850 => x"fead7bd5",
			7851 => x"00045308",
			7852 => x"08032c04",
			7853 => x"00007bd5",
			7854 => x"029b7bd5",
			7855 => x"0b04af08",
			7856 => x"06013e04",
			7857 => x"ff5b7bd5",
			7858 => x"01a37bd5",
			7859 => x"06014604",
			7860 => x"01237bd5",
			7861 => x"ff017bd5",
			7862 => x"0100550c",
			7863 => x"0b04b908",
			7864 => x"03054304",
			7865 => x"02157bd5",
			7866 => x"fff27bd5",
			7867 => x"030f7bd5",
			7868 => x"0e049634",
			7869 => x"0b04b214",
			7870 => x"00040804",
			7871 => x"01607bd5",
			7872 => x"00045808",
			7873 => x"01005804",
			7874 => x"fffc7bd5",
			7875 => x"fd5e7bd5",
			7876 => x"0e047804",
			7877 => x"02227bd5",
			7878 => x"00207bd5",
			7879 => x"0f06c110",
			7880 => x"03050008",
			7881 => x"0003d504",
			7882 => x"ff037bd5",
			7883 => x"018e7bd5",
			7884 => x"08035e04",
			7885 => x"004f7bd5",
			7886 => x"fd8d7bd5",
			7887 => x"02080908",
			7888 => x"0f06ca04",
			7889 => x"01a07bd5",
			7890 => x"02f97bd5",
			7891 => x"00044204",
			7892 => x"ff527bd5",
			7893 => x"01677bd5",
			7894 => x"02080920",
			7895 => x"06012b10",
			7896 => x"0e04d308",
			7897 => x"0a023e04",
			7898 => x"00007bd5",
			7899 => x"02497bd5",
			7900 => x"0a023304",
			7901 => x"00cd7bd5",
			7902 => x"ff107bd5",
			7903 => x"06014508",
			7904 => x"0305b604",
			7905 => x"ff0c7bd5",
			7906 => x"00887bd5",
			7907 => x"03057904",
			7908 => x"fd667bd5",
			7909 => x"fe757bd5",
			7910 => x"0704c410",
			7911 => x"0704c108",
			7912 => x"02093a04",
			7913 => x"00287bd5",
			7914 => x"fe1c7bd5",
			7915 => x"0704c204",
			7916 => x"01c57bd5",
			7917 => x"00437bd5",
			7918 => x"0b04d008",
			7919 => x"0704d704",
			7920 => x"fe757bd5",
			7921 => x"00007bd5",
			7922 => x"0900b704",
			7923 => x"ffc07bd5",
			7924 => x"00337bd5",
			7925 => x"0e053bcc",
			7926 => x"0f071f70",
			7927 => x"03054340",
			7928 => x"09009920",
			7929 => x"01005c10",
			7930 => x"09009308",
			7931 => x"00041004",
			7932 => x"00657eab",
			7933 => x"fff27eab",
			7934 => x"0704a604",
			7935 => x"ff447eab",
			7936 => x"014d7eab",
			7937 => x"03051008",
			7938 => x"0207c304",
			7939 => x"fe9f7eab",
			7940 => x"008c7eab",
			7941 => x"0704aa04",
			7942 => x"fff87eab",
			7943 => x"fe4a7eab",
			7944 => x"0f06a510",
			7945 => x"0c04b208",
			7946 => x"0f067a04",
			7947 => x"01e97eab",
			7948 => x"ffba7eab",
			7949 => x"0704c004",
			7950 => x"fd567eab",
			7951 => x"ff477eab",
			7952 => x"0f070908",
			7953 => x"0207e504",
			7954 => x"02a97eab",
			7955 => x"009f7eab",
			7956 => x"02085204",
			7957 => x"03937eab",
			7958 => x"01757eab",
			7959 => x"0d05a920",
			7960 => x"0e04e910",
			7961 => x"01006208",
			7962 => x"02084404",
			7963 => x"ffd17eab",
			7964 => x"fdd47eab",
			7965 => x"0f06d604",
			7966 => x"fe107eab",
			7967 => x"00cb7eab",
			7968 => x"0c04b108",
			7969 => x"00040704",
			7970 => x"ffbd7eab",
			7971 => x"fe9f7eab",
			7972 => x"0e051004",
			7973 => x"fdac7eab",
			7974 => x"ff177eab",
			7975 => x"040bcc0c",
			7976 => x"040b1508",
			7977 => x"0505af04",
			7978 => x"00f77eab",
			7979 => x"feef7eab",
			7980 => x"027a7eab",
			7981 => x"ff397eab",
			7982 => x"00044b38",
			7983 => x"0d055a1c",
			7984 => x"0704910c",
			7985 => x"05052d08",
			7986 => x"0c047204",
			7987 => x"fecf7eab",
			7988 => x"023d7eab",
			7989 => x"fe3c7eab",
			7990 => x"040b8a08",
			7991 => x"06013d04",
			7992 => x"01db7eab",
			7993 => x"03f37eab",
			7994 => x"040b9d04",
			7995 => x"ffdd7eab",
			7996 => x"01ab7eab",
			7997 => x"0b04bf0c",
			7998 => x"03057908",
			7999 => x"0d056804",
			8000 => x"fec87eab",
			8001 => x"00bb7eab",
			8002 => x"fd897eab",
			8003 => x"02083808",
			8004 => x"0900ad04",
			8005 => x"feaf7eab",
			8006 => x"002d7eab",
			8007 => x"0704eb04",
			8008 => x"009d7eab",
			8009 => x"02217eab",
			8010 => x"0b05311c",
			8011 => x"09009c0c",
			8012 => x"01006208",
			8013 => x"040bf704",
			8014 => x"fed07eab",
			8015 => x"001d7eab",
			8016 => x"fd3d7eab",
			8017 => x"0704a608",
			8018 => x"0e051604",
			8019 => x"02ca7eab",
			8020 => x"00957eab",
			8021 => x"00045b04",
			8022 => x"ff5b7eab",
			8023 => x"007d7eab",
			8024 => x"07051a04",
			8025 => x"fbf57eab",
			8026 => x"00007eab",
			8027 => x"0900ad38",
			8028 => x"0f07f230",
			8029 => x"06014b1c",
			8030 => x"0f079d10",
			8031 => x"040bb708",
			8032 => x"03057904",
			8033 => x"00787eab",
			8034 => x"fe2c7eab",
			8035 => x"0e054b04",
			8036 => x"010d7eab",
			8037 => x"fe6f7eab",
			8038 => x"0d058d08",
			8039 => x"00043104",
			8040 => x"01757eab",
			8041 => x"ff1c7eab",
			8042 => x"02567eab",
			8043 => x"040c9a0c",
			8044 => x"02088904",
			8045 => x"00a97eab",
			8046 => x"05058504",
			8047 => x"feb47eab",
			8048 => x"fd967eab",
			8049 => x"0e054b04",
			8050 => x"014e7eab",
			8051 => x"ffb87eab",
			8052 => x"0305e104",
			8053 => x"02287eab",
			8054 => x"003c7eab",
			8055 => x"0003ea34",
			8056 => x"0100791c",
			8057 => x"0704d40c",
			8058 => x"02085b08",
			8059 => x"06014104",
			8060 => x"fec67eab",
			8061 => x"01777eab",
			8062 => x"02097eab",
			8063 => x"0704ef08",
			8064 => x"040aa904",
			8065 => x"00e97eab",
			8066 => x"030e7eab",
			8067 => x"0505b104",
			8068 => x"fe647eab",
			8069 => x"01577eab",
			8070 => x"0900cd08",
			8071 => x"0003b304",
			8072 => x"00007eab",
			8073 => x"fe067eab",
			8074 => x"09014308",
			8075 => x"040ad504",
			8076 => x"00187eab",
			8077 => x"022d7eab",
			8078 => x"0601ad04",
			8079 => x"fe737eab",
			8080 => x"00007eab",
			8081 => x"040b3614",
			8082 => x"0c050710",
			8083 => x"0704d708",
			8084 => x"0c04ce04",
			8085 => x"ff217eab",
			8086 => x"024f7eab",
			8087 => x"0c04e704",
			8088 => x"fe3a7eab",
			8089 => x"ff7f7eab",
			8090 => x"02257eab",
			8091 => x"0900c410",
			8092 => x"01006f08",
			8093 => x"0505a304",
			8094 => x"ffd97eab",
			8095 => x"017d7eab",
			8096 => x"0c04b404",
			8097 => x"ffd97eab",
			8098 => x"ff0a7eab",
			8099 => x"03061908",
			8100 => x"040c9a04",
			8101 => x"01547eab",
			8102 => x"fdb37eab",
			8103 => x"040b8504",
			8104 => x"00947eab",
			8105 => x"ffa07eab",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(2753, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(5446, initial_addr_3'length));
	end generate gen_rom_7;

	gen_rom_8: if SELECT_ROM = 8 generate
		bank <= (
			0 => x"00000005",
			1 => x"00000009",
			2 => x"05095e04",
			3 => x"00000015",
			4 => x"fed00015",
			5 => x"040bf104",
			6 => x"fffd0029",
			7 => x"040e2304",
			8 => x"00270029",
			9 => x"00000029",
			10 => x"040c8504",
			11 => x"fffd003d",
			12 => x"040e2304",
			13 => x"000e003d",
			14 => x"0000003d",
			15 => x"08034d08",
			16 => x"0802eb04",
			17 => x"00000051",
			18 => x"000e0051",
			19 => x"00000051",
			20 => x"0b083808",
			21 => x"0901bc04",
			22 => x"00000065",
			23 => x"00010065",
			24 => x"ff540065",
			25 => x"0707640c",
			26 => x"040c5e04",
			27 => x"00000081",
			28 => x"040e2304",
			29 => x"002f0081",
			30 => x"00000081",
			31 => x"ff740081",
			32 => x"0707640c",
			33 => x"040c3e04",
			34 => x"0000009d",
			35 => x"040e2304",
			36 => x"0019009d",
			37 => x"0000009d",
			38 => x"ff9a009d",
			39 => x"0a02880c",
			40 => x"0a027704",
			41 => x"000000c1",
			42 => x"06017d04",
			43 => x"000000c1",
			44 => x"001800c1",
			45 => x"0a02cc04",
			46 => x"ffd900c1",
			47 => x"000000c1",
			48 => x"0101500c",
			49 => x"0a02d108",
			50 => x"0a026504",
			51 => x"000000e5",
			52 => x"ffdf00e5",
			53 => x"000000e5",
			54 => x"0a02a104",
			55 => x"003600e5",
			56 => x"000000e5",
			57 => x"0c06dc0c",
			58 => x"0901bc04",
			59 => x"00000109",
			60 => x"09026b04",
			61 => x"000a0109",
			62 => x"00000109",
			63 => x"0c06e504",
			64 => x"ff560109",
			65 => x"00000109",
			66 => x"0a02880c",
			67 => x"00038504",
			68 => x"00000135",
			69 => x"06017d04",
			70 => x"00000135",
			71 => x"00570135",
			72 => x"06019904",
			73 => x"00000135",
			74 => x"0003cc04",
			75 => x"00000135",
			76 => x"ffdb0135",
			77 => x"08033f0c",
			78 => x"040b6b04",
			79 => x"00000161",
			80 => x"040c9a04",
			81 => x"001a0161",
			82 => x"00000161",
			83 => x"0e0c8c08",
			84 => x"040df504",
			85 => x"ff920161",
			86 => x"00000161",
			87 => x"00000161",
			88 => x"07076410",
			89 => x"0901bc04",
			90 => x"00000185",
			91 => x"040b6b04",
			92 => x"00000185",
			93 => x"0c061404",
			94 => x"00000185",
			95 => x"004a0185",
			96 => x"ff020185",
			97 => x"0509ab10",
			98 => x"0706c904",
			99 => x"000001a9",
			100 => x"05088604",
			101 => x"000001a9",
			102 => x"0b076304",
			103 => x"000001a9",
			104 => x"003101a9",
			105 => x"fffb01a9",
			106 => x"0f0b1704",
			107 => x"000001cd",
			108 => x"0101810c",
			109 => x"06018a04",
			110 => x"000001cd",
			111 => x"030cdd04",
			112 => x"ff9001cd",
			113 => x"000001cd",
			114 => x"000001cd",
			115 => x"0c06dc10",
			116 => x"0901bc04",
			117 => x"000001f9",
			118 => x"0c063004",
			119 => x"000001f9",
			120 => x"09026b04",
			121 => x"002001f9",
			122 => x"000001f9",
			123 => x"0c06e504",
			124 => x"ff4b01f9",
			125 => x"000001f9",
			126 => x"07076414",
			127 => x"040c4708",
			128 => x"01016004",
			129 => x"fff80225",
			130 => x"00000225",
			131 => x"0901bc04",
			132 => x"00000225",
			133 => x"0c063004",
			134 => x"00000225",
			135 => x"00560225",
			136 => x"ff1b0225",
			137 => x"040c470c",
			138 => x"040b1404",
			139 => x"00000259",
			140 => x"0f0be504",
			141 => x"ffec0259",
			142 => x"00000259",
			143 => x"040e230c",
			144 => x"020a2d04",
			145 => x"00000259",
			146 => x"020b0f04",
			147 => x"00330259",
			148 => x"00000259",
			149 => x"00000259",
			150 => x"0b07b514",
			151 => x"05075604",
			152 => x"0000028d",
			153 => x"0a02dd0c",
			154 => x"0a026204",
			155 => x"0000028d",
			156 => x"030ba604",
			157 => x"0053028d",
			158 => x"0000028d",
			159 => x"0000028d",
			160 => x"0d095b04",
			161 => x"0000028d",
			162 => x"ffed028d",
			163 => x"08035e14",
			164 => x"020a9904",
			165 => x"000002c1",
			166 => x"0c061404",
			167 => x"000002c1",
			168 => x"0c06dc08",
			169 => x"00038104",
			170 => x"000002c1",
			171 => x"001c02c1",
			172 => x"000002c1",
			173 => x"020ad104",
			174 => x"000002c1",
			175 => x"ff9f02c1",
			176 => x"07076414",
			177 => x"0c05f604",
			178 => x"000002ed",
			179 => x"0601ca0c",
			180 => x"020a2d04",
			181 => x"000002ed",
			182 => x"06017c04",
			183 => x"000002ed",
			184 => x"001a02ed",
			185 => x"000002ed",
			186 => x"ffd202ed",
			187 => x"040c470c",
			188 => x"06018a04",
			189 => x"00000329",
			190 => x"0f0be504",
			191 => x"ffd90329",
			192 => x"00000329",
			193 => x"0601b210",
			194 => x"05075604",
			195 => x"00000329",
			196 => x"0d091c08",
			197 => x"040e2304",
			198 => x"00510329",
			199 => x"00000329",
			200 => x"00000329",
			201 => x"00000329",
			202 => x"07072814",
			203 => x"0901bc04",
			204 => x"00000365",
			205 => x"020a9904",
			206 => x"00000365",
			207 => x"08036b08",
			208 => x"0c063004",
			209 => x"00000365",
			210 => x"00480365",
			211 => x"00000365",
			212 => x"06019204",
			213 => x"00000365",
			214 => x"0b07c304",
			215 => x"00000365",
			216 => x"ff340365",
			217 => x"07067114",
			218 => x"07061304",
			219 => x"000003a9",
			220 => x"040b8e04",
			221 => x"000003a9",
			222 => x"0a02e408",
			223 => x"0f0af504",
			224 => x"014a03a9",
			225 => x"000003a9",
			226 => x"000003a9",
			227 => x"08034a04",
			228 => x"000003a9",
			229 => x"0e0c8c08",
			230 => x"06019904",
			231 => x"000003a9",
			232 => x"ff6f03a9",
			233 => x"000003a9",
			234 => x"020aad10",
			235 => x"020a2d04",
			236 => x"000003ed",
			237 => x"06019608",
			238 => x"06017c04",
			239 => x"000003ed",
			240 => x"004f03ed",
			241 => x"000003ed",
			242 => x"0802e304",
			243 => x"000003ed",
			244 => x"06018a04",
			245 => x"000003ed",
			246 => x"040b1404",
			247 => x"000003ed",
			248 => x"0a026104",
			249 => x"000003ed",
			250 => x"ffcf03ed",
			251 => x"0901fa0c",
			252 => x"0f0b1008",
			253 => x"040d2e04",
			254 => x"ff770439",
			255 => x"00000439",
			256 => x"00000439",
			257 => x"0f0b2d0c",
			258 => x"0c06ac08",
			259 => x"07069b04",
			260 => x"00000439",
			261 => x"00d10439",
			262 => x"00000439",
			263 => x"040c470c",
			264 => x"09024f08",
			265 => x"040b5d04",
			266 => x"00000439",
			267 => x"ffc40439",
			268 => x"00000439",
			269 => x"00000439",
			270 => x"0a028714",
			271 => x"0a026404",
			272 => x"0000048d",
			273 => x"020a9904",
			274 => x"0000048d",
			275 => x"05091b08",
			276 => x"0c063204",
			277 => x"0000048d",
			278 => x"0113048d",
			279 => x"0000048d",
			280 => x"040d420c",
			281 => x"09024f08",
			282 => x"08030d04",
			283 => x"0000048d",
			284 => x"ffc1048d",
			285 => x"0000048d",
			286 => x"0a02dd08",
			287 => x"0a02bc04",
			288 => x"0000048d",
			289 => x"001c048d",
			290 => x"0000048d",
			291 => x"0601a518",
			292 => x"0d097514",
			293 => x"06017c04",
			294 => x"000004c9",
			295 => x"0d079604",
			296 => x"000004c9",
			297 => x"0a025404",
			298 => x"000004c9",
			299 => x"06019904",
			300 => x"005e04c9",
			301 => x"000004c9",
			302 => x"000004c9",
			303 => x"08032604",
			304 => x"000004c9",
			305 => x"ffff04c9",
			306 => x"08034d18",
			307 => x"040b1604",
			308 => x"00000505",
			309 => x"0c063204",
			310 => x"00000505",
			311 => x"0707280c",
			312 => x"01011504",
			313 => x"00000505",
			314 => x"0802e004",
			315 => x"00000505",
			316 => x"00600505",
			317 => x"00000505",
			318 => x"040d0e04",
			319 => x"ff440505",
			320 => x"00000505",
			321 => x"040df520",
			322 => x"0901dd08",
			323 => x"040d2e04",
			324 => x"ffb90559",
			325 => x"00000559",
			326 => x"06018e08",
			327 => x"09020504",
			328 => x"00000559",
			329 => x"00640559",
			330 => x"040c4708",
			331 => x"09023904",
			332 => x"ffbd0559",
			333 => x"00000559",
			334 => x"09026b04",
			335 => x"001f0559",
			336 => x"00000559",
			337 => x"0a02dd08",
			338 => x"0c05a204",
			339 => x"00000559",
			340 => x"01db0559",
			341 => x"00000559",
			342 => x"040c5e18",
			343 => x"01016014",
			344 => x"0802d804",
			345 => x"000005a5",
			346 => x"0508fd0c",
			347 => x"00037d04",
			348 => x"000005a5",
			349 => x"0b07c304",
			350 => x"ff8205a5",
			351 => x"000005a5",
			352 => x"000005a5",
			353 => x"000005a5",
			354 => x"08036e0c",
			355 => x"01010b04",
			356 => x"000005a5",
			357 => x"00040c04",
			358 => x"000005a5",
			359 => x"006a05a5",
			360 => x"000005a5",
			361 => x"040c4718",
			362 => x"0b078214",
			363 => x"0706e110",
			364 => x"0c06870c",
			365 => x"01016708",
			366 => x"0802d504",
			367 => x"000005f1",
			368 => x"ffad05f1",
			369 => x"000005f1",
			370 => x"000005f1",
			371 => x"000005f1",
			372 => x"000005f1",
			373 => x"08035e0c",
			374 => x"01010b04",
			375 => x"000005f1",
			376 => x"07073c04",
			377 => x"00b705f1",
			378 => x"000005f1",
			379 => x"000005f1",
			380 => x"0508ee1c",
			381 => x"0c063008",
			382 => x"040df504",
			383 => x"ffee0645",
			384 => x"00000645",
			385 => x"08036b10",
			386 => x"0e0b070c",
			387 => x"040b1604",
			388 => x"00000645",
			389 => x"0901bc04",
			390 => x"00000645",
			391 => x"00d80645",
			392 => x"00000645",
			393 => x"00000645",
			394 => x"06018e04",
			395 => x"00000645",
			396 => x"0b07b504",
			397 => x"00000645",
			398 => x"07070b04",
			399 => x"00000645",
			400 => x"ffc50645",
			401 => x"05080f10",
			402 => x"0100e504",
			403 => x"000006a1",
			404 => x"040c9304",
			405 => x"000006a1",
			406 => x"0c05b404",
			407 => x"000006a1",
			408 => x"01a706a1",
			409 => x"01015910",
			410 => x"07068804",
			411 => x"000006a1",
			412 => x"0a026504",
			413 => x"000006a1",
			414 => x"0802e304",
			415 => x"000006a1",
			416 => x"ff9706a1",
			417 => x"0803730c",
			418 => x"0706a104",
			419 => x"000006a1",
			420 => x"00039a04",
			421 => x"000006a1",
			422 => x"005206a1",
			423 => x"000006a1",
			424 => x"0901fa0c",
			425 => x"0f0b1008",
			426 => x"040d2e04",
			427 => x"ff8006fd",
			428 => x"000006fd",
			429 => x"000006fd",
			430 => x"0e0b0714",
			431 => x"0c06ac10",
			432 => x"0601bb0c",
			433 => x"05082e04",
			434 => x"000006fd",
			435 => x"0b071004",
			436 => x"000006fd",
			437 => x"00c406fd",
			438 => x"000006fd",
			439 => x"000006fd",
			440 => x"09024f0c",
			441 => x"0c063304",
			442 => x"000006fd",
			443 => x"07073804",
			444 => x"ffba06fd",
			445 => x"000006fd",
			446 => x"000006fd",
			447 => x"020aad14",
			448 => x"020a2d04",
			449 => x"00000761",
			450 => x"0c05d804",
			451 => x"00000761",
			452 => x"09016b04",
			453 => x"00000761",
			454 => x"0f0a8a04",
			455 => x"01780761",
			456 => x"00000761",
			457 => x"0d09500c",
			458 => x"01015004",
			459 => x"00000761",
			460 => x"08035604",
			461 => x"002f0761",
			462 => x"00000761",
			463 => x"09024f10",
			464 => x"0c068904",
			465 => x"00000761",
			466 => x"030b1304",
			467 => x"00000761",
			468 => x"01015304",
			469 => x"00000761",
			470 => x"ffa80761",
			471 => x"00000761",
			472 => x"0d097520",
			473 => x"0c063008",
			474 => x"040df504",
			475 => x"fff107ad",
			476 => x"000007ad",
			477 => x"040b1604",
			478 => x"000007ad",
			479 => x"08036b10",
			480 => x"0e0b070c",
			481 => x"0c06c208",
			482 => x"01011504",
			483 => x"000007ad",
			484 => x"00cb07ad",
			485 => x"000007ad",
			486 => x"000007ad",
			487 => x"000007ad",
			488 => x"01015f04",
			489 => x"000007ad",
			490 => x"ffd707ad",
			491 => x"0d09501c",
			492 => x"07061304",
			493 => x"000007f9",
			494 => x"06019f14",
			495 => x"09022810",
			496 => x"06017804",
			497 => x"000007f9",
			498 => x"09016b04",
			499 => x"000007f9",
			500 => x"020a1004",
			501 => x"000007f9",
			502 => x"008407f9",
			503 => x"000007f9",
			504 => x"000007f9",
			505 => x"020ad604",
			506 => x"000007f9",
			507 => x"06018d04",
			508 => x"000007f9",
			509 => x"fff207f9",
			510 => x"040d5524",
			511 => x"08034718",
			512 => x"0901dd04",
			513 => x"00000855",
			514 => x"0b07b510",
			515 => x"0e0b070c",
			516 => x"030a3904",
			517 => x"00000855",
			518 => x"0b071004",
			519 => x"00000855",
			520 => x"00a80855",
			521 => x"00000855",
			522 => x"00000855",
			523 => x"040d1b08",
			524 => x"030c2504",
			525 => x"ff880855",
			526 => x"00000855",
			527 => x"00000855",
			528 => x"08039c08",
			529 => x"06019404",
			530 => x"00000855",
			531 => x"01910855",
			532 => x"00000855",
			533 => x"0e0aa21c",
			534 => x"0c063004",
			535 => x"000008a9",
			536 => x"08036b14",
			537 => x"0309c004",
			538 => x"000008a9",
			539 => x"0c06a10c",
			540 => x"020a8304",
			541 => x"000008a9",
			542 => x"0d092204",
			543 => x"00cd08a9",
			544 => x"000008a9",
			545 => x"000008a9",
			546 => x"000008a9",
			547 => x"040b4604",
			548 => x"000008a9",
			549 => x"0a026104",
			550 => x"000008a9",
			551 => x"0f0af304",
			552 => x"000008a9",
			553 => x"ffc608a9",
			554 => x"040d5528",
			555 => x"01015914",
			556 => x"030b2310",
			557 => x"0802d804",
			558 => x"0000090d",
			559 => x"040ce108",
			560 => x"09022b04",
			561 => x"ff7a090d",
			562 => x"0000090d",
			563 => x"0000090d",
			564 => x"0000090d",
			565 => x"0d097510",
			566 => x"0f0c090c",
			567 => x"040b1504",
			568 => x"0000090d",
			569 => x"05084d04",
			570 => x"0000090d",
			571 => x"00c0090d",
			572 => x"0000090d",
			573 => x"0000090d",
			574 => x"0a02dd08",
			575 => x"0100e504",
			576 => x"0000090d",
			577 => x"0264090d",
			578 => x"0000090d",
			579 => x"01013f14",
			580 => x"040d2e04",
			581 => x"ff020981",
			582 => x"0803810c",
			583 => x"00043904",
			584 => x"00000981",
			585 => x"0100eb04",
			586 => x"00000981",
			587 => x"00960981",
			588 => x"00000981",
			589 => x"030b530c",
			590 => x"0c06aa08",
			591 => x"07069b04",
			592 => x"00000981",
			593 => x"00f50981",
			594 => x"00000981",
			595 => x"0c06a410",
			596 => x"0f0b4a04",
			597 => x"00000981",
			598 => x"0a027004",
			599 => x"00000981",
			600 => x"07070e04",
			601 => x"ff6b0981",
			602 => x"00000981",
			603 => x"01018a08",
			604 => x"0c06a704",
			605 => x"00000981",
			606 => x"005c0981",
			607 => x"00000981",
			608 => x"040d552c",
			609 => x"01015918",
			610 => x"0b079510",
			611 => x"0802d804",
			612 => x"000009ed",
			613 => x"0706e208",
			614 => x"08030804",
			615 => x"ff6709ed",
			616 => x"000009ed",
			617 => x"000009ed",
			618 => x"08030604",
			619 => x"001109ed",
			620 => x"000009ed",
			621 => x"0d097510",
			622 => x"0e0b940c",
			623 => x"0508fb08",
			624 => x"0706a104",
			625 => x"000009ed",
			626 => x"00ac09ed",
			627 => x"000009ed",
			628 => x"000009ed",
			629 => x"000009ed",
			630 => x"0a02dd08",
			631 => x"0100e504",
			632 => x"000009ed",
			633 => x"023909ed",
			634 => x"000009ed",
			635 => x"08030f1c",
			636 => x"0b079310",
			637 => x"0101590c",
			638 => x"00039a04",
			639 => x"00000a61",
			640 => x"0003c804",
			641 => x"ffac0a61",
			642 => x"00000a61",
			643 => x"00000a61",
			644 => x"01016608",
			645 => x"09020a04",
			646 => x"00000a61",
			647 => x"00bc0a61",
			648 => x"00000a61",
			649 => x"040c4c08",
			650 => x"09024f04",
			651 => x"ff750a61",
			652 => x"00000a61",
			653 => x"00047d14",
			654 => x"0601c210",
			655 => x"0003f304",
			656 => x"00000a61",
			657 => x"06018a04",
			658 => x"00000a61",
			659 => x"0601b404",
			660 => x"00590a61",
			661 => x"00000a61",
			662 => x"00000a61",
			663 => x"00000a61",
			664 => x"0004a728",
			665 => x"0706e118",
			666 => x"01015914",
			667 => x"0a029310",
			668 => x"0802d804",
			669 => x"00000abd",
			670 => x"0b079508",
			671 => x"00037d04",
			672 => x"00000abd",
			673 => x"ff750abd",
			674 => x"00000abd",
			675 => x"00000abd",
			676 => x"00000abd",
			677 => x"0707280c",
			678 => x"08036808",
			679 => x"06017d04",
			680 => x"00000abd",
			681 => x"00390abd",
			682 => x"00000abd",
			683 => x"00000abd",
			684 => x"0004ab04",
			685 => x"00f70abd",
			686 => x"00000abd",
			687 => x"01013f14",
			688 => x"040d2e04",
			689 => x"ff170b39",
			690 => x"0803810c",
			691 => x"00043904",
			692 => x"00000b39",
			693 => x"0100eb04",
			694 => x"00000b39",
			695 => x"007f0b39",
			696 => x"00000b39",
			697 => x"0e0b0714",
			698 => x"0c06aa10",
			699 => x"07069b04",
			700 => x"00000b39",
			701 => x"0b07b508",
			702 => x"0c063304",
			703 => x"00000b39",
			704 => x"00fc0b39",
			705 => x"00000b39",
			706 => x"00000b39",
			707 => x"0c06a710",
			708 => x"09023f0c",
			709 => x"0a027004",
			710 => x"00000b39",
			711 => x"01016904",
			712 => x"ff610b39",
			713 => x"00000b39",
			714 => x"00000b39",
			715 => x"01018a04",
			716 => x"004e0b39",
			717 => x"00000b39",
			718 => x"040df530",
			719 => x"0601a524",
			720 => x"020ae614",
			721 => x"040d2e10",
			722 => x"0802e304",
			723 => x"00000bad",
			724 => x"01016008",
			725 => x"0f0b0904",
			726 => x"ff870bad",
			727 => x"00000bad",
			728 => x"00000bad",
			729 => x"00000bad",
			730 => x"0d09750c",
			731 => x"01012304",
			732 => x"00000bad",
			733 => x"0f0b9804",
			734 => x"00c00bad",
			735 => x"00000bad",
			736 => x"00000bad",
			737 => x"09023f08",
			738 => x"040cce04",
			739 => x"ff9c0bad",
			740 => x"00000bad",
			741 => x"00000bad",
			742 => x"0a02dd08",
			743 => x"0100e504",
			744 => x"00000bad",
			745 => x"023b0bad",
			746 => x"00000bad",
			747 => x"0c063a10",
			748 => x"05086a0c",
			749 => x"0a02cb04",
			750 => x"fea00c39",
			751 => x"0a02cc04",
			752 => x"00000c39",
			753 => x"ffaf0c39",
			754 => x"00000c39",
			755 => x"09020e14",
			756 => x"020b390c",
			757 => x"030ae508",
			758 => x"06018504",
			759 => x"00000c39",
			760 => x"ff560c39",
			761 => x"00000c39",
			762 => x"0d090104",
			763 => x"00490c39",
			764 => x"00000c39",
			765 => x"0d09500c",
			766 => x"030ba608",
			767 => x"01014d04",
			768 => x"00000c39",
			769 => x"013a0c39",
			770 => x"00000c39",
			771 => x"07070c0c",
			772 => x"030b2a04",
			773 => x"00000c39",
			774 => x"0802ee04",
			775 => x"ff2d0c39",
			776 => x"00000c39",
			777 => x"0601cc08",
			778 => x"0e0ac904",
			779 => x"00000c39",
			780 => x"01280c39",
			781 => x"ffaa0c39",
			782 => x"020a5b0c",
			783 => x"00037d04",
			784 => x"00000cb5",
			785 => x"05086a04",
			786 => x"ff770cb5",
			787 => x"00000cb5",
			788 => x"0e0aa218",
			789 => x"0c06c014",
			790 => x"00048110",
			791 => x"020a8304",
			792 => x"00000cb5",
			793 => x"0100f804",
			794 => x"00000cb5",
			795 => x"0c05d804",
			796 => x"00000cb5",
			797 => x"00830cb5",
			798 => x"00000cb5",
			799 => x"00000cb5",
			800 => x"01016110",
			801 => x"09022a04",
			802 => x"00000cb5",
			803 => x"0f0afc04",
			804 => x"00000cb5",
			805 => x"0003a304",
			806 => x"ff700cb5",
			807 => x"00000cb5",
			808 => x"00043108",
			809 => x"00039504",
			810 => x"00000cb5",
			811 => x"00340cb5",
			812 => x"00000cb5",
			813 => x"0100f804",
			814 => x"febb0d21",
			815 => x"0601a124",
			816 => x"09022a18",
			817 => x"09021210",
			818 => x"0003f30c",
			819 => x"06018504",
			820 => x"00000d21",
			821 => x"030ae504",
			822 => x"ff6c0d21",
			823 => x"00000d21",
			824 => x"00c60d21",
			825 => x"05083e04",
			826 => x"00000d21",
			827 => x"011e0d21",
			828 => x"0a026708",
			829 => x"030b1b04",
			830 => x"00000d21",
			831 => x"fed40d21",
			832 => x"00bd0d21",
			833 => x"07068804",
			834 => x"00000d21",
			835 => x"01015f04",
			836 => x"ff140d21",
			837 => x"08036804",
			838 => x"00580d21",
			839 => x"ffae0d21",
			840 => x"09020524",
			841 => x"0902021c",
			842 => x"09018b04",
			843 => x"fe510dbd",
			844 => x"07067208",
			845 => x"09019004",
			846 => x"ff430dbd",
			847 => x"fe5a0dbd",
			848 => x"0e0a700c",
			849 => x"06018e04",
			850 => x"fe600dbd",
			851 => x"0601a104",
			852 => x"043a0dbd",
			853 => x"ffd80dbd",
			854 => x"fe610dbd",
			855 => x"07068604",
			856 => x"fe640dbd",
			857 => x"02a60dbd",
			858 => x"0706a110",
			859 => x"05086a0c",
			860 => x"0c063204",
			861 => x"fe4e0dbd",
			862 => x"0b071e04",
			863 => x"00600dbd",
			864 => x"fe6a0dbd",
			865 => x"015d0dbd",
			866 => x"08036818",
			867 => x"0a02a910",
			868 => x"0706b408",
			869 => x"0003aa04",
			870 => x"029b0dbd",
			871 => x"01250dbd",
			872 => x"0003f304",
			873 => x"02a00dbd",
			874 => x"03150dbd",
			875 => x"00041404",
			876 => x"00820dbd",
			877 => x"028a0dbd",
			878 => x"fe760dbd",
			879 => x"09018b04",
			880 => x"feff0e31",
			881 => x"040c8524",
			882 => x"06018c0c",
			883 => x"09020504",
			884 => x"00000e31",
			885 => x"0b071004",
			886 => x"00000e31",
			887 => x"009e0e31",
			888 => x"01016010",
			889 => x"0707380c",
			890 => x"040c4408",
			891 => x"0802d804",
			892 => x"00000e31",
			893 => x"ff6a0e31",
			894 => x"00000e31",
			895 => x"00000e31",
			896 => x"08032504",
			897 => x"00090e31",
			898 => x"00000e31",
			899 => x"0a02db10",
			900 => x"0d08f404",
			901 => x"010f0e31",
			902 => x"0d097704",
			903 => x"00000e31",
			904 => x"01015b04",
			905 => x"00000e31",
			906 => x"00670e31",
			907 => x"00000e31",
			908 => x"0101492c",
			909 => x"0901fa18",
			910 => x"01010f04",
			911 => x"fe5e0ec5",
			912 => x"07065a04",
			913 => x"fe630ec5",
			914 => x"0d083104",
			915 => x"02990ec5",
			916 => x"0e09fd08",
			917 => x"0c063404",
			918 => x"fe7a0ec5",
			919 => x"00e80ec5",
			920 => x"fe6b0ec5",
			921 => x"07068604",
			922 => x"fe620ec5",
			923 => x"0e0a8608",
			924 => x"01014504",
			925 => x"02a20ec5",
			926 => x"011d0ec5",
			927 => x"0601a604",
			928 => x"00000ec5",
			929 => x"fe5e0ec5",
			930 => x"0d089a04",
			931 => x"fe760ec5",
			932 => x"08034c14",
			933 => x"0706a104",
			934 => x"004c0ec5",
			935 => x"0c06cb0c",
			936 => x"0b07d608",
			937 => x"0b077104",
			938 => x"017c0ec5",
			939 => x"01d30ec5",
			940 => x"00d30ec5",
			941 => x"00430ec5",
			942 => x"040d2e04",
			943 => x"fec20ec5",
			944 => x"00b10ec5",
			945 => x"09018b04",
			946 => x"feb20f49",
			947 => x"0c06521c",
			948 => x"0a029e0c",
			949 => x"05086a08",
			950 => x"0802d404",
			951 => x"00000f49",
			952 => x"ff080f49",
			953 => x"00000f49",
			954 => x"020b6908",
			955 => x"040c9a04",
			956 => x"00000f49",
			957 => x"00930f49",
			958 => x"08033604",
			959 => x"00000f49",
			960 => x"ffcb0f49",
			961 => x"040b3608",
			962 => x"09020504",
			963 => x"00000f49",
			964 => x"01020f49",
			965 => x"020ae60c",
			966 => x"0706de04",
			967 => x"00000f49",
			968 => x"01016004",
			969 => x"ff300f49",
			970 => x"00000f49",
			971 => x"08036e0c",
			972 => x"00039a04",
			973 => x"00000f49",
			974 => x"01014104",
			975 => x"00000f49",
			976 => x"00f90f49",
			977 => x"ffc00f49",
			978 => x"01014934",
			979 => x"09020e2c",
			980 => x"09020220",
			981 => x"0100f804",
			982 => x"fe3d0fe5",
			983 => x"0c06330c",
			984 => x"09019004",
			985 => x"ffa40fe5",
			986 => x"0901bf04",
			987 => x"fe880fe5",
			988 => x"fe430fe5",
			989 => x"0e09fd08",
			990 => x"020ad604",
			991 => x"fe600fe5",
			992 => x"047f0fe5",
			993 => x"0901fa04",
			994 => x"fe570fe5",
			995 => x"ff5e0fe5",
			996 => x"0c065008",
			997 => x"05082e04",
			998 => x"fe430fe5",
			999 => x"006a0fe5",
			1000 => x"04f80fe5",
			1001 => x"06018d04",
			1002 => x"065c0fe5",
			1003 => x"fe630fe5",
			1004 => x"05086a08",
			1005 => x"0706a104",
			1006 => x"fe440fe5",
			1007 => x"04020fe5",
			1008 => x"08035e0c",
			1009 => x"08034508",
			1010 => x"09021204",
			1011 => x"055f0fe5",
			1012 => x"063b0fe5",
			1013 => x"04720fe5",
			1014 => x"07072604",
			1015 => x"fe600fe5",
			1016 => x"01180fe5",
			1017 => x"020a5b08",
			1018 => x"0c063a04",
			1019 => x"ff5e1079",
			1020 => x"00001079",
			1021 => x"0508dc24",
			1022 => x"01015018",
			1023 => x"040d1b10",
			1024 => x"0f0b880c",
			1025 => x"00039504",
			1026 => x"00001079",
			1027 => x"0f0a7c04",
			1028 => x"00001079",
			1029 => x"ffc01079",
			1030 => x"00001079",
			1031 => x"00048104",
			1032 => x"006a1079",
			1033 => x"00001079",
			1034 => x"0e0b6308",
			1035 => x"0c063004",
			1036 => x"00001079",
			1037 => x"00ca1079",
			1038 => x"00001079",
			1039 => x"0c06a414",
			1040 => x"09022a04",
			1041 => x"00001079",
			1042 => x"030b1b04",
			1043 => x"00001079",
			1044 => x"07072508",
			1045 => x"0d094e04",
			1046 => x"00001079",
			1047 => x"ff3c1079",
			1048 => x"00001079",
			1049 => x"0601ca08",
			1050 => x"0e0ac904",
			1051 => x"00001079",
			1052 => x"00b61079",
			1053 => x"00001079",
			1054 => x"0901ce04",
			1055 => x"fef610ed",
			1056 => x"040b6320",
			1057 => x"0706df14",
			1058 => x"01015910",
			1059 => x"06018804",
			1060 => x"000010ed",
			1061 => x"0b079308",
			1062 => x"0a025604",
			1063 => x"000010ed",
			1064 => x"feee10ed",
			1065 => x"000010ed",
			1066 => x"000010ed",
			1067 => x"0d096908",
			1068 => x"00039e04",
			1069 => x"00a710ed",
			1070 => x"000010ed",
			1071 => x"000010ed",
			1072 => x"0601c214",
			1073 => x"0c06dc10",
			1074 => x"0c063004",
			1075 => x"000010ed",
			1076 => x"0e0b5108",
			1077 => x"07066e04",
			1078 => x"000010ed",
			1079 => x"00c510ed",
			1080 => x"000010ed",
			1081 => x"000010ed",
			1082 => x"ffd610ed",
			1083 => x"020a5b0c",
			1084 => x"0802d804",
			1085 => x"00001171",
			1086 => x"0c065004",
			1087 => x"ff651171",
			1088 => x"00001171",
			1089 => x"0601ca34",
			1090 => x"0003a318",
			1091 => x"0802e308",
			1092 => x"09020504",
			1093 => x"00001171",
			1094 => x"00461171",
			1095 => x"09022a04",
			1096 => x"00001171",
			1097 => x"030b1304",
			1098 => x"00001171",
			1099 => x"09023904",
			1100 => x"ff471171",
			1101 => x"00001171",
			1102 => x"09021b14",
			1103 => x"040d1b0c",
			1104 => x"0f0b8808",
			1105 => x"0f0a8a04",
			1106 => x"00001171",
			1107 => x"ffda1171",
			1108 => x"00001171",
			1109 => x"040df504",
			1110 => x"00331171",
			1111 => x"00001171",
			1112 => x"0c066c04",
			1113 => x"00001171",
			1114 => x"00c81171",
			1115 => x"ffd61171",
			1116 => x"0901dd08",
			1117 => x"040da904",
			1118 => x"fe961215",
			1119 => x"00001215",
			1120 => x"0e0b0734",
			1121 => x"040b4a20",
			1122 => x"06019110",
			1123 => x"05086a08",
			1124 => x"06017d04",
			1125 => x"00001215",
			1126 => x"ff3c1215",
			1127 => x"040b4604",
			1128 => x"01191215",
			1129 => x"00001215",
			1130 => x"07070b0c",
			1131 => x"040b3c08",
			1132 => x"0c068d04",
			1133 => x"ff1a1215",
			1134 => x"00001215",
			1135 => x"00001215",
			1136 => x"00001215",
			1137 => x"0601a90c",
			1138 => x"0b071004",
			1139 => x"00001215",
			1140 => x"0c06c404",
			1141 => x"01181215",
			1142 => x"00001215",
			1143 => x"0c06a104",
			1144 => x"00001215",
			1145 => x"ffcb1215",
			1146 => x"09023f0c",
			1147 => x"07070d08",
			1148 => x"0c06a404",
			1149 => x"fee71215",
			1150 => x"00001215",
			1151 => x"00001215",
			1152 => x"0601cc08",
			1153 => x"0c068a04",
			1154 => x"00001215",
			1155 => x"00e51215",
			1156 => x"ff9d1215",
			1157 => x"0902051c",
			1158 => x"020a2d04",
			1159 => x"fe6312c9",
			1160 => x"0e0a7014",
			1161 => x"0c05f604",
			1162 => x"fe8612c9",
			1163 => x"07062c04",
			1164 => x"03d612c9",
			1165 => x"0901a904",
			1166 => x"fe7e12c9",
			1167 => x"0601a704",
			1168 => x"013a12c9",
			1169 => x"ff4e12c9",
			1170 => x"fe6a12c9",
			1171 => x"05086a14",
			1172 => x"040b8e08",
			1173 => x"0802d704",
			1174 => x"000a12c9",
			1175 => x"fe3412c9",
			1176 => x"040b9d04",
			1177 => x"099c12c9",
			1178 => x"0f0b3b04",
			1179 => x"019b12c9",
			1180 => x"fee712c9",
			1181 => x"0601b71c",
			1182 => x"09021208",
			1183 => x"0a027504",
			1184 => x"019212c9",
			1185 => x"ff6312c9",
			1186 => x"0d09750c",
			1187 => x"0d095004",
			1188 => x"01a712c9",
			1189 => x"0706e304",
			1190 => x"ff1012c9",
			1191 => x"016d12c9",
			1192 => x"0003a704",
			1193 => x"feed12c9",
			1194 => x"018c12c9",
			1195 => x"040c4704",
			1196 => x"fec612c9",
			1197 => x"08036e08",
			1198 => x"0c068b04",
			1199 => x"ffd012c9",
			1200 => x"01ec12c9",
			1201 => x"fec212c9",
			1202 => x"0c061304",
			1203 => x"ff5d134d",
			1204 => x"0601b62c",
			1205 => x"040b631c",
			1206 => x"0b078210",
			1207 => x"06018904",
			1208 => x"0000134d",
			1209 => x"01015908",
			1210 => x"0706e204",
			1211 => x"ff3d134d",
			1212 => x"0000134d",
			1213 => x"0000134d",
			1214 => x"0b07b508",
			1215 => x"01014704",
			1216 => x"0000134d",
			1217 => x"006e134d",
			1218 => x"0000134d",
			1219 => x"0901ce04",
			1220 => x"0000134d",
			1221 => x"020bbc08",
			1222 => x"07066e04",
			1223 => x"0000134d",
			1224 => x"00b6134d",
			1225 => x"0000134d",
			1226 => x"0e0c8c10",
			1227 => x"0101850c",
			1228 => x"020b5304",
			1229 => x"0000134d",
			1230 => x"0a02ae04",
			1231 => x"0000134d",
			1232 => x"ff48134d",
			1233 => x"0000134d",
			1234 => x"0000134d",
			1235 => x"01012308",
			1236 => x"040da904",
			1237 => x"fe9013f9",
			1238 => x"000013f9",
			1239 => x"0003a324",
			1240 => x"0f0b0314",
			1241 => x"0706c910",
			1242 => x"0802d804",
			1243 => x"000013f9",
			1244 => x"040b1608",
			1245 => x"0b077104",
			1246 => x"feef13f9",
			1247 => x"000013f9",
			1248 => x"000013f9",
			1249 => x"010713f9",
			1250 => x"01015808",
			1251 => x"0508cf04",
			1252 => x"000013f9",
			1253 => x"002013f9",
			1254 => x"0d094e04",
			1255 => x"000013f9",
			1256 => x"feb813f9",
			1257 => x"0601a110",
			1258 => x"0b071004",
			1259 => x"000013f9",
			1260 => x"040b5b04",
			1261 => x"000013f9",
			1262 => x"05091b04",
			1263 => x"013313f9",
			1264 => x"000013f9",
			1265 => x"040c470c",
			1266 => x"0a028d04",
			1267 => x"000013f9",
			1268 => x"01017904",
			1269 => x"fefb13f9",
			1270 => x"000013f9",
			1271 => x"00042908",
			1272 => x"08033304",
			1273 => x"000013f9",
			1274 => x"00c013f9",
			1275 => x"040d4204",
			1276 => x"ff2d13f9",
			1277 => x"001213f9",
			1278 => x"0c061304",
			1279 => x"ff49147d",
			1280 => x"0e0aa218",
			1281 => x"020a8304",
			1282 => x"0000147d",
			1283 => x"08036b10",
			1284 => x"01010b04",
			1285 => x"0000147d",
			1286 => x"0c06a108",
			1287 => x"0a025104",
			1288 => x"0000147d",
			1289 => x"00c1147d",
			1290 => x"0000147d",
			1291 => x"0000147d",
			1292 => x"0c068d14",
			1293 => x"0802e304",
			1294 => x"0000147d",
			1295 => x"09023b0c",
			1296 => x"07072408",
			1297 => x"01014304",
			1298 => x"0000147d",
			1299 => x"ff57147d",
			1300 => x"0000147d",
			1301 => x"0000147d",
			1302 => x"0803420c",
			1303 => x"07072808",
			1304 => x"01014904",
			1305 => x"0000147d",
			1306 => x"0099147d",
			1307 => x"0000147d",
			1308 => x"01017904",
			1309 => x"ffb5147d",
			1310 => x"0000147d",
			1311 => x"01013f20",
			1312 => x"06018a04",
			1313 => x"fe651551",
			1314 => x"0f0aa610",
			1315 => x"040d2e08",
			1316 => x"0f0a9204",
			1317 => x"fec91551",
			1318 => x"00001551",
			1319 => x"0100d804",
			1320 => x"ff8a1551",
			1321 => x"02191551",
			1322 => x"06019408",
			1323 => x"020afb04",
			1324 => x"ff6a1551",
			1325 => x"00991551",
			1326 => x"fe8e1551",
			1327 => x"01015028",
			1328 => x"06018c14",
			1329 => x"030a3904",
			1330 => x"feca1551",
			1331 => x"040b5d0c",
			1332 => x"040b1504",
			1333 => x"017c1551",
			1334 => x"040b2204",
			1335 => x"ffd51551",
			1336 => x"00a51551",
			1337 => x"036a1551",
			1338 => x"040c2c10",
			1339 => x"0e0a5108",
			1340 => x"0b070104",
			1341 => x"ffdc1551",
			1342 => x"00de1551",
			1343 => x"040b0204",
			1344 => x"00001551",
			1345 => x"fdb41551",
			1346 => x"00fd1551",
			1347 => x"08034d1c",
			1348 => x"0d097514",
			1349 => x"0706a10c",
			1350 => x"0e0a9a08",
			1351 => x"020ab704",
			1352 => x"00001551",
			1353 => x"01301551",
			1354 => x"fed21551",
			1355 => x"07073804",
			1356 => x"01941551",
			1357 => x"00001551",
			1358 => x"0e0b0e04",
			1359 => x"fe641551",
			1360 => x"01931551",
			1361 => x"07072504",
			1362 => x"feb11551",
			1363 => x"00001551",
			1364 => x"0901fc24",
			1365 => x"06018a04",
			1366 => x"fe68162d",
			1367 => x"0f0a7c0c",
			1368 => x"09016b04",
			1369 => x"ff67162d",
			1370 => x"040be904",
			1371 => x"0000162d",
			1372 => x"01c8162d",
			1373 => x"01012304",
			1374 => x"fe82162d",
			1375 => x"01012a08",
			1376 => x"0601a604",
			1377 => x"010d162d",
			1378 => x"0000162d",
			1379 => x"06019d04",
			1380 => x"0000162d",
			1381 => x"feec162d",
			1382 => x"01014e28",
			1383 => x"01014514",
			1384 => x"040b8e08",
			1385 => x"06018304",
			1386 => x"0000162d",
			1387 => x"ff2c162d",
			1388 => x"0508a308",
			1389 => x"0b071004",
			1390 => x"0000162d",
			1391 => x"01d1162d",
			1392 => x"ffa2162d",
			1393 => x"0802dd08",
			1394 => x"030a3904",
			1395 => x"0000162d",
			1396 => x"00d8162d",
			1397 => x"00040808",
			1398 => x"09021904",
			1399 => x"fe8a162d",
			1400 => x"0000162d",
			1401 => x"0000162d",
			1402 => x"05086a08",
			1403 => x"0e0a2a04",
			1404 => x"001b162d",
			1405 => x"fe90162d",
			1406 => x"0d094e08",
			1407 => x"0e0b6304",
			1408 => x"0191162d",
			1409 => x"0000162d",
			1410 => x"0706df04",
			1411 => x"fdfa162d",
			1412 => x"00039a08",
			1413 => x"09022e04",
			1414 => x"011d162d",
			1415 => x"ff0f162d",
			1416 => x"08036804",
			1417 => x"0149162d",
			1418 => x"ff0e162d",
			1419 => x"0101280c",
			1420 => x"0100f804",
			1421 => x"fe6916e1",
			1422 => x"040d2e04",
			1423 => x"fea316e1",
			1424 => x"007816e1",
			1425 => x"01015c3c",
			1426 => x"0f0b031c",
			1427 => x"0d087f08",
			1428 => x"08033a04",
			1429 => x"fec616e1",
			1430 => x"000016e1",
			1431 => x"0c06c410",
			1432 => x"0f0a6e08",
			1433 => x"0c063a04",
			1434 => x"fea316e1",
			1435 => x"00f316e1",
			1436 => x"0f0af304",
			1437 => x"017116e1",
			1438 => x"007816e1",
			1439 => x"ff5416e1",
			1440 => x"0706f514",
			1441 => x"040c6610",
			1442 => x"0f0b0908",
			1443 => x"020af104",
			1444 => x"f99d16e1",
			1445 => x"000016e1",
			1446 => x"0b07a104",
			1447 => x"fddf16e1",
			1448 => x"000016e1",
			1449 => x"006616e1",
			1450 => x"0601b008",
			1451 => x"01014704",
			1452 => x"000016e1",
			1453 => x"016716e1",
			1454 => x"fee116e1",
			1455 => x"0a026408",
			1456 => x"030b1304",
			1457 => x"014816e1",
			1458 => x"feb416e1",
			1459 => x"0601c208",
			1460 => x"0b075f04",
			1461 => x"000016e1",
			1462 => x"019616e1",
			1463 => x"002e16e1",
			1464 => x"09018b04",
			1465 => x"ff09176d",
			1466 => x"040c8530",
			1467 => x"06018c0c",
			1468 => x"09020504",
			1469 => x"0000176d",
			1470 => x"0b071004",
			1471 => x"0000176d",
			1472 => x"0091176d",
			1473 => x"01015008",
			1474 => x"0f0a8a04",
			1475 => x"0000176d",
			1476 => x"ff2b176d",
			1477 => x"0b07b510",
			1478 => x"0802e008",
			1479 => x"0706df04",
			1480 => x"ff9f176d",
			1481 => x"0000176d",
			1482 => x"020b6904",
			1483 => x"00c0176d",
			1484 => x"0000176d",
			1485 => x"09022e04",
			1486 => x"0000176d",
			1487 => x"0f0afc04",
			1488 => x"0000176d",
			1489 => x"ff6f176d",
			1490 => x"0a02db10",
			1491 => x"0d08f404",
			1492 => x"0103176d",
			1493 => x"0d097704",
			1494 => x"0000176d",
			1495 => x"09022e04",
			1496 => x"0000176d",
			1497 => x"0062176d",
			1498 => x"0000176d",
			1499 => x"0c05d804",
			1500 => x"fe8d17f1",
			1501 => x"040d4238",
			1502 => x"0601a528",
			1503 => x"040b6318",
			1504 => x"0802e30c",
			1505 => x"0b073304",
			1506 => x"000017f1",
			1507 => x"040b4604",
			1508 => x"011617f1",
			1509 => x"000017f1",
			1510 => x"01016008",
			1511 => x"0c068d04",
			1512 => x"ff1117f1",
			1513 => x"000017f1",
			1514 => x"004a17f1",
			1515 => x"0c061404",
			1516 => x"ffbc17f1",
			1517 => x"0f0b9808",
			1518 => x"01010b04",
			1519 => x"000017f1",
			1520 => x"014017f1",
			1521 => x"000017f1",
			1522 => x"01015f08",
			1523 => x"040cce04",
			1524 => x"fee717f1",
			1525 => x"000017f1",
			1526 => x"08035604",
			1527 => x"009717f1",
			1528 => x"ffa917f1",
			1529 => x"0a02dd04",
			1530 => x"01a117f1",
			1531 => x"fff417f1",
			1532 => x"01014740",
			1533 => x"01013f30",
			1534 => x"0100f804",
			1535 => x"fe5418a5",
			1536 => x"0c063314",
			1537 => x"0100fa08",
			1538 => x"07064604",
			1539 => x"01a418a5",
			1540 => x"fe8e18a5",
			1541 => x"0c061404",
			1542 => x"fe5718a5",
			1543 => x"01011904",
			1544 => x"000018a5",
			1545 => x"fe5b18a5",
			1546 => x"07069b0c",
			1547 => x"06019104",
			1548 => x"fe8d18a5",
			1549 => x"030a9904",
			1550 => x"034518a5",
			1551 => x"fed018a5",
			1552 => x"0c065208",
			1553 => x"01012304",
			1554 => x"fe8218a5",
			1555 => x"01a518a5",
			1556 => x"fe5418a5",
			1557 => x"0706a108",
			1558 => x"0c063204",
			1559 => x"fe5a18a5",
			1560 => x"000018a5",
			1561 => x"030ac504",
			1562 => x"039a18a5",
			1563 => x"00cf18a5",
			1564 => x"0d08b304",
			1565 => x"fe4c18a5",
			1566 => x"0601cc14",
			1567 => x"040d0e10",
			1568 => x"08034d0c",
			1569 => x"05086a04",
			1570 => x"010118a5",
			1571 => x"01015004",
			1572 => x"023318a5",
			1573 => x"026618a5",
			1574 => x"ff0218a5",
			1575 => x"045c18a5",
			1576 => x"fe6b18a5",
			1577 => x"020a2d08",
			1578 => x"030a3904",
			1579 => x"fe6d1949",
			1580 => x"00001949",
			1581 => x"0f0adf18",
			1582 => x"0c05d804",
			1583 => x"ff7d1949",
			1584 => x"0c06c310",
			1585 => x"09016b04",
			1586 => x"00001949",
			1587 => x"040a9504",
			1588 => x"00001949",
			1589 => x"06017d04",
			1590 => x"00001949",
			1591 => x"01471949",
			1592 => x"ffce1949",
			1593 => x"01016128",
			1594 => x"0b07b51c",
			1595 => x"0706e210",
			1596 => x"0508a308",
			1597 => x"0601b204",
			1598 => x"00381949",
			1599 => x"ff231949",
			1600 => x"01015c04",
			1601 => x"fe701949",
			1602 => x"00001949",
			1603 => x"01014e08",
			1604 => x"0c068a04",
			1605 => x"00001949",
			1606 => x"ff671949",
			1607 => x"014f1949",
			1608 => x"09022e08",
			1609 => x"040bbd04",
			1610 => x"00d01949",
			1611 => x"fef71949",
			1612 => x"fdca1949",
			1613 => x"0a02cb08",
			1614 => x"0706b704",
			1615 => x"00001949",
			1616 => x"01711949",
			1617 => x"00001949",
			1618 => x"020a1004",
			1619 => x"fe8619d5",
			1620 => x"040d4238",
			1621 => x"0601a52c",
			1622 => x"040b631c",
			1623 => x"0003950c",
			1624 => x"0706a104",
			1625 => x"000019d5",
			1626 => x"01014704",
			1627 => x"000019d5",
			1628 => x"012019d5",
			1629 => x"0706f508",
			1630 => x"01015c04",
			1631 => x"fed219d5",
			1632 => x"000019d5",
			1633 => x"07072204",
			1634 => x"00b519d5",
			1635 => x"000019d5",
			1636 => x"0c061404",
			1637 => x"ff9b19d5",
			1638 => x"0e0b5108",
			1639 => x"01010b04",
			1640 => x"000019d5",
			1641 => x"014e19d5",
			1642 => x"000019d5",
			1643 => x"01015f04",
			1644 => x"fee519d5",
			1645 => x"08035604",
			1646 => x"00ac19d5",
			1647 => x"ff8e19d5",
			1648 => x"0a02dd08",
			1649 => x"06019104",
			1650 => x"000019d5",
			1651 => x"01c319d5",
			1652 => x"ffcb19d5",
			1653 => x"0901fa10",
			1654 => x"0901b204",
			1655 => x"fe671aa1",
			1656 => x"040cc604",
			1657 => x"fe961aa1",
			1658 => x"0601b604",
			1659 => x"01811aa1",
			1660 => x"ffee1aa1",
			1661 => x"0706c924",
			1662 => x"0f0bae20",
			1663 => x"040b8010",
			1664 => x"0b07710c",
			1665 => x"09022908",
			1666 => x"06017d04",
			1667 => x"00001aa1",
			1668 => x"fe6a1aa1",
			1669 => x"00441aa1",
			1670 => x"010d1aa1",
			1671 => x"0601b20c",
			1672 => x"0b071004",
			1673 => x"00001aa1",
			1674 => x"030b4b04",
			1675 => x"01c21aa1",
			1676 => x"00001aa1",
			1677 => x"ffc41aa1",
			1678 => x"fe1e1aa1",
			1679 => x"0508dc0c",
			1680 => x"09021208",
			1681 => x"09020e04",
			1682 => x"004a1aa1",
			1683 => x"ffff1aa1",
			1684 => x"01991aa1",
			1685 => x"0706f510",
			1686 => x"0508de08",
			1687 => x"0a026904",
			1688 => x"f9431aa1",
			1689 => x"00001aa1",
			1690 => x"0508f804",
			1691 => x"00df1aa1",
			1692 => x"00001aa1",
			1693 => x"0a02a910",
			1694 => x"00039a08",
			1695 => x"030b2304",
			1696 => x"00db1aa1",
			1697 => x"fe5d1aa1",
			1698 => x"09021804",
			1699 => x"00001aa1",
			1700 => x"018a1aa1",
			1701 => x"09025b04",
			1702 => x"fe631aa1",
			1703 => x"005b1aa1",
			1704 => x"09018b04",
			1705 => x"fee31b3d",
			1706 => x"0d08da14",
			1707 => x"040d2e10",
			1708 => x"0901dd04",
			1709 => x"ffd01b3d",
			1710 => x"0c063004",
			1711 => x"00001b3d",
			1712 => x"0c064d04",
			1713 => x"006b1b3d",
			1714 => x"00001b3d",
			1715 => x"00d71b3d",
			1716 => x"0b078210",
			1717 => x"0101590c",
			1718 => x"06018904",
			1719 => x"00001b3d",
			1720 => x"0c068704",
			1721 => x"fec01b3d",
			1722 => x"00001b3d",
			1723 => x"00001b3d",
			1724 => x"0d094110",
			1725 => x"020bbc0c",
			1726 => x"01013b04",
			1727 => x"00001b3d",
			1728 => x"0c06c204",
			1729 => x"00971b3d",
			1730 => x"00001b3d",
			1731 => x"00001b3d",
			1732 => x"08034710",
			1733 => x"020ae608",
			1734 => x"020ad604",
			1735 => x"00001b3d",
			1736 => x"ff8f1b3d",
			1737 => x"00039a04",
			1738 => x"00001b3d",
			1739 => x"00a61b3d",
			1740 => x"01018304",
			1741 => x"ff811b3d",
			1742 => x"00001b3d",
			1743 => x"0c061304",
			1744 => x"fe7d1bf1",
			1745 => x"0b07b538",
			1746 => x"09021f24",
			1747 => x"0e0a9214",
			1748 => x"0901a904",
			1749 => x"ff861bf1",
			1750 => x"040b7608",
			1751 => x"0706a104",
			1752 => x"ff341bf1",
			1753 => x"009d1bf1",
			1754 => x"0601a904",
			1755 => x"01521bf1",
			1756 => x"00001bf1",
			1757 => x"06018d04",
			1758 => x"00001bf1",
			1759 => x"0508df08",
			1760 => x"040c6604",
			1761 => x"fe931bf1",
			1762 => x"00001bf1",
			1763 => x"00001bf1",
			1764 => x"0c06520c",
			1765 => x"0c063404",
			1766 => x"001e1bf1",
			1767 => x"0706c904",
			1768 => x"ff431bf1",
			1769 => x"00001bf1",
			1770 => x"09026404",
			1771 => x"015a1bf1",
			1772 => x"00001bf1",
			1773 => x"09023918",
			1774 => x"0802e808",
			1775 => x"09022e04",
			1776 => x"00291bf1",
			1777 => x"00001bf1",
			1778 => x"0c068c04",
			1779 => x"00001bf1",
			1780 => x"06018e04",
			1781 => x"00001bf1",
			1782 => x"0d094104",
			1783 => x"00001bf1",
			1784 => x"fead1bf1",
			1785 => x"08036804",
			1786 => x"00b71bf1",
			1787 => x"00001bf1",
			1788 => x"020a5b08",
			1789 => x"0c063a04",
			1790 => x"fe6d1cbd",
			1791 => x"00001cbd",
			1792 => x"01015c48",
			1793 => x"0f0adf1c",
			1794 => x"0902020c",
			1795 => x"040cb604",
			1796 => x"ff521cbd",
			1797 => x"08037f04",
			1798 => x"00d51cbd",
			1799 => x"00001cbd",
			1800 => x"0f0a8a08",
			1801 => x"0c065204",
			1802 => x"ff801cbd",
			1803 => x"005b1cbd",
			1804 => x"0c063204",
			1805 => x"00001cbd",
			1806 => x"017b1cbd",
			1807 => x"020ae610",
			1808 => x"0508dd0c",
			1809 => x"00039504",
			1810 => x"00001cbd",
			1811 => x"0f0aed04",
			1812 => x"00001cbd",
			1813 => x"fe381cbd",
			1814 => x"000c1cbd",
			1815 => x"0a028d10",
			1816 => x"09022a08",
			1817 => x"0901fa04",
			1818 => x"00001cbd",
			1819 => x"012e1cbd",
			1820 => x"0a026d04",
			1821 => x"ff6e1cbd",
			1822 => x"00001cbd",
			1823 => x"0d091b08",
			1824 => x"01014104",
			1825 => x"ff111cbd",
			1826 => x"00881cbd",
			1827 => x"fed71cbd",
			1828 => x"0d09750c",
			1829 => x"05086a04",
			1830 => x"00001cbd",
			1831 => x"0f0c0904",
			1832 => x"01711cbd",
			1833 => x"00001cbd",
			1834 => x"09025204",
			1835 => x"ff2f1cbd",
			1836 => x"08037704",
			1837 => x"012a1cbd",
			1838 => x"ff9d1cbd",
			1839 => x"020a2d08",
			1840 => x"0b074404",
			1841 => x"fe671d89",
			1842 => x"00001d89",
			1843 => x"01014e34",
			1844 => x"0601a728",
			1845 => x"040b8e14",
			1846 => x"0b07710c",
			1847 => x"06018308",
			1848 => x"06017c04",
			1849 => x"00001d89",
			1850 => x"00131d89",
			1851 => x"fe621d89",
			1852 => x"01014504",
			1853 => x"00001d89",
			1854 => x"01061d89",
			1855 => x"09016b04",
			1856 => x"ff3e1d89",
			1857 => x"06019908",
			1858 => x"06018904",
			1859 => x"00001d89",
			1860 => x"01fd1d89",
			1861 => x"01012304",
			1862 => x"ff531d89",
			1863 => x"01091d89",
			1864 => x"0706a108",
			1865 => x"07068604",
			1866 => x"ff401d89",
			1867 => x"00001d89",
			1868 => x"fe6e1d89",
			1869 => x"05086a0c",
			1870 => x"01015208",
			1871 => x"040ba404",
			1872 => x"00001d89",
			1873 => x"006d1d89",
			1874 => x"fe561d89",
			1875 => x"0d094e0c",
			1876 => x"020b7704",
			1877 => x"01971d89",
			1878 => x"0706ce04",
			1879 => x"ffcc1d89",
			1880 => x"00871d89",
			1881 => x"0706df04",
			1882 => x"fdbd1d89",
			1883 => x"01016008",
			1884 => x"01015f04",
			1885 => x"00e01d89",
			1886 => x"fe741d89",
			1887 => x"08036804",
			1888 => x"018b1d89",
			1889 => x"ff2c1d89",
			1890 => x"0100e504",
			1891 => x"fe6f1e25",
			1892 => x"01016144",
			1893 => x"030b1324",
			1894 => x"0101501c",
			1895 => x"040c0410",
			1896 => x"0c066d08",
			1897 => x"0706e104",
			1898 => x"fe8e1e25",
			1899 => x"00001e25",
			1900 => x"0a027204",
			1901 => x"007c1e25",
			1902 => x"ffbf1e25",
			1903 => x"0601b708",
			1904 => x"030a8104",
			1905 => x"01391e25",
			1906 => x"00001e25",
			1907 => x"ff751e25",
			1908 => x"05084d04",
			1909 => x"00001e25",
			1910 => x"017a1e25",
			1911 => x"0706f50c",
			1912 => x"01015304",
			1913 => x"00001e25",
			1914 => x"01015c04",
			1915 => x"fdef1e25",
			1916 => x"00001e25",
			1917 => x"0a027008",
			1918 => x"01015f04",
			1919 => x"011b1e25",
			1920 => x"ffb61e25",
			1921 => x"0b07a504",
			1922 => x"00001e25",
			1923 => x"0c06a104",
			1924 => x"00001e25",
			1925 => x"fede1e25",
			1926 => x"08036504",
			1927 => x"01701e25",
			1928 => x"00001e25",
			1929 => x"020a2d08",
			1930 => x"0b074404",
			1931 => x"fe6a1ef3",
			1932 => x"00001ef3",
			1933 => x"0101594c",
			1934 => x"0e0aa22c",
			1935 => x"05086a18",
			1936 => x"0003e20c",
			1937 => x"0f0af508",
			1938 => x"0802d404",
			1939 => x"00001ef3",
			1940 => x"fe681ef3",
			1941 => x"00001ef3",
			1942 => x"0c05f604",
			1943 => x"ff5e1ef3",
			1944 => x"09016b04",
			1945 => x"00001ef3",
			1946 => x"012f1ef3",
			1947 => x"09020e10",
			1948 => x"0b077308",
			1949 => x"0c066c04",
			1950 => x"00001ef3",
			1951 => x"00aa1ef3",
			1952 => x"020aa104",
			1953 => x"00001ef3",
			1954 => x"fefc1ef3",
			1955 => x"016b1ef3",
			1956 => x"0706e214",
			1957 => x"040c6610",
			1958 => x"0b079308",
			1959 => x"0f0aed04",
			1960 => x"00001ef3",
			1961 => x"fdf01ef3",
			1962 => x"0003b304",
			1963 => x"002a1ef3",
			1964 => x"00001ef3",
			1965 => x"00001ef3",
			1966 => x"08030204",
			1967 => x"01501ef3",
			1968 => x"0b078404",
			1969 => x"00001ef3",
			1970 => x"fec21ef3",
			1971 => x"0e0adc04",
			1972 => x"01861ef3",
			1973 => x"00039e04",
			1974 => x"fe8c1ef3",
			1975 => x"08036e08",
			1976 => x"0c065204",
			1977 => x"ffda1ef3",
			1978 => x"01921ef3",
			1979 => x"ff291ef3",
			1980 => x"00001ef5",
			1981 => x"0b083804",
			1982 => x"00001f01",
			1983 => x"fcf81f01",
			1984 => x"05095e04",
			1985 => x"00001f0d",
			1986 => x"fee31f0d",
			1987 => x"040bf104",
			1988 => x"00001f21",
			1989 => x"040e2304",
			1990 => x"00291f21",
			1991 => x"00001f21",
			1992 => x"0c06a108",
			1993 => x"0c05d804",
			1994 => x"00001f35",
			1995 => x"00271f35",
			1996 => x"fffa1f35",
			1997 => x"0509d604",
			1998 => x"00001f49",
			1999 => x"0d0a5304",
			2000 => x"f22d1f49",
			2001 => x"00001f49",
			2002 => x"040d2e08",
			2003 => x"08034704",
			2004 => x"00001f5d",
			2005 => x"ff671f5d",
			2006 => x"00001f5d",
			2007 => x"0d0a110c",
			2008 => x"040c3e04",
			2009 => x"fffc1f79",
			2010 => x"040e2304",
			2011 => x"001a1f79",
			2012 => x"00001f79",
			2013 => x"ff8c1f79",
			2014 => x"040bf108",
			2015 => x"040b1404",
			2016 => x"00001f9d",
			2017 => x"fff71f9d",
			2018 => x"040e2308",
			2019 => x"040c8504",
			2020 => x"00001f9d",
			2021 => x"002e1f9d",
			2022 => x"00001f9d",
			2023 => x"0a02880c",
			2024 => x"0a026204",
			2025 => x"00001fc1",
			2026 => x"06017d04",
			2027 => x"00001fc1",
			2028 => x"004a1fc1",
			2029 => x"06019904",
			2030 => x"00001fc1",
			2031 => x"ffe61fc1",
			2032 => x"0101500c",
			2033 => x"0a02d108",
			2034 => x"0a026504",
			2035 => x"00001fe5",
			2036 => x"ffe11fe5",
			2037 => x"00001fe5",
			2038 => x"0a02a904",
			2039 => x"002d1fe5",
			2040 => x"00001fe5",
			2041 => x"0c06dc0c",
			2042 => x"040c5e04",
			2043 => x"00002009",
			2044 => x"040e2304",
			2045 => x"001c2009",
			2046 => x"00002009",
			2047 => x"07072804",
			2048 => x"00002009",
			2049 => x"ff692009",
			2050 => x"0a02880c",
			2051 => x"0a026204",
			2052 => x"00002035",
			2053 => x"06017d04",
			2054 => x"00002035",
			2055 => x"00532035",
			2056 => x"06019904",
			2057 => x"00002035",
			2058 => x"0003cc04",
			2059 => x"00002035",
			2060 => x"ffde2035",
			2061 => x"08033f0c",
			2062 => x"0003a304",
			2063 => x"00002061",
			2064 => x"00041404",
			2065 => x"000a2061",
			2066 => x"00002061",
			2067 => x"01017908",
			2068 => x"0004a704",
			2069 => x"ffa52061",
			2070 => x"00002061",
			2071 => x"00002061",
			2072 => x"040d2e10",
			2073 => x"0803470c",
			2074 => x"040bfa08",
			2075 => x"040ac204",
			2076 => x"00002085",
			2077 => x"fffc2085",
			2078 => x"00002085",
			2079 => x"ff5a2085",
			2080 => x"00002085",
			2081 => x"07076410",
			2082 => x"0706c904",
			2083 => x"000020a9",
			2084 => x"0b077104",
			2085 => x"000020a9",
			2086 => x"0d08f404",
			2087 => x"000020a9",
			2088 => x"002720a9",
			2089 => x"fffc20a9",
			2090 => x"020ad604",
			2091 => x"000020cd",
			2092 => x"0101810c",
			2093 => x"040d0e08",
			2094 => x"08032504",
			2095 => x"000020cd",
			2096 => x"ff9120cd",
			2097 => x"000020cd",
			2098 => x"000020cd",
			2099 => x"09020a10",
			2100 => x"07066f08",
			2101 => x"0c05d804",
			2102 => x"00002101",
			2103 => x"00052101",
			2104 => x"05080104",
			2105 => x"00002101",
			2106 => x"ffbf2101",
			2107 => x"0c065204",
			2108 => x"00002101",
			2109 => x"07072804",
			2110 => x"00602101",
			2111 => x"00002101",
			2112 => x"040c5e10",
			2113 => x"040b3604",
			2114 => x"00002135",
			2115 => x"020af408",
			2116 => x"09023204",
			2117 => x"ffd32135",
			2118 => x"00002135",
			2119 => x"00002135",
			2120 => x"0901bc04",
			2121 => x"00002135",
			2122 => x"0601cc04",
			2123 => x"00522135",
			2124 => x"00002135",
			2125 => x"0c06dc14",
			2126 => x"01014e08",
			2127 => x"0f0a6e04",
			2128 => x"00002169",
			2129 => x"fff72169",
			2130 => x"0706df04",
			2131 => x"00002169",
			2132 => x"01018904",
			2133 => x"00352169",
			2134 => x"00002169",
			2135 => x"0b082804",
			2136 => x"00002169",
			2137 => x"fd9d2169",
			2138 => x"0c06dc14",
			2139 => x"09021f04",
			2140 => x"0000219d",
			2141 => x"06018d04",
			2142 => x"0000219d",
			2143 => x"09027408",
			2144 => x"05084d04",
			2145 => x"0000219d",
			2146 => x"003e219d",
			2147 => x"0000219d",
			2148 => x"0b082804",
			2149 => x"0000219d",
			2150 => x"fdfb219d",
			2151 => x"08035e14",
			2152 => x"0c063004",
			2153 => x"000021d1",
			2154 => x"00038504",
			2155 => x"000021d1",
			2156 => x"0d086604",
			2157 => x"000021d1",
			2158 => x"0c06dc04",
			2159 => x"001b21d1",
			2160 => x"000021d1",
			2161 => x"0004a704",
			2162 => x"ffac21d1",
			2163 => x"000021d1",
			2164 => x"0509ab14",
			2165 => x"0b077104",
			2166 => x"000021fd",
			2167 => x"05088604",
			2168 => x"000021fd",
			2169 => x"0c065004",
			2170 => x"000021fd",
			2171 => x"0c06de04",
			2172 => x"002f21fd",
			2173 => x"000021fd",
			2174 => x"fffb21fd",
			2175 => x"07072814",
			2176 => x"0901bc04",
			2177 => x"00002239",
			2178 => x"020a9904",
			2179 => x"00002239",
			2180 => x"08036b08",
			2181 => x"07065a04",
			2182 => x"00002239",
			2183 => x"004c2239",
			2184 => x"00002239",
			2185 => x"06019204",
			2186 => x"00002239",
			2187 => x"0b07c304",
			2188 => x"00002239",
			2189 => x"ff1c2239",
			2190 => x"040da918",
			2191 => x"01016010",
			2192 => x"00039504",
			2193 => x"0000227d",
			2194 => x"040d0e08",
			2195 => x"0a026104",
			2196 => x"0000227d",
			2197 => x"ffbc227d",
			2198 => x"0000227d",
			2199 => x"0601c204",
			2200 => x"0048227d",
			2201 => x"0000227d",
			2202 => x"0a02dd08",
			2203 => x"0100e504",
			2204 => x"0000227d",
			2205 => x"015d227d",
			2206 => x"0000227d",
			2207 => x"040c4714",
			2208 => x"0706df10",
			2209 => x"0c06870c",
			2210 => x"01016808",
			2211 => x"0802d704",
			2212 => x"000022c1",
			2213 => x"ffbf22c1",
			2214 => x"000022c1",
			2215 => x"000022c1",
			2216 => x"000022c1",
			2217 => x"08035e0c",
			2218 => x"01010b04",
			2219 => x"000022c1",
			2220 => x"0003f304",
			2221 => x"000022c1",
			2222 => x"00b022c1",
			2223 => x"000022c1",
			2224 => x"040c4714",
			2225 => x"00039204",
			2226 => x"00002305",
			2227 => x"09024f0c",
			2228 => x"07073808",
			2229 => x"0802e304",
			2230 => x"00002305",
			2231 => x"ffb22305",
			2232 => x"00002305",
			2233 => x"00002305",
			2234 => x"08036e0c",
			2235 => x"01010b04",
			2236 => x"00002305",
			2237 => x"0003f104",
			2238 => x"00002305",
			2239 => x"00442305",
			2240 => x"00002305",
			2241 => x"040da91c",
			2242 => x"01016010",
			2243 => x"0802d804",
			2244 => x"00002351",
			2245 => x"040d0e08",
			2246 => x"00037d04",
			2247 => x"00002351",
			2248 => x"ffb42351",
			2249 => x"00002351",
			2250 => x"08035608",
			2251 => x"0d090104",
			2252 => x"00002351",
			2253 => x"006d2351",
			2254 => x"00002351",
			2255 => x"0a02dd08",
			2256 => x"0100e504",
			2257 => x"00002351",
			2258 => x"016f2351",
			2259 => x"00002351",
			2260 => x"040c471c",
			2261 => x"0b078210",
			2262 => x"00037d04",
			2263 => x"000023a5",
			2264 => x"09022b08",
			2265 => x"0706f604",
			2266 => x"ffa223a5",
			2267 => x"000023a5",
			2268 => x"000023a5",
			2269 => x"0a029608",
			2270 => x"06017d04",
			2271 => x"000023a5",
			2272 => x"000a23a5",
			2273 => x"000023a5",
			2274 => x"0a02dd0c",
			2275 => x"09016b04",
			2276 => x"000023a5",
			2277 => x"07068604",
			2278 => x"00e123a5",
			2279 => x"000023a5",
			2280 => x"000023a5",
			2281 => x"0c06de18",
			2282 => x"0a026a04",
			2283 => x"000023e1",
			2284 => x"09016b04",
			2285 => x"000023e1",
			2286 => x"0a02dd0c",
			2287 => x"09026b08",
			2288 => x"0c05d804",
			2289 => x"000023e1",
			2290 => x"003823e1",
			2291 => x"000023e1",
			2292 => x"000023e1",
			2293 => x"08034a04",
			2294 => x"000023e1",
			2295 => x"fe7623e1",
			2296 => x"040d551c",
			2297 => x"09020a04",
			2298 => x"ffb6242d",
			2299 => x"030b130c",
			2300 => x"0b07c308",
			2301 => x"0d08b304",
			2302 => x"0000242d",
			2303 => x"0077242d",
			2304 => x"0000242d",
			2305 => x"09024f08",
			2306 => x"08032504",
			2307 => x"0000242d",
			2308 => x"ffb6242d",
			2309 => x"0000242d",
			2310 => x"0a02dd08",
			2311 => x"06019404",
			2312 => x"0000242d",
			2313 => x"0184242d",
			2314 => x"0000242d",
			2315 => x"07076418",
			2316 => x"0c066d04",
			2317 => x"00002461",
			2318 => x"0601ca10",
			2319 => x"0e0a3904",
			2320 => x"00002461",
			2321 => x"020ae604",
			2322 => x"00002461",
			2323 => x"0a02dd04",
			2324 => x"003d2461",
			2325 => x"00002461",
			2326 => x"00002461",
			2327 => x"ffbb2461",
			2328 => x"0f0a6e10",
			2329 => x"0100e504",
			2330 => x"000024ad",
			2331 => x"020a1004",
			2332 => x"000024ad",
			2333 => x"01015704",
			2334 => x"00d324ad",
			2335 => x"000024ad",
			2336 => x"0802e304",
			2337 => x"000024ad",
			2338 => x"030aa904",
			2339 => x"000024ad",
			2340 => x"06018a04",
			2341 => x"000024ad",
			2342 => x"040b1404",
			2343 => x"000024ad",
			2344 => x"0a026104",
			2345 => x"000024ad",
			2346 => x"ffac24ad",
			2347 => x"0a028718",
			2348 => x"0a026404",
			2349 => x"00002501",
			2350 => x"0c063204",
			2351 => x"00002501",
			2352 => x"05091b0c",
			2353 => x"040b0404",
			2354 => x"00002501",
			2355 => x"01011504",
			2356 => x"00002501",
			2357 => x"012d2501",
			2358 => x"00002501",
			2359 => x"040d4208",
			2360 => x"08034704",
			2361 => x"00002501",
			2362 => x"ffae2501",
			2363 => x"0a02dd08",
			2364 => x"0a02bc04",
			2365 => x"00002501",
			2366 => x"00262501",
			2367 => x"00002501",
			2368 => x"040d1b20",
			2369 => x"0802e310",
			2370 => x"0b073304",
			2371 => x"0000255d",
			2372 => x"030b3208",
			2373 => x"01014304",
			2374 => x"0000255d",
			2375 => x"0082255d",
			2376 => x"0000255d",
			2377 => x"0101610c",
			2378 => x"040ce108",
			2379 => x"00039504",
			2380 => x"0000255d",
			2381 => x"ff67255d",
			2382 => x"0000255d",
			2383 => x"0000255d",
			2384 => x"08037c0c",
			2385 => x"00042e04",
			2386 => x"0000255d",
			2387 => x"0100f804",
			2388 => x"0000255d",
			2389 => x"00f7255d",
			2390 => x"ffd4255d",
			2391 => x"040c4720",
			2392 => x"0b078214",
			2393 => x"0802d804",
			2394 => x"000025b9",
			2395 => x"0101590c",
			2396 => x"0706f608",
			2397 => x"0a024f04",
			2398 => x"000025b9",
			2399 => x"ffa725b9",
			2400 => x"000025b9",
			2401 => x"000025b9",
			2402 => x"0a029608",
			2403 => x"06017d04",
			2404 => x"000025b9",
			2405 => x"000925b9",
			2406 => x"000025b9",
			2407 => x"08035e0c",
			2408 => x"0c061404",
			2409 => x"000025b9",
			2410 => x"0003f104",
			2411 => x"000025b9",
			2412 => x"00d725b9",
			2413 => x"000025b9",
			2414 => x"0b071e14",
			2415 => x"0c05d804",
			2416 => x"00002615",
			2417 => x"0003f304",
			2418 => x"00002615",
			2419 => x"0601a208",
			2420 => x"09016b04",
			2421 => x"00002615",
			2422 => x"00f02615",
			2423 => x"00002615",
			2424 => x"01015914",
			2425 => x"0802d804",
			2426 => x"00002615",
			2427 => x"030b230c",
			2428 => x"09022b08",
			2429 => x"05082e04",
			2430 => x"00002615",
			2431 => x"ff932615",
			2432 => x"00002615",
			2433 => x"00002615",
			2434 => x"08036504",
			2435 => x"00232615",
			2436 => x"00002615",
			2437 => x"0601b61c",
			2438 => x"09018b04",
			2439 => x"ffc92661",
			2440 => x"0c06dc14",
			2441 => x"06018e04",
			2442 => x"00002661",
			2443 => x"020b5b0c",
			2444 => x"0d097508",
			2445 => x"0601a104",
			2446 => x"00ce2661",
			2447 => x"00002661",
			2448 => x"00002661",
			2449 => x"00002661",
			2450 => x"00002661",
			2451 => x"08034704",
			2452 => x"00002661",
			2453 => x"0f0afc04",
			2454 => x"00002661",
			2455 => x"ff902661",
			2456 => x"0803471c",
			2457 => x"0d097518",
			2458 => x"020a8c04",
			2459 => x"000026ad",
			2460 => x"0c06ac10",
			2461 => x"0901bc04",
			2462 => x"000026ad",
			2463 => x"0e0bab08",
			2464 => x"0c063004",
			2465 => x"000026ad",
			2466 => x"008626ad",
			2467 => x"000026ad",
			2468 => x"000026ad",
			2469 => x"000026ad",
			2470 => x"020aa104",
			2471 => x"000026ad",
			2472 => x"0e0c8c04",
			2473 => x"ffdb26ad",
			2474 => x"000026ad",
			2475 => x"08030f1c",
			2476 => x"0b079310",
			2477 => x"0101590c",
			2478 => x"00039a04",
			2479 => x"00002721",
			2480 => x"0003c804",
			2481 => x"ffa42721",
			2482 => x"00002721",
			2483 => x"00002721",
			2484 => x"01016608",
			2485 => x"09020a04",
			2486 => x"00002721",
			2487 => x"00d42721",
			2488 => x"00002721",
			2489 => x"040c4c0c",
			2490 => x"09024f08",
			2491 => x"08032004",
			2492 => x"00002721",
			2493 => x"ff642721",
			2494 => x"00002721",
			2495 => x"08038110",
			2496 => x"0601c20c",
			2497 => x"0b068b04",
			2498 => x"00002721",
			2499 => x"0003f304",
			2500 => x"00002721",
			2501 => x"00582721",
			2502 => x"00002721",
			2503 => x"ffe72721",
			2504 => x"0e09510c",
			2505 => x"0100e504",
			2506 => x"0000277d",
			2507 => x"040c9304",
			2508 => x"0000277d",
			2509 => x"0202277d",
			2510 => x"0601900c",
			2511 => x"07068604",
			2512 => x"0000277d",
			2513 => x"0901fc04",
			2514 => x"0000277d",
			2515 => x"0014277d",
			2516 => x"0f0acb04",
			2517 => x"0000277d",
			2518 => x"01016110",
			2519 => x"0e0ae10c",
			2520 => x"0b072f04",
			2521 => x"0000277d",
			2522 => x"0802e304",
			2523 => x"0000277d",
			2524 => x"ff77277d",
			2525 => x"0000277d",
			2526 => x"0000277d",
			2527 => x"0f0a6e10",
			2528 => x"0d079604",
			2529 => x"000027d1",
			2530 => x"020a2d04",
			2531 => x"000027d1",
			2532 => x"06017c04",
			2533 => x"000027d1",
			2534 => x"001f27d1",
			2535 => x"0a026104",
			2536 => x"000027d1",
			2537 => x"0e0c8c14",
			2538 => x"0b071e04",
			2539 => x"000027d1",
			2540 => x"040b1404",
			2541 => x"000027d1",
			2542 => x"00039204",
			2543 => x"000027d1",
			2544 => x"030cdd04",
			2545 => x"ffc727d1",
			2546 => x"000027d1",
			2547 => x"000027d1",
			2548 => x"0e09510c",
			2549 => x"0100e504",
			2550 => x"00002835",
			2551 => x"040c9304",
			2552 => x"00002835",
			2553 => x"02552835",
			2554 => x"08036520",
			2555 => x"020ae610",
			2556 => x"00039504",
			2557 => x"00002835",
			2558 => x"0f0ad704",
			2559 => x"00002835",
			2560 => x"040b1404",
			2561 => x"00002835",
			2562 => x"ffa02835",
			2563 => x"0c063a04",
			2564 => x"00002835",
			2565 => x"040b3004",
			2566 => x"00002835",
			2567 => x"0c06dc04",
			2568 => x"00842835",
			2569 => x"00002835",
			2570 => x"0b070104",
			2571 => x"00002835",
			2572 => x"ff932835",
			2573 => x"01013f14",
			2574 => x"040d2e04",
			2575 => x"ff0c28a9",
			2576 => x"0803810c",
			2577 => x"00043904",
			2578 => x"000028a9",
			2579 => x"0100eb04",
			2580 => x"000028a9",
			2581 => x"008828a9",
			2582 => x"000028a9",
			2583 => x"030b530c",
			2584 => x"0c06aa08",
			2585 => x"07069b04",
			2586 => x"000028a9",
			2587 => x"00e728a9",
			2588 => x"000028a9",
			2589 => x"0c06a410",
			2590 => x"0f0b4a04",
			2591 => x"000028a9",
			2592 => x"0a027004",
			2593 => x"000028a9",
			2594 => x"01016904",
			2595 => x"ff6128a9",
			2596 => x"000028a9",
			2597 => x"01018a08",
			2598 => x"09021d04",
			2599 => x"000028a9",
			2600 => x"005b28a9",
			2601 => x"000028a9",
			2602 => x"040d5528",
			2603 => x"01015918",
			2604 => x"0706e114",
			2605 => x"040c4710",
			2606 => x"0802d804",
			2607 => x"0000290d",
			2608 => x"0b079508",
			2609 => x"0a025104",
			2610 => x"0000290d",
			2611 => x"ff4a290d",
			2612 => x"0000290d",
			2613 => x"0000290d",
			2614 => x"0000290d",
			2615 => x"0707280c",
			2616 => x"0706a104",
			2617 => x"0000290d",
			2618 => x"08034d04",
			2619 => x"0044290d",
			2620 => x"0000290d",
			2621 => x"0000290d",
			2622 => x"0a02dd08",
			2623 => x"06019104",
			2624 => x"0000290d",
			2625 => x"013d290d",
			2626 => x"0000290d",
			2627 => x"0c063a08",
			2628 => x"0a02cb04",
			2629 => x"ff882969",
			2630 => x"00002969",
			2631 => x"0d094110",
			2632 => x"05084d04",
			2633 => x"00002969",
			2634 => x"0c06c208",
			2635 => x"01012304",
			2636 => x"00002969",
			2637 => x"007e2969",
			2638 => x"00002969",
			2639 => x"07070c14",
			2640 => x"01015804",
			2641 => x"00002969",
			2642 => x"0c06a40c",
			2643 => x"0508dc04",
			2644 => x"00002969",
			2645 => x"0d094e04",
			2646 => x"00002969",
			2647 => x"ff812969",
			2648 => x"00002969",
			2649 => x"00002969",
			2650 => x"05080f10",
			2651 => x"0c05d804",
			2652 => x"000029d5",
			2653 => x"040c9304",
			2654 => x"000029d5",
			2655 => x"0803d004",
			2656 => x"01d929d5",
			2657 => x"000029d5",
			2658 => x"01015918",
			2659 => x"06018a04",
			2660 => x"000029d5",
			2661 => x"07068804",
			2662 => x"000029d5",
			2663 => x"09022b0c",
			2664 => x"0508f808",
			2665 => x"0802d804",
			2666 => x"000029d5",
			2667 => x"ff7729d5",
			2668 => x"000029d5",
			2669 => x"000029d5",
			2670 => x"0601ca0c",
			2671 => x"0706a104",
			2672 => x"000029d5",
			2673 => x"0a026204",
			2674 => x"000029d5",
			2675 => x"004d29d5",
			2676 => x"000029d5",
			2677 => x"0101492c",
			2678 => x"0902021c",
			2679 => x"0100f804",
			2680 => x"fe482a51",
			2681 => x"07067208",
			2682 => x"09019004",
			2683 => x"ffd92a51",
			2684 => x"fe512a51",
			2685 => x"0e0a700c",
			2686 => x"06018e04",
			2687 => x"fe572a51",
			2688 => x"0c066604",
			2689 => x"07252a51",
			2690 => x"00362a51",
			2691 => x"fe5d2a51",
			2692 => x"07069b08",
			2693 => x"0c063204",
			2694 => x"fe452a51",
			2695 => x"00002a51",
			2696 => x"06019f04",
			2697 => x"05612a51",
			2698 => x"004b2a51",
			2699 => x"0b072f04",
			2700 => x"fe4d2a51",
			2701 => x"0803680c",
			2702 => x"0706a104",
			2703 => x"01202a51",
			2704 => x"0c06de04",
			2705 => x"03832a51",
			2706 => x"023b2a51",
			2707 => x"fe5d2a51",
			2708 => x"0309d810",
			2709 => x"09016b04",
			2710 => x"00002ac5",
			2711 => x"040c9304",
			2712 => x"00002ac5",
			2713 => x"0c05a204",
			2714 => x"00002ac5",
			2715 => x"022b2ac5",
			2716 => x"06019014",
			2717 => x"0c063a04",
			2718 => x"00002ac5",
			2719 => x"0c06ac0c",
			2720 => x"0b073304",
			2721 => x"00002ac5",
			2722 => x"09020204",
			2723 => x"00002ac5",
			2724 => x"006e2ac5",
			2725 => x"00002ac5",
			2726 => x"0f0acb04",
			2727 => x"00002ac5",
			2728 => x"09023d10",
			2729 => x"0b072f04",
			2730 => x"00002ac5",
			2731 => x"0802e304",
			2732 => x"00002ac5",
			2733 => x"040b1404",
			2734 => x"00002ac5",
			2735 => x"ff932ac5",
			2736 => x"00002ac5",
			2737 => x"0f0a6e18",
			2738 => x"0100e504",
			2739 => x"00002b29",
			2740 => x"020a2d04",
			2741 => x"00002b29",
			2742 => x"06019f0c",
			2743 => x"06017c04",
			2744 => x"00002b29",
			2745 => x"09021d04",
			2746 => x"00282b29",
			2747 => x"00002b29",
			2748 => x"00002b29",
			2749 => x"0802e304",
			2750 => x"00002b29",
			2751 => x"0e0c8c14",
			2752 => x"0b071e04",
			2753 => x"00002b29",
			2754 => x"0a026104",
			2755 => x"00002b29",
			2756 => x"040b0204",
			2757 => x"00002b29",
			2758 => x"00039204",
			2759 => x"00002b29",
			2760 => x"ffb62b29",
			2761 => x"00002b29",
			2762 => x"0e0a2a18",
			2763 => x"0c05d804",
			2764 => x"00002ba5",
			2765 => x"0601ad10",
			2766 => x"020a2d04",
			2767 => x"00002ba5",
			2768 => x"06017804",
			2769 => x"00002ba5",
			2770 => x"0c066604",
			2771 => x"01052ba5",
			2772 => x"00002ba5",
			2773 => x"00002ba5",
			2774 => x"01015918",
			2775 => x"030b2314",
			2776 => x"0a025b04",
			2777 => x"00002ba5",
			2778 => x"09022b0c",
			2779 => x"0802d804",
			2780 => x"00002ba5",
			2781 => x"06018904",
			2782 => x"00002ba5",
			2783 => x"ff822ba5",
			2784 => x"00002ba5",
			2785 => x"00002ba5",
			2786 => x"0803610c",
			2787 => x"00039a04",
			2788 => x"00002ba5",
			2789 => x"0b074404",
			2790 => x"00002ba5",
			2791 => x"00402ba5",
			2792 => x"00002ba5",
			2793 => x"01014934",
			2794 => x"09020224",
			2795 => x"0100f804",
			2796 => x"fe4d2c31",
			2797 => x"0c063410",
			2798 => x"09019004",
			2799 => x"ffd82c31",
			2800 => x"0c061404",
			2801 => x"fe512c31",
			2802 => x"0c061504",
			2803 => x"ff812c31",
			2804 => x"fe792c31",
			2805 => x"0e0a700c",
			2806 => x"0901ce04",
			2807 => x"fe542c31",
			2808 => x"020ad604",
			2809 => x"fe962c31",
			2810 => x"048f2c31",
			2811 => x"fe602c31",
			2812 => x"0b072f08",
			2813 => x"0c063204",
			2814 => x"fe4a2c31",
			2815 => x"004f2c31",
			2816 => x"06019f04",
			2817 => x"03f22c31",
			2818 => x"004e2c31",
			2819 => x"0b072f04",
			2820 => x"fe522c31",
			2821 => x"0803680c",
			2822 => x"0c063a04",
			2823 => x"01012c31",
			2824 => x"0c06de04",
			2825 => x"02fa2c31",
			2826 => x"01ca2c31",
			2827 => x"fe672c31",
			2828 => x"0901fa10",
			2829 => x"020a9b04",
			2830 => x"fe6f2ccd",
			2831 => x"020b0f08",
			2832 => x"040c6004",
			2833 => x"ffc12ccd",
			2834 => x"00d62ccd",
			2835 => x"fec82ccd",
			2836 => x"040b6328",
			2837 => x"0b077110",
			2838 => x"0a025704",
			2839 => x"00002ccd",
			2840 => x"01015a08",
			2841 => x"01014504",
			2842 => x"00002ccd",
			2843 => x"fe472ccd",
			2844 => x"00002ccd",
			2845 => x"030b1304",
			2846 => x"01732ccd",
			2847 => x"0e0ac908",
			2848 => x"0e0ac404",
			2849 => x"00002ccd",
			2850 => x"fdbf2ccd",
			2851 => x"0706df04",
			2852 => x"ff3a2ccd",
			2853 => x"040b3004",
			2854 => x"ffce2ccd",
			2855 => x"011a2ccd",
			2856 => x"0a02a90c",
			2857 => x"0b071004",
			2858 => x"00002ccd",
			2859 => x"0b07e604",
			2860 => x"01732ccd",
			2861 => x"00002ccd",
			2862 => x"040c8504",
			2863 => x"fede2ccd",
			2864 => x"08036e04",
			2865 => x"01482ccd",
			2866 => x"ff402ccd",
			2867 => x"09018b04",
			2868 => x"ff682d49",
			2869 => x"0f0b2d20",
			2870 => x"0b07b514",
			2871 => x"0601b210",
			2872 => x"0802e504",
			2873 => x"00002d49",
			2874 => x"020a8304",
			2875 => x"00002d49",
			2876 => x"0c05d804",
			2877 => x"00002d49",
			2878 => x"00c42d49",
			2879 => x"00002d49",
			2880 => x"06019104",
			2881 => x"00002d49",
			2882 => x"0802eb04",
			2883 => x"ffda2d49",
			2884 => x"00002d49",
			2885 => x"09024f10",
			2886 => x"0707380c",
			2887 => x"0e0b0704",
			2888 => x"00002d49",
			2889 => x"06018a04",
			2890 => x"00002d49",
			2891 => x"ff402d49",
			2892 => x"00002d49",
			2893 => x"0601ca08",
			2894 => x"0c067304",
			2895 => x"00002d49",
			2896 => x"00892d49",
			2897 => x"00002d49",
			2898 => x"09020520",
			2899 => x"06018a08",
			2900 => x"09020204",
			2901 => x"fe642e05",
			2902 => x"00002e05",
			2903 => x"0e0a7014",
			2904 => x"040c2404",
			2905 => x"fe902e05",
			2906 => x"06019908",
			2907 => x"0c05f604",
			2908 => x"ff292e05",
			2909 => x"02732e05",
			2910 => x"0901dd04",
			2911 => x"fe892e05",
			2912 => x"009f2e05",
			2913 => x"fe6d2e05",
			2914 => x"0b07631c",
			2915 => x"040b6310",
			2916 => x"06018908",
			2917 => x"05084d04",
			2918 => x"fedb2e05",
			2919 => x"016c2e05",
			2920 => x"01015704",
			2921 => x"fe112e05",
			2922 => x"ff802e05",
			2923 => x"0e0a9c04",
			2924 => x"02a12e05",
			2925 => x"09022e04",
			2926 => x"fec32e05",
			2927 => x"000a2e05",
			2928 => x"0b07b510",
			2929 => x"0601bc0c",
			2930 => x"0c06ac04",
			2931 => x"01a52e05",
			2932 => x"0c06ae04",
			2933 => x"00002e05",
			2934 => x"01762e05",
			2935 => x"ffae2e05",
			2936 => x"00039a08",
			2937 => x"0f0afc04",
			2938 => x"01552e05",
			2939 => x"fe022e05",
			2940 => x"0e0ab804",
			2941 => x"fee52e05",
			2942 => x"0601ca04",
			2943 => x"019f2e05",
			2944 => x"fec12e05",
			2945 => x"0901ce04",
			2946 => x"ff042e89",
			2947 => x"0f0b1720",
			2948 => x"020aaf10",
			2949 => x"0706c90c",
			2950 => x"0802d804",
			2951 => x"00002e89",
			2952 => x"0003e104",
			2953 => x"ff862e89",
			2954 => x"00002e89",
			2955 => x"00002e89",
			2956 => x"0706e00c",
			2957 => x"0601b708",
			2958 => x"0d087f04",
			2959 => x"00002e89",
			2960 => x"00d52e89",
			2961 => x"00002e89",
			2962 => x"00002e89",
			2963 => x"0706df10",
			2964 => x"09023f0c",
			2965 => x"040c6608",
			2966 => x"01016704",
			2967 => x"ff1e2e89",
			2968 => x"00002e89",
			2969 => x"00002e89",
			2970 => x"00002e89",
			2971 => x"0803610c",
			2972 => x"040b3c04",
			2973 => x"00002e89",
			2974 => x"01014704",
			2975 => x"00002e89",
			2976 => x"00c42e89",
			2977 => x"00002e89",
			2978 => x"0901fa14",
			2979 => x"06018a04",
			2980 => x"fe702f35",
			2981 => x"0f0a9e0c",
			2982 => x"0c05d804",
			2983 => x"00002f35",
			2984 => x"040c1804",
			2985 => x"00002f35",
			2986 => x"00ba2f35",
			2987 => x"fecd2f35",
			2988 => x"040b6328",
			2989 => x"0b077110",
			2990 => x"06018908",
			2991 => x"05084d04",
			2992 => x"00002f35",
			2993 => x"00912f35",
			2994 => x"01015a04",
			2995 => x"fe4d2f35",
			2996 => x"00002f35",
			2997 => x"0f0b0304",
			2998 => x"016e2f35",
			2999 => x"09022a08",
			3000 => x"0c06aa04",
			3001 => x"00f92f35",
			3002 => x"fff02f35",
			3003 => x"0802eb08",
			3004 => x"0d094e04",
			3005 => x"00002f35",
			3006 => x"fdf92f35",
			3007 => x"00562f35",
			3008 => x"0601b20c",
			3009 => x"0b071004",
			3010 => x"00002f35",
			3011 => x"0f0be504",
			3012 => x"016a2f35",
			3013 => x"00002f35",
			3014 => x"09023004",
			3015 => x"fee42f35",
			3016 => x"0601cc08",
			3017 => x"0c067004",
			3018 => x"00002f35",
			3019 => x"01602f35",
			3020 => x"ff2e2f35",
			3021 => x"0004a740",
			3022 => x"040d2e30",
			3023 => x"0706c910",
			3024 => x"0802d804",
			3025 => x"00002fc9",
			3026 => x"09023b08",
			3027 => x"0c068904",
			3028 => x"ff832fc9",
			3029 => x"00002fc9",
			3030 => x"00002fc9",
			3031 => x"0c06a110",
			3032 => x"0901e804",
			3033 => x"00002fc9",
			3034 => x"07072208",
			3035 => x"0706ca04",
			3036 => x"00002fc9",
			3037 => x"007c2fc9",
			3038 => x"00002fc9",
			3039 => x"0a027004",
			3040 => x"00002fc9",
			3041 => x"040b6904",
			3042 => x"00002fc9",
			3043 => x"020bf304",
			3044 => x"ffc32fc9",
			3045 => x"00002fc9",
			3046 => x"0803810c",
			3047 => x"00042e04",
			3048 => x"00002fc9",
			3049 => x"09018b04",
			3050 => x"00002fc9",
			3051 => x"00b52fc9",
			3052 => x"00002fc9",
			3053 => x"0004ab08",
			3054 => x"040d1b04",
			3055 => x"00002fc9",
			3056 => x"03612fc9",
			3057 => x"00002fc9",
			3058 => x"01014934",
			3059 => x"09020e2c",
			3060 => x"09020220",
			3061 => x"0100f804",
			3062 => x"fe43306d",
			3063 => x"0c06330c",
			3064 => x"09019004",
			3065 => x"ffba306d",
			3066 => x"0901bf04",
			3067 => x"fe96306d",
			3068 => x"fe48306d",
			3069 => x"0e09fd08",
			3070 => x"0901ce04",
			3071 => x"fe56306d",
			3072 => x"03b1306d",
			3073 => x"0901fa04",
			3074 => x"fe5a306d",
			3075 => x"ff6d306d",
			3076 => x"0c065008",
			3077 => x"05082e04",
			3078 => x"fe49306d",
			3079 => x"0066306d",
			3080 => x"0381306d",
			3081 => x"06018d04",
			3082 => x"0479306d",
			3083 => x"fe6e306d",
			3084 => x"0d08b308",
			3085 => x"040bcc04",
			3086 => x"fe47306d",
			3087 => x"0000306d",
			3088 => x"0a02c710",
			3089 => x"0c063a04",
			3090 => x"021a306d",
			3091 => x"0706a104",
			3092 => x"02df306d",
			3093 => x"0c06de04",
			3094 => x"046a306d",
			3095 => x"0321306d",
			3096 => x"07072604",
			3097 => x"fe6c306d",
			3098 => x"00e8306d",
			3099 => x"0101492c",
			3100 => x"0100f80c",
			3101 => x"0100e504",
			3102 => x"fe603131",
			3103 => x"0100e704",
			3104 => x"00833131",
			3105 => x"fe6f3131",
			3106 => x"040c6014",
			3107 => x"0706b708",
			3108 => x"05088604",
			3109 => x"fe5d3131",
			3110 => x"ffeb3131",
			3111 => x"06019408",
			3112 => x"01013b04",
			3113 => x"fee93131",
			3114 => x"01cc3131",
			3115 => x"fe763131",
			3116 => x"020b4904",
			3117 => x"02ec3131",
			3118 => x"0601a904",
			3119 => x"01103131",
			3120 => x"fe753131",
			3121 => x"0c063a0c",
			3122 => x"06019e08",
			3123 => x"0f0abc04",
			3124 => x"fe0a3131",
			3125 => x"00fe3131",
			3126 => x"fe383131",
			3127 => x"0601c224",
			3128 => x"0b07630c",
			3129 => x"0c066c08",
			3130 => x"0802f804",
			3131 => x"019b3131",
			3132 => x"fe883131",
			3133 => x"02093131",
			3134 => x"0601ad10",
			3135 => x"0d097508",
			3136 => x"0b077104",
			3137 => x"01383131",
			3138 => x"01b63131",
			3139 => x"0d097704",
			3140 => x"00003131",
			3141 => x"01b53131",
			3142 => x"01016c04",
			3143 => x"ff3f3131",
			3144 => x"01d03131",
			3145 => x"00045404",
			3146 => x"fef43131",
			3147 => x"00433131",
			3148 => x"040d1b3c",
			3149 => x"08034734",
			3150 => x"040b6b20",
			3151 => x"0802e310",
			3152 => x"0706a104",
			3153 => x"000031c5",
			3154 => x"030b2a08",
			3155 => x"01014304",
			3156 => x"000031c5",
			3157 => x"007931c5",
			3158 => x"000031c5",
			3159 => x"0c06a40c",
			3160 => x"07072408",
			3161 => x"09023904",
			3162 => x"ff6631c5",
			3163 => x"000031c5",
			3164 => x"000031c5",
			3165 => x"000031c5",
			3166 => x"0c063204",
			3167 => x"000031c5",
			3168 => x"0c06dc0c",
			3169 => x"0e0bc508",
			3170 => x"01012304",
			3171 => x"000031c5",
			3172 => x"009731c5",
			3173 => x"000031c5",
			3174 => x"000031c5",
			3175 => x"020bf304",
			3176 => x"ff2131c5",
			3177 => x"000031c5",
			3178 => x"08037c0c",
			3179 => x"00042e04",
			3180 => x"000031c5",
			3181 => x"0100f804",
			3182 => x"000031c5",
			3183 => x"00ee31c5",
			3184 => x"ffd931c5",
			3185 => x"020a830c",
			3186 => x"0802d804",
			3187 => x"00003279",
			3188 => x"05086a04",
			3189 => x"fed63279",
			3190 => x"00003279",
			3191 => x"0e0aa220",
			3192 => x"01012310",
			3193 => x"020ad10c",
			3194 => x"040d2e04",
			3195 => x"00003279",
			3196 => x"06017c04",
			3197 => x"00003279",
			3198 => x"006a3279",
			3199 => x"ff783279",
			3200 => x"0c06a10c",
			3201 => x"0d087404",
			3202 => x"00003279",
			3203 => x"0c063004",
			3204 => x"00003279",
			3205 => x"00e03279",
			3206 => x"00003279",
			3207 => x"0706f514",
			3208 => x"01015c0c",
			3209 => x"0b079308",
			3210 => x"00039504",
			3211 => x"00003279",
			3212 => x"fed63279",
			3213 => x"00003279",
			3214 => x"08033c04",
			3215 => x"000c3279",
			3216 => x"00003279",
			3217 => x"030b5b0c",
			3218 => x"040b1504",
			3219 => x"00003279",
			3220 => x"01014304",
			3221 => x"00003279",
			3222 => x"00ac3279",
			3223 => x"0101790c",
			3224 => x"0a027004",
			3225 => x"00003279",
			3226 => x"0c06a104",
			3227 => x"00003279",
			3228 => x"ff7e3279",
			3229 => x"00003279",
			3230 => x"01014928",
			3231 => x"0100f804",
			3232 => x"fe613325",
			3233 => x"040c6014",
			3234 => x"0706b708",
			3235 => x"05088604",
			3236 => x"fe5b3325",
			3237 => x"ffdf3325",
			3238 => x"0901fa04",
			3239 => x"fe823325",
			3240 => x"0508a504",
			3241 => x"01df3325",
			3242 => x"00003325",
			3243 => x"0508b30c",
			3244 => x"08037f08",
			3245 => x"0b071e04",
			3246 => x"03a73325",
			3247 => x"01ef3325",
			3248 => x"00003325",
			3249 => x"fe7b3325",
			3250 => x"0c063a0c",
			3251 => x"0a027a08",
			3252 => x"040b2e04",
			3253 => x"fe063325",
			3254 => x"01153325",
			3255 => x"fe2d3325",
			3256 => x"08037320",
			3257 => x"0101500c",
			3258 => x"0a026904",
			3259 => x"01c23325",
			3260 => x"0e0aa204",
			3261 => x"01843325",
			3262 => x"fdbd3325",
			3263 => x"0d095004",
			3264 => x"01c43325",
			3265 => x"00039d08",
			3266 => x"0f0afc04",
			3267 => x"019b3325",
			3268 => x"fe913325",
			3269 => x"0a02a904",
			3270 => x"01c63325",
			3271 => x"008f3325",
			3272 => x"fea93325",
			3273 => x"0100f804",
			3274 => x"fec233a9",
			3275 => x"020b5b34",
			3276 => x"0508dc1c",
			3277 => x"09021214",
			3278 => x"040c600c",
			3279 => x"0802e904",
			3280 => x"000033a9",
			3281 => x"0706e304",
			3282 => x"ff4633a9",
			3283 => x"000033a9",
			3284 => x"07069b04",
			3285 => x"00d833a9",
			3286 => x"000033a9",
			3287 => x"0d08b304",
			3288 => x"000033a9",
			3289 => x"012833a9",
			3290 => x"0c068d10",
			3291 => x"09022a04",
			3292 => x"000033a9",
			3293 => x"0a026708",
			3294 => x"0d094e04",
			3295 => x"000033a9",
			3296 => x"fed533a9",
			3297 => x"000033a9",
			3298 => x"0003c404",
			3299 => x"00a933a9",
			3300 => x"000033a9",
			3301 => x"08031204",
			3302 => x"000033a9",
			3303 => x"01016d04",
			3304 => x"ff4333a9",
			3305 => x"000033a9",
			3306 => x"020a1004",
			3307 => x"fe893425",
			3308 => x"040d4230",
			3309 => x"0a02b424",
			3310 => x"0101601c",
			3311 => x"0003950c",
			3312 => x"0706a104",
			3313 => x"00003425",
			3314 => x"01014704",
			3315 => x"00003425",
			3316 => x"010e3425",
			3317 => x"040b6308",
			3318 => x"0706f504",
			3319 => x"ff073425",
			3320 => x"00003425",
			3321 => x"0a028d04",
			3322 => x"00b13425",
			3323 => x"00003425",
			3324 => x"0d08f404",
			3325 => x"00003425",
			3326 => x"012c3425",
			3327 => x"020a8604",
			3328 => x"00003425",
			3329 => x"08034804",
			3330 => x"00003425",
			3331 => x"ff013425",
			3332 => x"0a02dd08",
			3333 => x"03088d04",
			3334 => x"00003425",
			3335 => x"01b23425",
			3336 => x"ffcf3425",
			3337 => x"09020224",
			3338 => x"06018a04",
			3339 => x"fe643501",
			3340 => x"0601960c",
			3341 => x"040c2404",
			3342 => x"feb43501",
			3343 => x"0c05d804",
			3344 => x"ff503501",
			3345 => x"024f3501",
			3346 => x"0901ce04",
			3347 => x"fe603501",
			3348 => x"040ce10c",
			3349 => x"0901df08",
			3350 => x"0901dd04",
			3351 => x"ffcc3501",
			3352 => x"00003501",
			3353 => x"fe753501",
			3354 => x"012c3501",
			3355 => x"0b077124",
			3356 => x"0e0aa214",
			3357 => x"040b8a10",
			3358 => x"05086a08",
			3359 => x"06018304",
			3360 => x"001e3501",
			3361 => x"fe463501",
			3362 => x"09021204",
			3363 => x"00003501",
			3364 => x"01793501",
			3365 => x"02963501",
			3366 => x"0e0aa404",
			3367 => x"f44d3501",
			3368 => x"0c066c08",
			3369 => x"09022d04",
			3370 => x"fe043501",
			3371 => x"ff6f3501",
			3372 => x"019a3501",
			3373 => x"0d094e10",
			3374 => x"0c06c208",
			3375 => x"0e0b6304",
			3376 => x"01a13501",
			3377 => x"00003501",
			3378 => x"0b07b104",
			3379 => x"00fd3501",
			3380 => x"ff933501",
			3381 => x"0706f508",
			3382 => x"0a026704",
			3383 => x"f92e3501",
			3384 => x"005f3501",
			3385 => x"0601cc0c",
			3386 => x"0e0ae108",
			3387 => x"07072204",
			3388 => x"018c3501",
			3389 => x"fee03501",
			3390 => x"01a33501",
			3391 => x"feef3501",
			3392 => x"0c06140c",
			3393 => x"020a9b04",
			3394 => x"fe6935bd",
			3395 => x"020aa104",
			3396 => x"009635bd",
			3397 => x"feb835bd",
			3398 => x"01015c40",
			3399 => x"030b1324",
			3400 => x"0901bc0c",
			3401 => x"0c061708",
			3402 => x"0100fa04",
			3403 => x"000035bd",
			3404 => x"005035bd",
			3405 => x"fec135bd",
			3406 => x"06018c08",
			3407 => x"0f0a4204",
			3408 => x"000035bd",
			3409 => x"019435bd",
			3410 => x"040bd808",
			3411 => x"01014f04",
			3412 => x"fea735bd",
			3413 => x"008c35bd",
			3414 => x"0601b204",
			3415 => x"016935bd",
			3416 => x"000035bd",
			3417 => x"0706f510",
			3418 => x"09021808",
			3419 => x"06019f04",
			3420 => x"002a35bd",
			3421 => x"000035bd",
			3422 => x"09022a04",
			3423 => x"fe9135bd",
			3424 => x"fc7d35bd",
			3425 => x"0a02a908",
			3426 => x"01014704",
			3427 => x"000035bd",
			3428 => x"015e35bd",
			3429 => x"feb535bd",
			3430 => x"0a026408",
			3431 => x"09023704",
			3432 => x"014235bd",
			3433 => x"fea035bd",
			3434 => x"0601c208",
			3435 => x"0d090104",
			3436 => x"000035bd",
			3437 => x"019235bd",
			3438 => x"002b35bd",
			3439 => x"09018b04",
			3440 => x"fe753659",
			3441 => x"0601a530",
			3442 => x"040b6320",
			3443 => x"05086a04",
			3444 => x"fee43659",
			3445 => x"0f0aed0c",
			3446 => x"01013f04",
			3447 => x"00003659",
			3448 => x"0802f804",
			3449 => x"015a3659",
			3450 => x"00003659",
			3451 => x"0a026c08",
			3452 => x"06019104",
			3453 => x"00003659",
			3454 => x"fea93659",
			3455 => x"0508a404",
			3456 => x"00003659",
			3457 => x"00b83659",
			3458 => x"020b7708",
			3459 => x"020a9b04",
			3460 => x"00003659",
			3461 => x"01463659",
			3462 => x"01016704",
			3463 => x"ffbb3659",
			3464 => x"00003659",
			3465 => x"040c5e0c",
			3466 => x"09024f08",
			3467 => x"0a028b04",
			3468 => x"00003659",
			3469 => x"fea43659",
			3470 => x"00003659",
			3471 => x"08036508",
			3472 => x"01014704",
			3473 => x"00003659",
			3474 => x"00fd3659",
			3475 => x"0601be04",
			3476 => x"002e3659",
			3477 => x"fee23659",
			3478 => x"0c05d804",
			3479 => x"ff1b36e5",
			3480 => x"040c8530",
			3481 => x"06018c0c",
			3482 => x"01013f04",
			3483 => x"000036e5",
			3484 => x"0b071004",
			3485 => x"000036e5",
			3486 => x"008936e5",
			3487 => x"01015008",
			3488 => x"0f0a8a04",
			3489 => x"000036e5",
			3490 => x"ff3b36e5",
			3491 => x"0802ee10",
			3492 => x"0b07b508",
			3493 => x"0802e004",
			3494 => x"ffd936e5",
			3495 => x"004b36e5",
			3496 => x"0802e804",
			3497 => x"000036e5",
			3498 => x"ff9836e5",
			3499 => x"020b7708",
			3500 => x"05086a04",
			3501 => x"000036e5",
			3502 => x"007f36e5",
			3503 => x"000036e5",
			3504 => x"0a02db10",
			3505 => x"0100f804",
			3506 => x"000036e5",
			3507 => x"0d08f404",
			3508 => x"00df36e5",
			3509 => x"0d097704",
			3510 => x"000036e5",
			3511 => x"004936e5",
			3512 => x"000036e5",
			3513 => x"09020828",
			3514 => x"020a2d04",
			3515 => x"fe6137a1",
			3516 => x"0601a520",
			3517 => x"040c240c",
			3518 => x"0c066604",
			3519 => x"fe5f37a1",
			3520 => x"0706c904",
			3521 => x"00b337a1",
			3522 => x"fef737a1",
			3523 => x"09016b04",
			3524 => x"fe9337a1",
			3525 => x"020b1f08",
			3526 => x"07061304",
			3527 => x"ff9137a1",
			3528 => x"037037a1",
			3529 => x"01012304",
			3530 => x"fe6f37a1",
			3531 => x"020137a1",
			3532 => x"fe6337a1",
			3533 => x"0c063a08",
			3534 => x"05086a04",
			3535 => x"fe4437a1",
			3536 => x"00c337a1",
			3537 => x"0803261c",
			3538 => x"0d097514",
			3539 => x"0b076308",
			3540 => x"01014f04",
			3541 => x"ff5a37a1",
			3542 => x"01b537a1",
			3543 => x"0d094e04",
			3544 => x"01b037a1",
			3545 => x"0b079304",
			3546 => x"ff4037a1",
			3547 => x"017d37a1",
			3548 => x"040b7004",
			3549 => x"feaf37a1",
			3550 => x"019e37a1",
			3551 => x"040c4708",
			3552 => x"01016c04",
			3553 => x"fdb937a1",
			3554 => x"00dc37a1",
			3555 => x"08036e08",
			3556 => x"08033404",
			3557 => x"003537a1",
			3558 => x"01e137a1",
			3559 => x"fec637a1",
			3560 => x"09020824",
			3561 => x"020a2d04",
			3562 => x"fe613855",
			3563 => x"0601a51c",
			3564 => x"040c240c",
			3565 => x"0c066604",
			3566 => x"fe5c3855",
			3567 => x"0706c904",
			3568 => x"00c63855",
			3569 => x"feec3855",
			3570 => x"09016b04",
			3571 => x"fe8b3855",
			3572 => x"0308b604",
			3573 => x"0a263855",
			3574 => x"020b5b04",
			3575 => x"02ad3855",
			3576 => x"005e3855",
			3577 => x"fe623855",
			3578 => x"05086a08",
			3579 => x"0c063a04",
			3580 => x"fe433855",
			3581 => x"00f13855",
			3582 => x"0601b724",
			3583 => x"0f0bae1c",
			3584 => x"0b07b50c",
			3585 => x"040c2c08",
			3586 => x"09021204",
			3587 => x"00e83855",
			3588 => x"01ae3855",
			3589 => x"02793855",
			3590 => x"0003a208",
			3591 => x"09022e04",
			3592 => x"01a13855",
			3593 => x"fe3e3855",
			3594 => x"0d094904",
			3595 => x"00003855",
			3596 => x"01b23855",
			3597 => x"0508de04",
			3598 => x"fe7d3855",
			3599 => x"01993855",
			3600 => x"01017704",
			3601 => x"fd773855",
			3602 => x"0601c604",
			3603 => x"01be3855",
			3604 => x"00003855",
			3605 => x"0c06140c",
			3606 => x"040dca04",
			3607 => x"fe753929",
			3608 => x"040df504",
			3609 => x"00003929",
			3610 => x"ff773929",
			3611 => x"0b07b53c",
			3612 => x"0c066c24",
			3613 => x"0706830c",
			3614 => x"040b8e04",
			3615 => x"00003929",
			3616 => x"0f0afc04",
			3617 => x"01543929",
			3618 => x"00003929",
			3619 => x"0706ca0c",
			3620 => x"0c061604",
			3621 => x"00003929",
			3622 => x"0802d804",
			3623 => x"00003929",
			3624 => x"fee73929",
			3625 => x"0b076304",
			3626 => x"00003929",
			3627 => x"0601a704",
			3628 => x"007e3929",
			3629 => x"00003929",
			3630 => x"09020208",
			3631 => x"0c066e04",
			3632 => x"00003929",
			3633 => x"ff923929",
			3634 => x"0e0b0704",
			3635 => x"016a3929",
			3636 => x"030b4104",
			3637 => x"ff953929",
			3638 => x"0f0be504",
			3639 => x"00793929",
			3640 => x"00003929",
			3641 => x"0c06a410",
			3642 => x"030b2a04",
			3643 => x"00003929",
			3644 => x"0b07c308",
			3645 => x"020b2c04",
			3646 => x"fe243929",
			3647 => x"00003929",
			3648 => x"00003929",
			3649 => x"0e0ac908",
			3650 => x"07071204",
			3651 => x"00003929",
			3652 => x"fef53929",
			3653 => x"0601ca08",
			3654 => x"09021d04",
			3655 => x"00003929",
			3656 => x"01563929",
			3657 => x"ff523929",
			3658 => x"01013f1c",
			3659 => x"06018a04",
			3660 => x"fe6539d5",
			3661 => x"030a8110",
			3662 => x"040c6004",
			3663 => x"fe9139d5",
			3664 => x"0706a108",
			3665 => x"0c05d804",
			3666 => x"fef839d5",
			3667 => x"021539d5",
			3668 => x"ff8839d5",
			3669 => x"06019404",
			3670 => x"fffc39d5",
			3671 => x"fe6b39d5",
			3672 => x"0c063004",
			3673 => x"fe9439d5",
			3674 => x"06018a08",
			3675 => x"0003ab04",
			3676 => x"019a39d5",
			3677 => x"042d39d5",
			3678 => x"01015918",
			3679 => x"0706e210",
			3680 => x"040b6308",
			3681 => x"0b078204",
			3682 => x"fd5939d5",
			3683 => x"000039d5",
			3684 => x"0e0aee04",
			3685 => x"017a39d5",
			3686 => x"feaf39d5",
			3687 => x"06019a04",
			3688 => x"018c39d5",
			3689 => x"feda39d5",
			3690 => x"0b07b50c",
			3691 => x"0e0bab08",
			3692 => x"0d08f404",
			3693 => x"005139d5",
			3694 => x"019e39d5",
			3695 => x"ff7039d5",
			3696 => x"0a026404",
			3697 => x"fd3039d5",
			3698 => x"0601cc04",
			3699 => x"015539d5",
			3700 => x"ff0539d5",
			3701 => x"020a5b08",
			3702 => x"05088604",
			3703 => x"fe8e3aa1",
			3704 => x"00003aa1",
			3705 => x"030b2a38",
			3706 => x"01015024",
			3707 => x"0f0ab214",
			3708 => x"0706830c",
			3709 => x"040b8e04",
			3710 => x"00003aa1",
			3711 => x"0100f804",
			3712 => x"00003aa1",
			3713 => x"00f83aa1",
			3714 => x"05086a04",
			3715 => x"ffac3aa1",
			3716 => x"00003aa1",
			3717 => x"030ae50c",
			3718 => x"040d0008",
			3719 => x"020aa104",
			3720 => x"00003aa1",
			3721 => x"ff093aa1",
			3722 => x"00003aa1",
			3723 => x"00003aa1",
			3724 => x"0707250c",
			3725 => x"0f0b5108",
			3726 => x"0d08b304",
			3727 => x"00003aa1",
			3728 => x"01513aa1",
			3729 => x"00003aa1",
			3730 => x"0508d104",
			3731 => x"00003aa1",
			3732 => x"fff73aa1",
			3733 => x"0003a20c",
			3734 => x"09021d04",
			3735 => x"00003aa1",
			3736 => x"0d095004",
			3737 => x"00003aa1",
			3738 => x"feae3aa1",
			3739 => x"040c1208",
			3740 => x"01014904",
			3741 => x"00003aa1",
			3742 => x"00e43aa1",
			3743 => x"09025208",
			3744 => x"0e0b1604",
			3745 => x"00003aa1",
			3746 => x"fef13aa1",
			3747 => x"08036e08",
			3748 => x"0c068804",
			3749 => x"00003aa1",
			3750 => x"00e53aa1",
			3751 => x"ffef3aa1",
			3752 => x"0c061410",
			3753 => x"040dca04",
			3754 => x"fe793b75",
			3755 => x"040df508",
			3756 => x"06017404",
			3757 => x"00003b75",
			3758 => x"002a3b75",
			3759 => x"ffa03b75",
			3760 => x"0b07b540",
			3761 => x"0c066c24",
			3762 => x"020b7720",
			3763 => x"040b6310",
			3764 => x"05086a08",
			3765 => x"06017d04",
			3766 => x"00003b75",
			3767 => x"fec93b75",
			3768 => x"0a027404",
			3769 => x"005e3b75",
			3770 => x"ffef3b75",
			3771 => x"06019908",
			3772 => x"020b2c04",
			3773 => x"013d3b75",
			3774 => x"00003b75",
			3775 => x"01013404",
			3776 => x"ffa63b75",
			3777 => x"002e3b75",
			3778 => x"feda3b75",
			3779 => x"01013508",
			3780 => x"0c066e04",
			3781 => x"00003b75",
			3782 => x"ffb13b75",
			3783 => x"0e0b0708",
			3784 => x"0d095e04",
			3785 => x"01613b75",
			3786 => x"00003b75",
			3787 => x"030b4104",
			3788 => x"ffa63b75",
			3789 => x"0f0be504",
			3790 => x"00613b75",
			3791 => x"00003b75",
			3792 => x"01016010",
			3793 => x"06018e04",
			3794 => x"00003b75",
			3795 => x"0e0b0e08",
			3796 => x"05090a04",
			3797 => x"fe733b75",
			3798 => x"00003b75",
			3799 => x"00003b75",
			3800 => x"0601ca08",
			3801 => x"0c068d04",
			3802 => x"00003b75",
			3803 => x"01343b75",
			3804 => x"ff5f3b75",
			3805 => x"0901fa28",
			3806 => x"06018a04",
			3807 => x"fe663c69",
			3808 => x"0f0aa618",
			3809 => x"0c05d804",
			3810 => x"fef53c69",
			3811 => x"0f0a6e08",
			3812 => x"0a028804",
			3813 => x"00003c69",
			3814 => x"01bf3c69",
			3815 => x"0f0a9208",
			3816 => x"06019404",
			3817 => x"00003c69",
			3818 => x"ff493c69",
			3819 => x"00b33c69",
			3820 => x"0d08b308",
			3821 => x"0d088204",
			3822 => x"fef63c69",
			3823 => x"00003c69",
			3824 => x"fe713c69",
			3825 => x"0101502c",
			3826 => x"0e0a8418",
			3827 => x"030a3908",
			3828 => x"08031b04",
			3829 => x"feb43c69",
			3830 => x"00003c69",
			3831 => x"07070d0c",
			3832 => x"020aad08",
			3833 => x"0706a104",
			3834 => x"fea93c69",
			3835 => x"016c3c69",
			3836 => x"01f73c69",
			3837 => x"ff6a3c69",
			3838 => x"0a026904",
			3839 => x"011e3c69",
			3840 => x"09020e0c",
			3841 => x"09020504",
			3842 => x"feda3c69",
			3843 => x"020b5304",
			3844 => x"00003c69",
			3845 => x"00043c69",
			3846 => x"fdc13c69",
			3847 => x"08034d20",
			3848 => x"0d097518",
			3849 => x"0706a10c",
			3850 => x"0e0a9a08",
			3851 => x"020ab704",
			3852 => x"00003c69",
			3853 => x"010d3c69",
			3854 => x"feec3c69",
			3855 => x"07073808",
			3856 => x"0c06ac04",
			3857 => x"019b3c69",
			3858 => x"00cf3c69",
			3859 => x"00003c69",
			3860 => x"020b2404",
			3861 => x"febc3c69",
			3862 => x"01813c69",
			3863 => x"0706f904",
			3864 => x"fea73c69",
			3865 => x"00003c69",
			3866 => x"0c05f604",
			3867 => x"fe6c3d0d",
			3868 => x"0101593c",
			3869 => x"040c472c",
			3870 => x"0b078218",
			3871 => x"0e0aa210",
			3872 => x"0c065008",
			3873 => x"040ba404",
			3874 => x"fe893d0d",
			3875 => x"00003d0d",
			3876 => x"0d08b304",
			3877 => x"00003d0d",
			3878 => x"00e13d0d",
			3879 => x"0c068704",
			3880 => x"fe113d0d",
			3881 => x"00003d0d",
			3882 => x"0c06ac08",
			3883 => x"09020804",
			3884 => x"00003d0d",
			3885 => x"01663d0d",
			3886 => x"0e0ae708",
			3887 => x"040b4604",
			3888 => x"00003d0d",
			3889 => x"feab3d0d",
			3890 => x"00003d0d",
			3891 => x"0601b20c",
			3892 => x"0d092208",
			3893 => x"09016b04",
			3894 => x"00003d0d",
			3895 => x"01693d0d",
			3896 => x"00003d0d",
			3897 => x"fef43d0d",
			3898 => x"030b2304",
			3899 => x"01803d0d",
			3900 => x"00039e04",
			3901 => x"fe763d0d",
			3902 => x"08036e08",
			3903 => x"0c065204",
			3904 => x"ffce3d0d",
			3905 => x"01873d0d",
			3906 => x"ff2d3d0d",
			3907 => x"09018b04",
			3908 => x"fe733dc9",
			3909 => x"030b132c",
			3910 => x"020a5b08",
			3911 => x"0b075f04",
			3912 => x"fef53dc9",
			3913 => x"00003dc9",
			3914 => x"0101501c",
			3915 => x"0e0a5110",
			3916 => x"01012308",
			3917 => x"0f0a6e04",
			3918 => x"00a13dc9",
			3919 => x"ff383dc9",
			3920 => x"0706eb04",
			3921 => x"01513dc9",
			3922 => x"00003dc9",
			3923 => x"040c2408",
			3924 => x"06018c04",
			3925 => x"00003dc9",
			3926 => x"fe913dc9",
			3927 => x"00313dc9",
			3928 => x"0c063004",
			3929 => x"00003dc9",
			3930 => x"016b3dc9",
			3931 => x"0706f514",
			3932 => x"01015f08",
			3933 => x"09021804",
			3934 => x"00003dc9",
			3935 => x"fe763dc9",
			3936 => x"0e0b5104",
			3937 => x"00ac3dc9",
			3938 => x"08032504",
			3939 => x"00003dc9",
			3940 => x"ff7b3dc9",
			3941 => x"07072814",
			3942 => x"09021d0c",
			3943 => x"0601b008",
			3944 => x"09020a04",
			3945 => x"00003dc9",
			3946 => x"00483dc9",
			3947 => x"ff5f3dc9",
			3948 => x"040b2e04",
			3949 => x"00003dc9",
			3950 => x"01383dc9",
			3951 => x"0c06aa04",
			3952 => x"00003dc9",
			3953 => x"ff273dc9",
			3954 => x"0c061404",
			3955 => x"fe8d3e95",
			3956 => x"0b07b544",
			3957 => x"0c066c28",
			3958 => x"07068310",
			3959 => x"07066e04",
			3960 => x"00003e95",
			3961 => x"0003c804",
			3962 => x"00003e95",
			3963 => x"0f0af304",
			3964 => x"013f3e95",
			3965 => x"00003e95",
			3966 => x"0601a110",
			3967 => x"0b076308",
			3968 => x"020ad904",
			3969 => x"ff2d3e95",
			3970 => x"00003e95",
			3971 => x"01013b04",
			3972 => x"00003e95",
			3973 => x"00e73e95",
			3974 => x"020b0f04",
			3975 => x"00003e95",
			3976 => x"feba3e95",
			3977 => x"01013508",
			3978 => x"0c066e04",
			3979 => x"00003e95",
			3980 => x"ffab3e95",
			3981 => x"0e0b0708",
			3982 => x"0f0b6404",
			3983 => x"01683e95",
			3984 => x"00003e95",
			3985 => x"030b4104",
			3986 => x"ff9e3e95",
			3987 => x"0f0be504",
			3988 => x"00683e95",
			3989 => x"00003e95",
			3990 => x"01016010",
			3991 => x"06018e04",
			3992 => x"00003e95",
			3993 => x"0e0b0e08",
			3994 => x"05090a04",
			3995 => x"fe5e3e95",
			3996 => x"00003e95",
			3997 => x"00003e95",
			3998 => x"0601ca0c",
			3999 => x"07070b08",
			4000 => x"0c068d04",
			4001 => x"fff03e95",
			4002 => x"00003e95",
			4003 => x"01443e95",
			4004 => x"ff573e95",
			4005 => x"09018b04",
			4006 => x"fe723f63",
			4007 => x"0601a54c",
			4008 => x"0003a328",
			4009 => x"06019014",
			4010 => x"0706df0c",
			4011 => x"01015908",
			4012 => x"0b079304",
			4013 => x"ff173f63",
			4014 => x"00003f63",
			4015 => x"00833f63",
			4016 => x"01014704",
			4017 => x"00003f63",
			4018 => x"015e3f63",
			4019 => x"0b07b50c",
			4020 => x"01015004",
			4021 => x"fecf3f63",
			4022 => x"030ac104",
			4023 => x"00003f63",
			4024 => x"00cb3f63",
			4025 => x"0f0b0304",
			4026 => x"00003f63",
			4027 => x"fe3f3f63",
			4028 => x"020b771c",
			4029 => x"0c06130c",
			4030 => x"0e08cb08",
			4031 => x"0308df04",
			4032 => x"00003f63",
			4033 => x"002c3f63",
			4034 => x"ff7c3f63",
			4035 => x"020ac808",
			4036 => x"01014f04",
			4037 => x"ffed3f63",
			4038 => x"00003f63",
			4039 => x"07065a04",
			4040 => x"00003f63",
			4041 => x"016e3f63",
			4042 => x"01016704",
			4043 => x"ffa43f63",
			4044 => x"00003f63",
			4045 => x"01015f0c",
			4046 => x"00044e08",
			4047 => x"07073a04",
			4048 => x"feb53f63",
			4049 => x"00003f63",
			4050 => x"00003f63",
			4051 => x"08035608",
			4052 => x"020b1f04",
			4053 => x"00003f63",
			4054 => x"00fd3f63",
			4055 => x"ff7b3f63",
			4056 => x"00003f65",
			4057 => x"05095e04",
			4058 => x"00003f71",
			4059 => x"febf3f71",
			4060 => x"0c06dc04",
			4061 => x"00003f7d",
			4062 => x"ff9a3f7d",
			4063 => x"040c8504",
			4064 => x"fffa3f91",
			4065 => x"040e2304",
			4066 => x"000c3f91",
			4067 => x"00003f91",
			4068 => x"08034d08",
			4069 => x"0802eb04",
			4070 => x"00003fa5",
			4071 => x"00133fa5",
			4072 => x"00003fa5",
			4073 => x"0509d604",
			4074 => x"00003fb9",
			4075 => x"0d0a5304",
			4076 => x"fb463fb9",
			4077 => x"00003fb9",
			4078 => x"0707640c",
			4079 => x"040c5e04",
			4080 => x"00003fd5",
			4081 => x"040e2304",
			4082 => x"00333fd5",
			4083 => x"00003fd5",
			4084 => x"ff6c3fd5",
			4085 => x"0707640c",
			4086 => x"040c3e04",
			4087 => x"00003ff1",
			4088 => x"040e2304",
			4089 => x"001a3ff1",
			4090 => x"00003ff1",
			4091 => x"ff953ff1",
			4092 => x"040c5e0c",
			4093 => x"040b1404",
			4094 => x"00004015",
			4095 => x"040c5204",
			4096 => x"fff14015",
			4097 => x"00004015",
			4098 => x"040e2304",
			4099 => x"001d4015",
			4100 => x"00004015",
			4101 => x"0101500c",
			4102 => x"0a02d108",
			4103 => x"0a026504",
			4104 => x"00004039",
			4105 => x"ffda4039",
			4106 => x"00004039",
			4107 => x"0a02a104",
			4108 => x"003c4039",
			4109 => x"00004039",
			4110 => x"0c06a10c",
			4111 => x"0c05d804",
			4112 => x"0000405d",
			4113 => x"0b07b504",
			4114 => x"0041405d",
			4115 => x"0000405d",
			4116 => x"0706de04",
			4117 => x"0000405d",
			4118 => x"fff5405d",
			4119 => x"040c5e0c",
			4120 => x"040b3604",
			4121 => x"00004089",
			4122 => x"09024f04",
			4123 => x"ffed4089",
			4124 => x"00004089",
			4125 => x"0901bc04",
			4126 => x"00004089",
			4127 => x"0601cc04",
			4128 => x"004b4089",
			4129 => x"00004089",
			4130 => x"09020a0c",
			4131 => x"07066f08",
			4132 => x"0c05d804",
			4133 => x"000040b5",
			4134 => x"000440b5",
			4135 => x"ffc740b5",
			4136 => x"0c065204",
			4137 => x"000040b5",
			4138 => x"07072804",
			4139 => x"005740b5",
			4140 => x"000040b5",
			4141 => x"0c06a110",
			4142 => x"0c05d804",
			4143 => x"000040d9",
			4144 => x"0d097508",
			4145 => x"0d079604",
			4146 => x"000040d9",
			4147 => x"003d40d9",
			4148 => x"000040d9",
			4149 => x"fff940d9",
			4150 => x"0d0a1110",
			4151 => x"0c05f604",
			4152 => x"000040fd",
			4153 => x"0601ca08",
			4154 => x"06017804",
			4155 => x"000040fd",
			4156 => x"001740fd",
			4157 => x"000040fd",
			4158 => x"ffd340fd",
			4159 => x"0f0b1704",
			4160 => x"00004121",
			4161 => x"0101810c",
			4162 => x"0a026104",
			4163 => x"00004121",
			4164 => x"030cdd04",
			4165 => x"ff854121",
			4166 => x"00004121",
			4167 => x"00004121",
			4168 => x"09020a08",
			4169 => x"0b071e04",
			4170 => x"0000414d",
			4171 => x"ffbd414d",
			4172 => x"0c065204",
			4173 => x"0000414d",
			4174 => x"08036e08",
			4175 => x"00039d04",
			4176 => x"0000414d",
			4177 => x"008e414d",
			4178 => x"0000414d",
			4179 => x"07076414",
			4180 => x"040c4708",
			4181 => x"01016004",
			4182 => x"fff94179",
			4183 => x"00004179",
			4184 => x"0901bc04",
			4185 => x"00004179",
			4186 => x"0601ca04",
			4187 => x"00514179",
			4188 => x"00004179",
			4189 => x"fef44179",
			4190 => x"040c470c",
			4191 => x"040b1404",
			4192 => x"000041ad",
			4193 => x"0f0be504",
			4194 => x"ffe841ad",
			4195 => x"000041ad",
			4196 => x"040e230c",
			4197 => x"020a2d04",
			4198 => x"000041ad",
			4199 => x"020b0f04",
			4200 => x"003841ad",
			4201 => x"000041ad",
			4202 => x"000041ad",
			4203 => x"08035e10",
			4204 => x"040c4704",
			4205 => x"000041e1",
			4206 => x"07065a04",
			4207 => x"000041e1",
			4208 => x"0003f104",
			4209 => x"000041e1",
			4210 => x"002c41e1",
			4211 => x"040df508",
			4212 => x"0a02b904",
			4213 => x"000041e1",
			4214 => x"ff8f41e1",
			4215 => x"000041e1",
			4216 => x"08034d14",
			4217 => x"040b1604",
			4218 => x"00004215",
			4219 => x"0c063204",
			4220 => x"00004215",
			4221 => x"07072808",
			4222 => x"01011504",
			4223 => x"00004215",
			4224 => x"00504215",
			4225 => x"00004215",
			4226 => x"040d0e04",
			4227 => x"ff4e4215",
			4228 => x"00004215",
			4229 => x"0b07b514",
			4230 => x"0b067a04",
			4231 => x"00004241",
			4232 => x"020b770c",
			4233 => x"020a1004",
			4234 => x"00004241",
			4235 => x"030b1b04",
			4236 => x"004f4241",
			4237 => x"00004241",
			4238 => x"00004241",
			4239 => x"00004241",
			4240 => x"0b071e10",
			4241 => x"0c05f604",
			4242 => x"00004285",
			4243 => x"040c6004",
			4244 => x"00004285",
			4245 => x"0803a304",
			4246 => x"01324285",
			4247 => x"00004285",
			4248 => x"08034a0c",
			4249 => x"0c065204",
			4250 => x"00004285",
			4251 => x"0c06aa04",
			4252 => x"00204285",
			4253 => x"00004285",
			4254 => x"0e0c8c04",
			4255 => x"ff854285",
			4256 => x"00004285",
			4257 => x"07072814",
			4258 => x"0901bc04",
			4259 => x"000042c1",
			4260 => x"020a9904",
			4261 => x"000042c1",
			4262 => x"08036b08",
			4263 => x"0c063004",
			4264 => x"000042c1",
			4265 => x"004f42c1",
			4266 => x"000042c1",
			4267 => x"06019204",
			4268 => x"000042c1",
			4269 => x"0b07c304",
			4270 => x"000042c1",
			4271 => x"ff2842c1",
			4272 => x"040c5e14",
			4273 => x"01016010",
			4274 => x"0802d804",
			4275 => x"00004305",
			4276 => x"0508fd08",
			4277 => x"06018a04",
			4278 => x"00004305",
			4279 => x"ff884305",
			4280 => x"00004305",
			4281 => x"00004305",
			4282 => x"08036e0c",
			4283 => x"01010b04",
			4284 => x"00004305",
			4285 => x"0a029e04",
			4286 => x"00004305",
			4287 => x"00684305",
			4288 => x"00004305",
			4289 => x"040c4714",
			4290 => x"0b078210",
			4291 => x"0706e10c",
			4292 => x"01016708",
			4293 => x"0802d504",
			4294 => x"00004349",
			4295 => x"ffc84349",
			4296 => x"00004349",
			4297 => x"00004349",
			4298 => x"00004349",
			4299 => x"08035e0c",
			4300 => x"01010b04",
			4301 => x"00004349",
			4302 => x"08032604",
			4303 => x"00004349",
			4304 => x"00a54349",
			4305 => x"00004349",
			4306 => x"0c06dc1c",
			4307 => x"09021f0c",
			4308 => x"0f0a6e04",
			4309 => x"0000438d",
			4310 => x"06018304",
			4311 => x"0000438d",
			4312 => x"fff1438d",
			4313 => x"06018d04",
			4314 => x"0000438d",
			4315 => x"09027408",
			4316 => x"0c063004",
			4317 => x"0000438d",
			4318 => x"0037438d",
			4319 => x"0000438d",
			4320 => x"0b082804",
			4321 => x"0000438d",
			4322 => x"fe40438d",
			4323 => x"07067114",
			4324 => x"0c05f604",
			4325 => x"000043e1",
			4326 => x"040b8e04",
			4327 => x"000043e1",
			4328 => x"0803a308",
			4329 => x"0f0afc04",
			4330 => x"015e43e1",
			4331 => x"000043e1",
			4332 => x"000043e1",
			4333 => x"08034a0c",
			4334 => x"0c063a04",
			4335 => x"000043e1",
			4336 => x"0c06aa04",
			4337 => x"002043e1",
			4338 => x"000043e1",
			4339 => x"06019904",
			4340 => x"000043e1",
			4341 => x"01017904",
			4342 => x"ff7543e1",
			4343 => x"000043e1",
			4344 => x"06019618",
			4345 => x"020a2d04",
			4346 => x"0000441d",
			4347 => x"0a026404",
			4348 => x"0000441d",
			4349 => x"09016b04",
			4350 => x"0000441d",
			4351 => x"0c06c408",
			4352 => x"0c05d804",
			4353 => x"0000441d",
			4354 => x"0128441d",
			4355 => x"0000441d",
			4356 => x"08035304",
			4357 => x"0000441d",
			4358 => x"ffc1441d",
			4359 => x"0c06de18",
			4360 => x"040b3c04",
			4361 => x"00004459",
			4362 => x"09016b04",
			4363 => x"00004459",
			4364 => x"020b690c",
			4365 => x"040b6304",
			4366 => x"00004459",
			4367 => x"0c05d804",
			4368 => x"00004459",
			4369 => x"005c4459",
			4370 => x"00004459",
			4371 => x"08034a04",
			4372 => x"00004459",
			4373 => x"fea84459",
			4374 => x"020ad614",
			4375 => x"020a2d04",
			4376 => x"000044a5",
			4377 => x"06019d0c",
			4378 => x"0100e504",
			4379 => x"000044a5",
			4380 => x"06017c04",
			4381 => x"000044a5",
			4382 => x"001144a5",
			4383 => x"000044a5",
			4384 => x"01016110",
			4385 => x"00039504",
			4386 => x"000044a5",
			4387 => x"06018a04",
			4388 => x"000044a5",
			4389 => x"0a026104",
			4390 => x"000044a5",
			4391 => x"ffb344a5",
			4392 => x"000044a5",
			4393 => x"0d0a1118",
			4394 => x"0c05f604",
			4395 => x"000044d9",
			4396 => x"0601ca10",
			4397 => x"020a2d04",
			4398 => x"000044d9",
			4399 => x"06017c04",
			4400 => x"000044d9",
			4401 => x"0b07b504",
			4402 => x"002244d9",
			4403 => x"000044d9",
			4404 => x"000044d9",
			4405 => x"ffcf44d9",
			4406 => x"020adf18",
			4407 => x"06017804",
			4408 => x"00004525",
			4409 => x"0f0ae610",
			4410 => x"0601a50c",
			4411 => x"0d079604",
			4412 => x"00004525",
			4413 => x"020a1004",
			4414 => x"00004525",
			4415 => x"00b74525",
			4416 => x"00004525",
			4417 => x"00004525",
			4418 => x"0c06a104",
			4419 => x"00004525",
			4420 => x"040b4604",
			4421 => x"00004525",
			4422 => x"06018d04",
			4423 => x"00004525",
			4424 => x"ffa44525",
			4425 => x"040c601c",
			4426 => x"0b078214",
			4427 => x"0802d804",
			4428 => x"00004579",
			4429 => x"09022b0c",
			4430 => x"0c068708",
			4431 => x"0706eb04",
			4432 => x"ff8b4579",
			4433 => x"00004579",
			4434 => x"00004579",
			4435 => x"00004579",
			4436 => x"0d097504",
			4437 => x"001a4579",
			4438 => x"00004579",
			4439 => x"08035e0c",
			4440 => x"0901a904",
			4441 => x"00004579",
			4442 => x"0c06cb04",
			4443 => x"00fa4579",
			4444 => x"00004579",
			4445 => x"00004579",
			4446 => x"0004a724",
			4447 => x"0601a518",
			4448 => x"0b07b50c",
			4449 => x"0b077104",
			4450 => x"000045d5",
			4451 => x"0601a104",
			4452 => x"008a45d5",
			4453 => x"000045d5",
			4454 => x"06018e04",
			4455 => x"000045d5",
			4456 => x"06019a04",
			4457 => x"ffe345d5",
			4458 => x"000045d5",
			4459 => x"0b082808",
			4460 => x"0b070104",
			4461 => x"000045d5",
			4462 => x"ffda45d5",
			4463 => x"000045d5",
			4464 => x"0004ab08",
			4465 => x"02095704",
			4466 => x"000045d5",
			4467 => x"020945d5",
			4468 => x"000045d5",
			4469 => x"040c4720",
			4470 => x"0b078214",
			4471 => x"0802d804",
			4472 => x"00004631",
			4473 => x"0101590c",
			4474 => x"0706f608",
			4475 => x"0a024f04",
			4476 => x"00004631",
			4477 => x"ffb04631",
			4478 => x"00004631",
			4479 => x"00004631",
			4480 => x"0a029608",
			4481 => x"0a025304",
			4482 => x"00004631",
			4483 => x"00044631",
			4484 => x"00004631",
			4485 => x"08035e0c",
			4486 => x"01010b04",
			4487 => x"00004631",
			4488 => x"08032604",
			4489 => x"00004631",
			4490 => x"00bd4631",
			4491 => x"00004631",
			4492 => x"040c4714",
			4493 => x"00039204",
			4494 => x"00004685",
			4495 => x"09024f0c",
			4496 => x"07073808",
			4497 => x"0a026104",
			4498 => x"00004685",
			4499 => x"ffa34685",
			4500 => x"00004685",
			4501 => x"00004685",
			4502 => x"0a02dd14",
			4503 => x"09016b04",
			4504 => x"00004685",
			4505 => x"0003f104",
			4506 => x"00004685",
			4507 => x"0601c208",
			4508 => x"07061304",
			4509 => x"00004685",
			4510 => x"00584685",
			4511 => x"00004685",
			4512 => x"00004685",
			4513 => x"0d097520",
			4514 => x"0c063008",
			4515 => x"040df504",
			4516 => x"ffef46d1",
			4517 => x"000046d1",
			4518 => x"040b1604",
			4519 => x"000046d1",
			4520 => x"08036b10",
			4521 => x"0e0b070c",
			4522 => x"0c06c208",
			4523 => x"01011504",
			4524 => x"000046d1",
			4525 => x"00d846d1",
			4526 => x"000046d1",
			4527 => x"000046d1",
			4528 => x"000046d1",
			4529 => x"01015f04",
			4530 => x"000046d1",
			4531 => x"ffd346d1",
			4532 => x"0d09751c",
			4533 => x"0901bc04",
			4534 => x"0000471d",
			4535 => x"0601b714",
			4536 => x"020a9904",
			4537 => x"0000471d",
			4538 => x"0c06ac0c",
			4539 => x"020bd708",
			4540 => x"0c063004",
			4541 => x"0000471d",
			4542 => x"0088471d",
			4543 => x"0000471d",
			4544 => x"0000471d",
			4545 => x"0000471d",
			4546 => x"0e0c8c08",
			4547 => x"06018e04",
			4548 => x"0000471d",
			4549 => x"ffeb471d",
			4550 => x"0000471d",
			4551 => x"040d5524",
			4552 => x"08034718",
			4553 => x"0901dd04",
			4554 => x"00004779",
			4555 => x"0b07b510",
			4556 => x"0e0b070c",
			4557 => x"030a3904",
			4558 => x"00004779",
			4559 => x"0b071004",
			4560 => x"00004779",
			4561 => x"00b34779",
			4562 => x"00004779",
			4563 => x"00004779",
			4564 => x"040d1b08",
			4565 => x"030c2504",
			4566 => x"ff7f4779",
			4567 => x"00004779",
			4568 => x"00004779",
			4569 => x"0a02dd08",
			4570 => x"06019404",
			4571 => x"00004779",
			4572 => x"01b64779",
			4573 => x"00004779",
			4574 => x"040c5e1c",
			4575 => x"0802d804",
			4576 => x"000047cd",
			4577 => x"0508fd14",
			4578 => x"09023d10",
			4579 => x"06018a04",
			4580 => x"000047cd",
			4581 => x"0b07c308",
			4582 => x"00037d04",
			4583 => x"000047cd",
			4584 => x"ff7247cd",
			4585 => x"000047cd",
			4586 => x"000047cd",
			4587 => x"000047cd",
			4588 => x"08036e0c",
			4589 => x"0901a904",
			4590 => x"000047cd",
			4591 => x"0a029e04",
			4592 => x"000047cd",
			4593 => x"006f47cd",
			4594 => x"000047cd",
			4595 => x"0c06de24",
			4596 => x"040c5e0c",
			4597 => x"0706df08",
			4598 => x"0b079504",
			4599 => x"ffd14821",
			4600 => x"00004821",
			4601 => x"00004821",
			4602 => x"0a02dd14",
			4603 => x"09016b04",
			4604 => x"00004821",
			4605 => x"020bd70c",
			4606 => x"0d093508",
			4607 => x"07061304",
			4608 => x"00004821",
			4609 => x"005d4821",
			4610 => x"00004821",
			4611 => x"00004821",
			4612 => x"00004821",
			4613 => x"08034a04",
			4614 => x"00004821",
			4615 => x"fe914821",
			4616 => x"0f0a6e18",
			4617 => x"0100e504",
			4618 => x"0000487d",
			4619 => x"020a2d04",
			4620 => x"0000487d",
			4621 => x"06019f0c",
			4622 => x"0c05d804",
			4623 => x"0000487d",
			4624 => x"01015704",
			4625 => x"002a487d",
			4626 => x"0000487d",
			4627 => x"0000487d",
			4628 => x"0802e304",
			4629 => x"0000487d",
			4630 => x"0e0c8c10",
			4631 => x"0a026104",
			4632 => x"0000487d",
			4633 => x"00039204",
			4634 => x"0000487d",
			4635 => x"030cdd04",
			4636 => x"ffb2487d",
			4637 => x"0000487d",
			4638 => x"0000487d",
			4639 => x"020aad18",
			4640 => x"020a2d04",
			4641 => x"000048f1",
			4642 => x"06019610",
			4643 => x"06017c04",
			4644 => x"000048f1",
			4645 => x"0c05d804",
			4646 => x"000048f1",
			4647 => x"00037804",
			4648 => x"000048f1",
			4649 => x"016448f1",
			4650 => x"000048f1",
			4651 => x"08035318",
			4652 => x"0003a20c",
			4653 => x"00039204",
			4654 => x"000048f1",
			4655 => x"00039d04",
			4656 => x"fff448f1",
			4657 => x"000048f1",
			4658 => x"0b071004",
			4659 => x"000048f1",
			4660 => x"0b07f604",
			4661 => x"001848f1",
			4662 => x"000048f1",
			4663 => x"0e0c8c08",
			4664 => x"030cdd04",
			4665 => x"ffc748f1",
			4666 => x"000048f1",
			4667 => x"000048f1",
			4668 => x"040d5528",
			4669 => x"01015918",
			4670 => x"0802d804",
			4671 => x"00004955",
			4672 => x"040d2e10",
			4673 => x"0b07b20c",
			4674 => x"0508de08",
			4675 => x"09022b04",
			4676 => x"ff804955",
			4677 => x"00004955",
			4678 => x"00004955",
			4679 => x"00004955",
			4680 => x"00004955",
			4681 => x"0b07d60c",
			4682 => x"08034d08",
			4683 => x"0b074404",
			4684 => x"00004955",
			4685 => x"00334955",
			4686 => x"00004955",
			4687 => x"00004955",
			4688 => x"0a02dd08",
			4689 => x"0100e504",
			4690 => x"00004955",
			4691 => x"01284955",
			4692 => x"00004955",
			4693 => x"0901fa08",
			4694 => x"0f0b1004",
			4695 => x"ff8949b1",
			4696 => x"000049b1",
			4697 => x"0e0b0718",
			4698 => x"0601bb14",
			4699 => x"0b071004",
			4700 => x"000049b1",
			4701 => x"030b320c",
			4702 => x"0b07b508",
			4703 => x"05082e04",
			4704 => x"000049b1",
			4705 => x"00de49b1",
			4706 => x"000049b1",
			4707 => x"000049b1",
			4708 => x"000049b1",
			4709 => x"09024f0c",
			4710 => x"07073808",
			4711 => x"040c5e04",
			4712 => x"ffb649b1",
			4713 => x"000049b1",
			4714 => x"000049b1",
			4715 => x"000049b1",
			4716 => x"05080f10",
			4717 => x"0c05d804",
			4718 => x"00004a1d",
			4719 => x"040c9304",
			4720 => x"00004a1d",
			4721 => x"0803d004",
			4722 => x"01bc4a1d",
			4723 => x"00004a1d",
			4724 => x"01015918",
			4725 => x"06018a04",
			4726 => x"00004a1d",
			4727 => x"07068804",
			4728 => x"00004a1d",
			4729 => x"09022b0c",
			4730 => x"0508f808",
			4731 => x"0802d804",
			4732 => x"00004a1d",
			4733 => x"ff814a1d",
			4734 => x"00004a1d",
			4735 => x"00004a1d",
			4736 => x"0601ca0c",
			4737 => x"0706a104",
			4738 => x"00004a1d",
			4739 => x"00039a04",
			4740 => x"00004a1d",
			4741 => x"00574a1d",
			4742 => x"00004a1d",
			4743 => x"0004a730",
			4744 => x"0c06a120",
			4745 => x"05086a0c",
			4746 => x"020a9b08",
			4747 => x"00037d04",
			4748 => x"00004a89",
			4749 => x"ffc74a89",
			4750 => x"00004a89",
			4751 => x"0601c010",
			4752 => x"0d095b0c",
			4753 => x"01013b04",
			4754 => x"00004a89",
			4755 => x"030ba604",
			4756 => x"00a04a89",
			4757 => x"00004a89",
			4758 => x"00004a89",
			4759 => x"00004a89",
			4760 => x"020adf04",
			4761 => x"00004a89",
			4762 => x"09024f08",
			4763 => x"06018d04",
			4764 => x"00004a89",
			4765 => x"ffa34a89",
			4766 => x"00004a89",
			4767 => x"0004ab04",
			4768 => x"01394a89",
			4769 => x"00004a89",
			4770 => x"020aad1c",
			4771 => x"020a2d04",
			4772 => x"00004afd",
			4773 => x"06019614",
			4774 => x"06017c04",
			4775 => x"00004afd",
			4776 => x"0c05d804",
			4777 => x"00004afd",
			4778 => x"040a9504",
			4779 => x"00004afd",
			4780 => x"0a024f04",
			4781 => x"00004afd",
			4782 => x"01884afd",
			4783 => x"00004afd",
			4784 => x"0d09270c",
			4785 => x"0901ce04",
			4786 => x"00004afd",
			4787 => x"01012304",
			4788 => x"00004afd",
			4789 => x"00144afd",
			4790 => x"09024f10",
			4791 => x"06019104",
			4792 => x"00004afd",
			4793 => x"0802e304",
			4794 => x"00004afd",
			4795 => x"040b1404",
			4796 => x"00004afd",
			4797 => x"ff934afd",
			4798 => x"00004afd",
			4799 => x"01014924",
			4800 => x"0901fa10",
			4801 => x"01010f04",
			4802 => x"fe5d4b91",
			4803 => x"020acb04",
			4804 => x"fe614b91",
			4805 => x"0e09fd04",
			4806 => x"01e14b91",
			4807 => x"fe644b91",
			4808 => x"07068604",
			4809 => x"fe5f4b91",
			4810 => x"0e0a8608",
			4811 => x"01014504",
			4812 => x"03044b91",
			4813 => x"01474b91",
			4814 => x"0c066c04",
			4815 => x"fe534b91",
			4816 => x"00004b91",
			4817 => x"0d08b30c",
			4818 => x"0e0a2a08",
			4819 => x"07066c04",
			4820 => x"ff1a4b91",
			4821 => x"009f4b91",
			4822 => x"fe664b91",
			4823 => x"0a02b414",
			4824 => x"0706a104",
			4825 => x"00684b91",
			4826 => x"0c06cb0c",
			4827 => x"0b07d608",
			4828 => x"09021204",
			4829 => x"01774b91",
			4830 => x"01e34b91",
			4831 => x"00f74b91",
			4832 => x"005f4b91",
			4833 => x"05091704",
			4834 => x"fe994b91",
			4835 => x"009a4b91",
			4836 => x"09020a20",
			4837 => x"09020214",
			4838 => x"0901b204",
			4839 => x"fe5b4c15",
			4840 => x"07065a04",
			4841 => x"fe5f4c15",
			4842 => x"0e0a7008",
			4843 => x"020acb04",
			4844 => x"fe6c4c15",
			4845 => x"02734c15",
			4846 => x"fe654c15",
			4847 => x"05084d04",
			4848 => x"fe5f4c15",
			4849 => x"030aa904",
			4850 => x"028d4c15",
			4851 => x"ff8e4c15",
			4852 => x"0b072004",
			4853 => x"fe624c15",
			4854 => x"08034c18",
			4855 => x"0706a108",
			4856 => x"05084d04",
			4857 => x"fe9d4c15",
			4858 => x"00f04c15",
			4859 => x"0c06cb0c",
			4860 => x"0b07d608",
			4861 => x"09021204",
			4862 => x"01874c15",
			4863 => x"01f84c15",
			4864 => x"011b4c15",
			4865 => x"007b4c15",
			4866 => x"040d2e04",
			4867 => x"fe9d4c15",
			4868 => x"00ca4c15",
			4869 => x"0101472c",
			4870 => x"0902021c",
			4871 => x"0100f804",
			4872 => x"fe594ca1",
			4873 => x"040cb610",
			4874 => x"040c2404",
			4875 => x"fe5b4ca1",
			4876 => x"040c2c04",
			4877 => x"01914ca1",
			4878 => x"0b073304",
			4879 => x"00004ca1",
			4880 => x"fe6f4ca1",
			4881 => x"0c066604",
			4882 => x"03384ca1",
			4883 => x"fe7d4ca1",
			4884 => x"0706a108",
			4885 => x"0c063204",
			4886 => x"fe644ca1",
			4887 => x"00344ca1",
			4888 => x"0e0aaa04",
			4889 => x"02db4ca1",
			4890 => x"00324ca1",
			4891 => x"0d08b304",
			4892 => x"fe554ca1",
			4893 => x"0601cc14",
			4894 => x"0c063a04",
			4895 => x"00b94ca1",
			4896 => x"0601c20c",
			4897 => x"040ca008",
			4898 => x"0601a904",
			4899 => x"02134ca1",
			4900 => x"01814ca1",
			4901 => x"03274ca1",
			4902 => x"00994ca1",
			4903 => x"fe7e4ca1",
			4904 => x"01014930",
			4905 => x"09020e28",
			4906 => x"0902021c",
			4907 => x"06018a04",
			4908 => x"db884d3d",
			4909 => x"0f0ac310",
			4910 => x"020acb08",
			4911 => x"07067004",
			4912 => x"dba74d3d",
			4913 => x"dcfd4d3d",
			4914 => x"01010f04",
			4915 => x"dbc44d3d",
			4916 => x"e5fc4d3d",
			4917 => x"06019404",
			4918 => x"dc924d3d",
			4919 => x"db8a4d3d",
			4920 => x"0c065008",
			4921 => x"05082e04",
			4922 => x"db8c4d3d",
			4923 => x"dd854d3d",
			4924 => x"e3a94d3d",
			4925 => x"06018d04",
			4926 => x"ea7f4d3d",
			4927 => x"dba64d3d",
			4928 => x"05086a08",
			4929 => x"0706a104",
			4930 => x"db8d4d3d",
			4931 => x"e3b44d3d",
			4932 => x"08035610",
			4933 => x"0706b408",
			4934 => x"0a027504",
			4935 => x"eaa04d3d",
			4936 => x"e47b4d3d",
			4937 => x"0c06dc04",
			4938 => x"eb414d3d",
			4939 => x"e77d4d3d",
			4940 => x"0601ca04",
			4941 => x"df964d3d",
			4942 => x"dbb64d3d",
			4943 => x"0c063a08",
			4944 => x"0a02cb04",
			4945 => x"ff764dc1",
			4946 => x"00004dc1",
			4947 => x"0d094e20",
			4948 => x"01015018",
			4949 => x"0d090110",
			4950 => x"0d088204",
			4951 => x"00004dc1",
			4952 => x"00046b08",
			4953 => x"00035b04",
			4954 => x"00004dc1",
			4955 => x"00344dc1",
			4956 => x"00004dc1",
			4957 => x"00039504",
			4958 => x"00004dc1",
			4959 => x"ffe34dc1",
			4960 => x"0b075f04",
			4961 => x"00004dc1",
			4962 => x"00af4dc1",
			4963 => x"09022a08",
			4964 => x"0c06ac04",
			4965 => x"00124dc1",
			4966 => x"00004dc1",
			4967 => x"0c06a410",
			4968 => x"0508fd0c",
			4969 => x"030b1b04",
			4970 => x"00004dc1",
			4971 => x"01018104",
			4972 => x"ff504dc1",
			4973 => x"00004dc1",
			4974 => x"00004dc1",
			4975 => x"00004dc1",
			4976 => x"0c061304",
			4977 => x"fec44e35",
			4978 => x"06018e0c",
			4979 => x"0f0a8a04",
			4980 => x"00004e35",
			4981 => x"01013f04",
			4982 => x"00004e35",
			4983 => x"00d14e35",
			4984 => x"00039a10",
			4985 => x"0f0aed04",
			4986 => x"00004e35",
			4987 => x"0c06a408",
			4988 => x"00039204",
			4989 => x"00004e35",
			4990 => x"ff1c4e35",
			4991 => x"00004e35",
			4992 => x"0601a910",
			4993 => x"040b3c04",
			4994 => x"00004e35",
			4995 => x"01010b04",
			4996 => x"00004e35",
			4997 => x"0e0b5104",
			4998 => x"00f14e35",
			4999 => x"00004e35",
			5000 => x"01015b04",
			5001 => x"ff4d4e35",
			5002 => x"0601ca04",
			5003 => x"004d4e35",
			5004 => x"ff964e35",
			5005 => x"01014734",
			5006 => x"09020224",
			5007 => x"0100f804",
			5008 => x"fe574ec9",
			5009 => x"040cb610",
			5010 => x"040c2404",
			5011 => x"fe594ec9",
			5012 => x"040c2c04",
			5013 => x"01bb4ec9",
			5014 => x"0b073304",
			5015 => x"00004ec9",
			5016 => x"fe694ec9",
			5017 => x"020b5304",
			5018 => x"04d34ec9",
			5019 => x"040ceb08",
			5020 => x"05090a04",
			5021 => x"01484ec9",
			5022 => x"ff8f4ec9",
			5023 => x"fe764ec9",
			5024 => x"0706a108",
			5025 => x"0c063204",
			5026 => x"fe604ec9",
			5027 => x"00264ec9",
			5028 => x"0e0aaa04",
			5029 => x"032a4ec9",
			5030 => x"002e4ec9",
			5031 => x"0d08b304",
			5032 => x"fe514ec9",
			5033 => x"08037310",
			5034 => x"0c063a04",
			5035 => x"00df4ec9",
			5036 => x"08035208",
			5037 => x"0c06de04",
			5038 => x"02354ec9",
			5039 => x"01744ec9",
			5040 => x"01454ec9",
			5041 => x"fe904ec9",
			5042 => x"01014924",
			5043 => x"0100f804",
			5044 => x"fe604f75",
			5045 => x"040c6014",
			5046 => x"0706b708",
			5047 => x"05088604",
			5048 => x"fe5a4f75",
			5049 => x"ffd34f75",
			5050 => x"06019408",
			5051 => x"01013b04",
			5052 => x"fed14f75",
			5053 => x"01eb4f75",
			5054 => x"fe654f75",
			5055 => x"020b4904",
			5056 => x"03824f75",
			5057 => x"0601a904",
			5058 => x"01704f75",
			5059 => x"fe614f75",
			5060 => x"0c063a0c",
			5061 => x"0a027a08",
			5062 => x"040b2e04",
			5063 => x"fe084f75",
			5064 => x"013a4f75",
			5065 => x"fe284f75",
			5066 => x"0601c220",
			5067 => x"0b07630c",
			5068 => x"0e0a9404",
			5069 => x"02084f75",
			5070 => x"09022e04",
			5071 => x"fe4f4f75",
			5072 => x"01a64f75",
			5073 => x"0601ad0c",
			5074 => x"0b07b804",
			5075 => x"01ca4f75",
			5076 => x"0b07c304",
			5077 => x"01234f75",
			5078 => x"01b34f75",
			5079 => x"01016c04",
			5080 => x"ff364f75",
			5081 => x"01e94f75",
			5082 => x"040d5504",
			5083 => x"fee54f75",
			5084 => x"00374f75",
			5085 => x"01012304",
			5086 => x"feee4ff1",
			5087 => x"040b6324",
			5088 => x"0b078210",
			5089 => x"0802d804",
			5090 => x"00004ff1",
			5091 => x"01015908",
			5092 => x"0c068704",
			5093 => x"fef24ff1",
			5094 => x"00004ff1",
			5095 => x"00004ff1",
			5096 => x"030b2a0c",
			5097 => x"0b07c508",
			5098 => x"0a027404",
			5099 => x"00b74ff1",
			5100 => x"00004ff1",
			5101 => x"00004ff1",
			5102 => x"0a026404",
			5103 => x"ffb94ff1",
			5104 => x"00004ff1",
			5105 => x"0601c214",
			5106 => x"0c06dc10",
			5107 => x"0c063004",
			5108 => x"00004ff1",
			5109 => x"0e0b5108",
			5110 => x"01014104",
			5111 => x"00004ff1",
			5112 => x"00f14ff1",
			5113 => x"00004ff1",
			5114 => x"00004ff1",
			5115 => x"ffc84ff1",
			5116 => x"020a5b08",
			5117 => x"0b075f04",
			5118 => x"fe9a508d",
			5119 => x"0000508d",
			5120 => x"0601a52c",
			5121 => x"0d095b1c",
			5122 => x"01015518",
			5123 => x"0e0aa20c",
			5124 => x"09018b04",
			5125 => x"0000508d",
			5126 => x"040b8e04",
			5127 => x"0000508d",
			5128 => x"00e0508d",
			5129 => x"0706e208",
			5130 => x"0003f304",
			5131 => x"ff09508d",
			5132 => x"0000508d",
			5133 => x"0000508d",
			5134 => x"0142508d",
			5135 => x"09022e08",
			5136 => x"01014904",
			5137 => x"0000508d",
			5138 => x"007c508d",
			5139 => x"0003a204",
			5140 => x"feea508d",
			5141 => x"0000508d",
			5142 => x"09024f0c",
			5143 => x"040cce08",
			5144 => x"0a028b04",
			5145 => x"0000508d",
			5146 => x"fee1508d",
			5147 => x"0000508d",
			5148 => x"09026b08",
			5149 => x"01017404",
			5150 => x"0000508d",
			5151 => x"00a0508d",
			5152 => x"0a02cb04",
			5153 => x"0000508d",
			5154 => x"ffe6508d",
			5155 => x"0100f804",
			5156 => x"fec95109",
			5157 => x"0601a12c",
			5158 => x"09022a18",
			5159 => x"09021210",
			5160 => x"0003f30c",
			5161 => x"06018504",
			5162 => x"00005109",
			5163 => x"01014d04",
			5164 => x"ff8b5109",
			5165 => x"00005109",
			5166 => x"00b15109",
			5167 => x"0d08b304",
			5168 => x"00005109",
			5169 => x"01165109",
			5170 => x"0a026710",
			5171 => x"0e0ac404",
			5172 => x"00005109",
			5173 => x"0c068f08",
			5174 => x"0d094904",
			5175 => x"00005109",
			5176 => x"fee35109",
			5177 => x"00005109",
			5178 => x"00ae5109",
			5179 => x"07068804",
			5180 => x"00005109",
			5181 => x"01015f04",
			5182 => x"ff285109",
			5183 => x"08036804",
			5184 => x"00505109",
			5185 => x"ffb65109",
			5186 => x"020a5b0c",
			5187 => x"0802d804",
			5188 => x"0000519d",
			5189 => x"0f0a6e04",
			5190 => x"ff52519d",
			5191 => x"0000519d",
			5192 => x"0508dc18",
			5193 => x"0601b214",
			5194 => x"09018b04",
			5195 => x"0000519d",
			5196 => x"0f0bae0c",
			5197 => x"040b1604",
			5198 => x"0000519d",
			5199 => x"06018504",
			5200 => x"0000519d",
			5201 => x"00b5519d",
			5202 => x"0000519d",
			5203 => x"0000519d",
			5204 => x"07070c14",
			5205 => x"09022a04",
			5206 => x"0000519d",
			5207 => x"030b1b04",
			5208 => x"0000519d",
			5209 => x"0b07c308",
			5210 => x"0d094e04",
			5211 => x"0000519d",
			5212 => x"ff49519d",
			5213 => x"0000519d",
			5214 => x"0601ca10",
			5215 => x"0f0b0904",
			5216 => x"0000519d",
			5217 => x"0e0ab804",
			5218 => x"0000519d",
			5219 => x"09020a04",
			5220 => x"0000519d",
			5221 => x"00d0519d",
			5222 => x"ffe2519d",
			5223 => x"0901ce08",
			5224 => x"040dca04",
			5225 => x"fea25221",
			5226 => x"00005221",
			5227 => x"0706a108",
			5228 => x"00040c04",
			5229 => x"ff435221",
			5230 => x"00005221",
			5231 => x"0b07b518",
			5232 => x"0c06ac10",
			5233 => x"0e0b940c",
			5234 => x"00038104",
			5235 => x"00005221",
			5236 => x"0901df04",
			5237 => x"00005221",
			5238 => x"011e5221",
			5239 => x"00005221",
			5240 => x"09021f04",
			5241 => x"fffd5221",
			5242 => x"00005221",
			5243 => x"0e0ac908",
			5244 => x"040b3604",
			5245 => x"00005221",
			5246 => x"ff475221",
			5247 => x"0601cc10",
			5248 => x"07070c08",
			5249 => x"0706fb04",
			5250 => x"00005221",
			5251 => x"ffdc5221",
			5252 => x"01014b04",
			5253 => x"00005221",
			5254 => x"010f5221",
			5255 => x"ffa05221",
			5256 => x"0c061304",
			5257 => x"ff53529d",
			5258 => x"0601ba30",
			5259 => x"040b631c",
			5260 => x"0b078210",
			5261 => x"06018904",
			5262 => x"0000529d",
			5263 => x"01015908",
			5264 => x"0c068804",
			5265 => x"ff2d529d",
			5266 => x"0000529d",
			5267 => x"0000529d",
			5268 => x"0b07b508",
			5269 => x"01014704",
			5270 => x"0000529d",
			5271 => x"0073529d",
			5272 => x"0000529d",
			5273 => x"0e0b9410",
			5274 => x"0901a904",
			5275 => x"0000529d",
			5276 => x"07065a04",
			5277 => x"0000529d",
			5278 => x"01010b04",
			5279 => x"0000529d",
			5280 => x"00b3529d",
			5281 => x"0000529d",
			5282 => x"01017904",
			5283 => x"ff74529d",
			5284 => x"08036e04",
			5285 => x"0017529d",
			5286 => x"0000529d",
			5287 => x"0c061304",
			5288 => x"febc5321",
			5289 => x"06018e10",
			5290 => x"030a3904",
			5291 => x"00005321",
			5292 => x"01013f04",
			5293 => x"00005321",
			5294 => x"0f0a8a04",
			5295 => x"00005321",
			5296 => x"00e25321",
			5297 => x"00039a10",
			5298 => x"0f0aed04",
			5299 => x"00005321",
			5300 => x"0c06a408",
			5301 => x"0802e304",
			5302 => x"00005321",
			5303 => x"ff035321",
			5304 => x"00005321",
			5305 => x"0601a910",
			5306 => x"0a026404",
			5307 => x"00005321",
			5308 => x"01010b04",
			5309 => x"00005321",
			5310 => x"0f0b9804",
			5311 => x"00f65321",
			5312 => x"00005321",
			5313 => x"01015b04",
			5314 => x"ff415321",
			5315 => x"0601ca08",
			5316 => x"00042904",
			5317 => x"00785321",
			5318 => x"00005321",
			5319 => x"ff8c5321",
			5320 => x"09018b04",
			5321 => x"fe9153b5",
			5322 => x"0601a530",
			5323 => x"0003a320",
			5324 => x"030b2a18",
			5325 => x"0706c90c",
			5326 => x"040b1608",
			5327 => x"0b077104",
			5328 => x"feeb53b5",
			5329 => x"000053b5",
			5330 => x"000053b5",
			5331 => x"07072508",
			5332 => x"01014304",
			5333 => x"000053b5",
			5334 => x"013353b5",
			5335 => x"000053b5",
			5336 => x"09022e04",
			5337 => x"000053b5",
			5338 => x"fea953b5",
			5339 => x"040b4a04",
			5340 => x"000053b5",
			5341 => x"0f0bc908",
			5342 => x"0f09e104",
			5343 => x"000053b5",
			5344 => x"010353b5",
			5345 => x"000053b5",
			5346 => x"09024f0c",
			5347 => x"040cce08",
			5348 => x"08031204",
			5349 => x"000053b5",
			5350 => x"fed653b5",
			5351 => x"000053b5",
			5352 => x"08036e08",
			5353 => x"0c067004",
			5354 => x"000053b5",
			5355 => x"00e553b5",
			5356 => x"fff253b5",
			5357 => x"01013f28",
			5358 => x"06018a04",
			5359 => x"fe665491",
			5360 => x"0f0aa610",
			5361 => x"040d2e08",
			5362 => x"030a1204",
			5363 => x"febe5491",
			5364 => x"00005491",
			5365 => x"09016704",
			5366 => x"ff915491",
			5367 => x"01f45491",
			5368 => x"06019408",
			5369 => x"06018e04",
			5370 => x"ff7b5491",
			5371 => x"008c5491",
			5372 => x"030a4908",
			5373 => x"030a3904",
			5374 => x"ff9c5491",
			5375 => x"00005491",
			5376 => x"fe885491",
			5377 => x"01015024",
			5378 => x"06018c10",
			5379 => x"030a3904",
			5380 => x"fed15491",
			5381 => x"0f0a8a08",
			5382 => x"020a6b04",
			5383 => x"01415491",
			5384 => x"ffb25491",
			5385 => x"01f55491",
			5386 => x"040c2c10",
			5387 => x"0e0a5108",
			5388 => x"0d088d04",
			5389 => x"fffa5491",
			5390 => x"00c75491",
			5391 => x"040b0204",
			5392 => x"00005491",
			5393 => x"fde15491",
			5394 => x"00ea5491",
			5395 => x"08034d1c",
			5396 => x"0d097514",
			5397 => x"05084d04",
			5398 => x"ff655491",
			5399 => x"0c06ac08",
			5400 => x"0e0b9404",
			5401 => x"019c5491",
			5402 => x"00005491",
			5403 => x"0d095004",
			5404 => x"01595491",
			5405 => x"00005491",
			5406 => x"0802ee04",
			5407 => x"fe975491",
			5408 => x"01895491",
			5409 => x"020bf304",
			5410 => x"00005491",
			5411 => x"fee15491",
			5412 => x"0c06140c",
			5413 => x"020a9b04",
			5414 => x"fe6a554d",
			5415 => x"020aa104",
			5416 => x"0091554d",
			5417 => x"fec1554d",
			5418 => x"01015c40",
			5419 => x"030b1324",
			5420 => x"0901bc0c",
			5421 => x"0c061708",
			5422 => x"0100fa04",
			5423 => x"0000554d",
			5424 => x"0050554d",
			5425 => x"fecc554d",
			5426 => x"06018c08",
			5427 => x"0f0a4204",
			5428 => x"0000554d",
			5429 => x"018f554d",
			5430 => x"040bc408",
			5431 => x"01014f04",
			5432 => x"feb5554d",
			5433 => x"0076554d",
			5434 => x"0601b204",
			5435 => x"0154554d",
			5436 => x"0000554d",
			5437 => x"0706f510",
			5438 => x"09021808",
			5439 => x"06019f04",
			5440 => x"001e554d",
			5441 => x"0000554d",
			5442 => x"09022a04",
			5443 => x"feb5554d",
			5444 => x"fccd554d",
			5445 => x"0a028704",
			5446 => x"014e554d",
			5447 => x"0d091b04",
			5448 => x"0000554d",
			5449 => x"fec0554d",
			5450 => x"0a026408",
			5451 => x"09023704",
			5452 => x"0138554d",
			5453 => x"feb4554d",
			5454 => x"0601c208",
			5455 => x"0d090104",
			5456 => x"0000554d",
			5457 => x"018f554d",
			5458 => x"002f554d",
			5459 => x"0c061304",
			5460 => x"fecd55f1",
			5461 => x"030b5334",
			5462 => x"040b3c1c",
			5463 => x"0601910c",
			5464 => x"09020a04",
			5465 => x"000055f1",
			5466 => x"0706a104",
			5467 => x"000055f1",
			5468 => x"00af55f1",
			5469 => x"0c068d0c",
			5470 => x"0f0aed04",
			5471 => x"000055f1",
			5472 => x"0802ed04",
			5473 => x"ff1e55f1",
			5474 => x"000055f1",
			5475 => x"000055f1",
			5476 => x"0901ce08",
			5477 => x"0f0a6e04",
			5478 => x"000055f1",
			5479 => x"ffcf55f1",
			5480 => x"0601bb0c",
			5481 => x"0c06c208",
			5482 => x"0c063004",
			5483 => x"000055f1",
			5484 => x"010855f1",
			5485 => x"000055f1",
			5486 => x"000055f1",
			5487 => x"0c06a410",
			5488 => x"0a027004",
			5489 => x"000055f1",
			5490 => x"0f0b4a04",
			5491 => x"000055f1",
			5492 => x"0e0b0704",
			5493 => x"000055f1",
			5494 => x"ff4655f1",
			5495 => x"0601ca08",
			5496 => x"01014b04",
			5497 => x"000055f1",
			5498 => x"00be55f1",
			5499 => x"ffd355f1",
			5500 => x"09020520",
			5501 => x"020a2d04",
			5502 => x"fe6356b5",
			5503 => x"0e0a7018",
			5504 => x"0c05f604",
			5505 => x"fe8156b5",
			5506 => x"040c2408",
			5507 => x"01014104",
			5508 => x"fe9656b5",
			5509 => x"000056b5",
			5510 => x"0c061a04",
			5511 => x"02e656b5",
			5512 => x"0901dd04",
			5513 => x"fe7356b5",
			5514 => x"010e56b5",
			5515 => x"fe6856b5",
			5516 => x"0b07631c",
			5517 => x"040b6310",
			5518 => x"06018908",
			5519 => x"05084d04",
			5520 => x"fec156b5",
			5521 => x"018656b5",
			5522 => x"01015704",
			5523 => x"fe0b56b5",
			5524 => x"ffa356b5",
			5525 => x"0e0a9a04",
			5526 => x"02f756b5",
			5527 => x"05088604",
			5528 => x"fea256b5",
			5529 => x"009b56b5",
			5530 => x"0c06dc24",
			5531 => x"0601bb18",
			5532 => x"0d097510",
			5533 => x"0c06ac08",
			5534 => x"0508fb04",
			5535 => x"01ab56b5",
			5536 => x"010656b5",
			5537 => x"0508cf04",
			5538 => x"000056b5",
			5539 => x"019856b5",
			5540 => x"020b2404",
			5541 => x"feeb56b5",
			5542 => x"019256b5",
			5543 => x"01017904",
			5544 => x"fef156b5",
			5545 => x"0c068b04",
			5546 => x"ffef56b5",
			5547 => x"019156b5",
			5548 => x"ff3b56b5",
			5549 => x"09020828",
			5550 => x"020a2d04",
			5551 => x"fe625771",
			5552 => x"0601a520",
			5553 => x"040c240c",
			5554 => x"0c066604",
			5555 => x"fe635771",
			5556 => x"0706c904",
			5557 => x"00a35771",
			5558 => x"ff035771",
			5559 => x"09016b04",
			5560 => x"fe9c5771",
			5561 => x"020b3208",
			5562 => x"07061304",
			5563 => x"ff9b5771",
			5564 => x"03035771",
			5565 => x"0901cc04",
			5566 => x"fe875771",
			5567 => x"01c85771",
			5568 => x"fe655771",
			5569 => x"0c063a08",
			5570 => x"05086a04",
			5571 => x"fe455771",
			5572 => x"00a95771",
			5573 => x"0a02961c",
			5574 => x"0d097514",
			5575 => x"0b076308",
			5576 => x"0e0a9404",
			5577 => x"017b5771",
			5578 => x"ffe75771",
			5579 => x"0d094e04",
			5580 => x"01ac5771",
			5581 => x"0b079304",
			5582 => x"ff2c5771",
			5583 => x"016f5771",
			5584 => x"0003a704",
			5585 => x"fe755771",
			5586 => x"01965771",
			5587 => x"040c5e08",
			5588 => x"09024104",
			5589 => x"fdaf5771",
			5590 => x"012c5771",
			5591 => x"0601ca08",
			5592 => x"0e0bab04",
			5593 => x"01eb5771",
			5594 => x"00f35771",
			5595 => x"fedc5771",
			5596 => x"020a2d08",
			5597 => x"030a3904",
			5598 => x"fe6c581d",
			5599 => x"0000581d",
			5600 => x"0f0adf20",
			5601 => x"0601a714",
			5602 => x"0c05d804",
			5603 => x"ffd6581d",
			5604 => x"09016b04",
			5605 => x"0000581d",
			5606 => x"040a9504",
			5607 => x"0000581d",
			5608 => x"06017d04",
			5609 => x"0000581d",
			5610 => x"015b581d",
			5611 => x"0f0aad08",
			5612 => x"01013004",
			5613 => x"0000581d",
			5614 => x"0068581d",
			5615 => x"ff52581d",
			5616 => x"01016128",
			5617 => x"0b07b51c",
			5618 => x"0e0b0710",
			5619 => x"09021f08",
			5620 => x"020af104",
			5621 => x"feb5581d",
			5622 => x"001f581d",
			5623 => x"05084d04",
			5624 => x"0000581d",
			5625 => x"0160581d",
			5626 => x"0d095008",
			5627 => x"0c06a504",
			5628 => x"fe69581d",
			5629 => x"0000581d",
			5630 => x"0000581d",
			5631 => x"09022e08",
			5632 => x"040bbd04",
			5633 => x"00db581d",
			5634 => x"fee9581d",
			5635 => x"fd97581d",
			5636 => x"08036504",
			5637 => x"0176581d",
			5638 => x"0000581d",
			5639 => x"09020224",
			5640 => x"06018a04",
			5641 => x"fe645911",
			5642 => x"0601960c",
			5643 => x"040c2404",
			5644 => x"fec15911",
			5645 => x"09016b04",
			5646 => x"ff5e5911",
			5647 => x"02245911",
			5648 => x"0901ce04",
			5649 => x"fe625911",
			5650 => x"040ce10c",
			5651 => x"0901df08",
			5652 => x"0901dd04",
			5653 => x"ffdf5911",
			5654 => x"00005911",
			5655 => x"fe7b5911",
			5656 => x"01135911",
			5657 => x"0b077128",
			5658 => x"0e0aa214",
			5659 => x"040b8a10",
			5660 => x"05086a08",
			5661 => x"0802d404",
			5662 => x"002b5911",
			5663 => x"fe525911",
			5664 => x"06019104",
			5665 => x"016c5911",
			5666 => x"00005911",
			5667 => x"02845911",
			5668 => x"0c066d10",
			5669 => x"040b5604",
			5670 => x"fc7a5911",
			5671 => x"0a028804",
			5672 => x"00675911",
			5673 => x"00041804",
			5674 => x"fe4b5911",
			5675 => x"00005911",
			5676 => x"017c5911",
			5677 => x"0d094e10",
			5678 => x"0c06c208",
			5679 => x"0e0b6304",
			5680 => x"019e5911",
			5681 => x"00005911",
			5682 => x"0b07b104",
			5683 => x"00e65911",
			5684 => x"ff935911",
			5685 => x"020af410",
			5686 => x"030b1b08",
			5687 => x"040b3c04",
			5688 => x"01835911",
			5689 => x"00005911",
			5690 => x"0a026704",
			5691 => x"fbe85911",
			5692 => x"01245911",
			5693 => x"08035208",
			5694 => x"0e0ad704",
			5695 => x"00005911",
			5696 => x"01a35911",
			5697 => x"040d5504",
			5698 => x"fe995911",
			5699 => x"00a35911",
			5700 => x"0c061304",
			5701 => x"fe7f59bd",
			5702 => x"0b07b538",
			5703 => x"09021f24",
			5704 => x"0e0aa214",
			5705 => x"0901a904",
			5706 => x"ff8d59bd",
			5707 => x"040b7608",
			5708 => x"0706a104",
			5709 => x"ff4259bd",
			5710 => x"007259bd",
			5711 => x"0601a904",
			5712 => x"014659bd",
			5713 => x"000059bd",
			5714 => x"06018d04",
			5715 => x"000059bd",
			5716 => x"01015408",
			5717 => x"0508f804",
			5718 => x"febf59bd",
			5719 => x"000059bd",
			5720 => x"000059bd",
			5721 => x"0c06520c",
			5722 => x"0c063404",
			5723 => x"002559bd",
			5724 => x"0706c904",
			5725 => x"ff5859bd",
			5726 => x"000059bd",
			5727 => x"09026404",
			5728 => x"015459bd",
			5729 => x"000059bd",
			5730 => x"01016010",
			5731 => x"09022e0c",
			5732 => x"0601a908",
			5733 => x"01014904",
			5734 => x"000059bd",
			5735 => x"008d59bd",
			5736 => x"ff4559bd",
			5737 => x"fea959bd",
			5738 => x"08036808",
			5739 => x"0b07b804",
			5740 => x"000059bd",
			5741 => x"00df59bd",
			5742 => x"fffc59bd",
			5743 => x"0901dd08",
			5744 => x"040da904",
			5745 => x"fe9b5a69",
			5746 => x"00005a69",
			5747 => x"06018a0c",
			5748 => x"07069b08",
			5749 => x"040b4a04",
			5750 => x"ffd15a69",
			5751 => x"00005a69",
			5752 => x"00ed5a69",
			5753 => x"0003a318",
			5754 => x"0f0b030c",
			5755 => x"0b077108",
			5756 => x"0706b704",
			5757 => x"00005a69",
			5758 => x"ff595a69",
			5759 => x"00a35a69",
			5760 => x"09022a04",
			5761 => x"00005a69",
			5762 => x"0d094e04",
			5763 => x"00005a69",
			5764 => x"feb15a69",
			5765 => x"0601a510",
			5766 => x"020ad604",
			5767 => x"00005a69",
			5768 => x"07068604",
			5769 => x"00005a69",
			5770 => x"07073c04",
			5771 => x"01145a69",
			5772 => x"00005a69",
			5773 => x"040c5e0c",
			5774 => x"09024f08",
			5775 => x"0a028b04",
			5776 => x"00005a69",
			5777 => x"ff145a69",
			5778 => x"00005a69",
			5779 => x"00042908",
			5780 => x"09020204",
			5781 => x"00005a69",
			5782 => x"009b5a69",
			5783 => x"040d4204",
			5784 => x"ff3d5a69",
			5785 => x"00125a69",
			5786 => x"0c061304",
			5787 => x"fe7a5b1d",
			5788 => x"0b07b538",
			5789 => x"020b7728",
			5790 => x"040b1614",
			5791 => x"0706c90c",
			5792 => x"06017d04",
			5793 => x"00005b1d",
			5794 => x"0b077104",
			5795 => x"fe8e5b1d",
			5796 => x"00005b1d",
			5797 => x"01014304",
			5798 => x"00005b1d",
			5799 => x"01095b1d",
			5800 => x"0c06ac0c",
			5801 => x"0901a904",
			5802 => x"fffc5b1d",
			5803 => x"07066e04",
			5804 => x"00005b1d",
			5805 => x"011b5b1d",
			5806 => x"0508cf04",
			5807 => x"ff765b1d",
			5808 => x"00005b1d",
			5809 => x"09023f08",
			5810 => x"0c06aa04",
			5811 => x"fef75b1d",
			5812 => x"00005b1d",
			5813 => x"0a02a604",
			5814 => x"00005b1d",
			5815 => x"00005b1d",
			5816 => x"01016014",
			5817 => x"06018e04",
			5818 => x"00005b1d",
			5819 => x"0c068904",
			5820 => x"00005b1d",
			5821 => x"0e0b0e08",
			5822 => x"0508dc04",
			5823 => x"00005b1d",
			5824 => x"fe815b1d",
			5825 => x"00005b1d",
			5826 => x"0a02cb08",
			5827 => x"0b07b804",
			5828 => x"00005b1d",
			5829 => x"00ea5b1d",
			5830 => x"ffec5b1d",
			5831 => x"020a2d08",
			5832 => x"0b074404",
			5833 => x"fe6b5be9",
			5834 => x"00005be9",
			5835 => x"09021f3c",
			5836 => x"0e0aa21c",
			5837 => x"09020e14",
			5838 => x"040c6008",
			5839 => x"06018504",
			5840 => x"00005be9",
			5841 => x"fe9d5be9",
			5842 => x"0a02dd08",
			5843 => x"0c065004",
			5844 => x"015a5be9",
			5845 => x"00005be9",
			5846 => x"ff835be9",
			5847 => x"0d08b304",
			5848 => x"00005be9",
			5849 => x"014a5be9",
			5850 => x"0c066d10",
			5851 => x"040c440c",
			5852 => x"0b078b08",
			5853 => x"0f0aed04",
			5854 => x"00005be9",
			5855 => x"fe0b5be9",
			5856 => x"00005be9",
			5857 => x"00005be9",
			5858 => x"0c06ac0c",
			5859 => x"0a02a908",
			5860 => x"09020204",
			5861 => x"00005be9",
			5862 => x"013c5be9",
			5863 => x"00005be9",
			5864 => x"fedd5be9",
			5865 => x"0c064d0c",
			5866 => x"0c063308",
			5867 => x"08032c04",
			5868 => x"00005be9",
			5869 => x"00615be9",
			5870 => x"fed05be9",
			5871 => x"0d094e04",
			5872 => x"01825be9",
			5873 => x"0c06a40c",
			5874 => x"030b1b04",
			5875 => x"008a5be9",
			5876 => x"0802ee04",
			5877 => x"fe825be9",
			5878 => x"00005be9",
			5879 => x"0c06dc04",
			5880 => x"01665be9",
			5881 => x"00005be9",
			5882 => x"01013f1c",
			5883 => x"020acb04",
			5884 => x"fe665cc5",
			5885 => x"0f0b1714",
			5886 => x"0c061304",
			5887 => x"fef75cc5",
			5888 => x"0c066608",
			5889 => x"040c2404",
			5890 => x"00005cc5",
			5891 => x"019d5cc5",
			5892 => x"0b075f04",
			5893 => x"00005cc5",
			5894 => x"fefa5cc5",
			5895 => x"fe875cc5",
			5896 => x"0c066a28",
			5897 => x"0e0b4224",
			5898 => x"040b5b10",
			5899 => x"0b07630c",
			5900 => x"06018908",
			5901 => x"0e09e004",
			5902 => x"ff445cc5",
			5903 => x"00395cc5",
			5904 => x"fe3a5cc5",
			5905 => x"013d5cc5",
			5906 => x"06019e08",
			5907 => x"0b071004",
			5908 => x"00005cc5",
			5909 => x"02005cc5",
			5910 => x"040c0408",
			5911 => x"0f0ae604",
			5912 => x"00005cc5",
			5913 => x"ff1f5cc5",
			5914 => x"00875cc5",
			5915 => x"fe105cc5",
			5916 => x"0b07b514",
			5917 => x"0601bc10",
			5918 => x"0b07820c",
			5919 => x"0e0b0708",
			5920 => x"0c066d04",
			5921 => x"00005cc5",
			5922 => x"01895cc5",
			5923 => x"fd265cc5",
			5924 => x"01975cc5",
			5925 => x"ffa85cc5",
			5926 => x"0706f504",
			5927 => x"fabd5cc5",
			5928 => x"00039a08",
			5929 => x"0f0afc04",
			5930 => x"00f25cc5",
			5931 => x"fe315cc5",
			5932 => x"0a02a904",
			5933 => x"017d5cc5",
			5934 => x"040d2e04",
			5935 => x"fee65cc5",
			5936 => x"00455cc5",
			5937 => x"020a2d08",
			5938 => x"0b074404",
			5939 => x"fe685d99",
			5940 => x"00005d99",
			5941 => x"01014e38",
			5942 => x"0601a52c",
			5943 => x"040b8e14",
			5944 => x"0c066a0c",
			5945 => x"06018304",
			5946 => x"00005d99",
			5947 => x"0802d804",
			5948 => x"00005d99",
			5949 => x"fe7e5d99",
			5950 => x"01013f04",
			5951 => x"00005d99",
			5952 => x"00f35d99",
			5953 => x"0101230c",
			5954 => x"0f0a7c08",
			5955 => x"09016b04",
			5956 => x"ffb45d99",
			5957 => x"01ae5d99",
			5958 => x"feb35d99",
			5959 => x"0b070e04",
			5960 => x"00005d99",
			5961 => x"0d090f04",
			5962 => x"01bc5d99",
			5963 => x"00005d99",
			5964 => x"0b077108",
			5965 => x"0b073304",
			5966 => x"fef35d99",
			5967 => x"00005d99",
			5968 => x"fe7b5d99",
			5969 => x"0c064d10",
			5970 => x"09022508",
			5971 => x"09022104",
			5972 => x"00005d99",
			5973 => x"00235d99",
			5974 => x"05089404",
			5975 => x"fe6d5d99",
			5976 => x"00005d99",
			5977 => x"0d094e08",
			5978 => x"0b075f04",
			5979 => x"00005d99",
			5980 => x"01945d99",
			5981 => x"0b079104",
			5982 => x"fe1e5d99",
			5983 => x"01016008",
			5984 => x"01015f04",
			5985 => x"00c75d99",
			5986 => x"fe9e5d99",
			5987 => x"08036804",
			5988 => x"017b5d99",
			5989 => x"ff425d99",
			5990 => x"09018b04",
			5991 => x"feeb5e4d",
			5992 => x"0e0aa224",
			5993 => x"040d0e20",
			5994 => x"0901fa08",
			5995 => x"0f0b0904",
			5996 => x"ff865e4d",
			5997 => x"00005e4d",
			5998 => x"0f0a8a0c",
			5999 => x"06017d04",
			6000 => x"00005e4d",
			6001 => x"0c065004",
			6002 => x"ff7e5e4d",
			6003 => x"00005e4d",
			6004 => x"0601a908",
			6005 => x"0d087f04",
			6006 => x"00005e4d",
			6007 => x"00b55e4d",
			6008 => x"00005e4d",
			6009 => x"00c95e4d",
			6010 => x"01016128",
			6011 => x"0b079310",
			6012 => x"0f0aed04",
			6013 => x"00005e4d",
			6014 => x"09020e04",
			6015 => x"00005e4d",
			6016 => x"06018a04",
			6017 => x"00005e4d",
			6018 => x"fed75e4d",
			6019 => x"09022e0c",
			6020 => x"040bbd08",
			6021 => x"01014304",
			6022 => x"00005e4d",
			6023 => x"00a05e4d",
			6024 => x"00005e4d",
			6025 => x"0b07c308",
			6026 => x"0f0afc04",
			6027 => x"00005e4d",
			6028 => x"ff6a5e4d",
			6029 => x"00005e4d",
			6030 => x"0601c208",
			6031 => x"030ada04",
			6032 => x"00005e4d",
			6033 => x"00c75e4d",
			6034 => x"ffd15e4d",
			6035 => x"0c061304",
			6036 => x"fe675ee3",
			6037 => x"01010f04",
			6038 => x"fe935ee3",
			6039 => x"0b07b528",
			6040 => x"0b078218",
			6041 => x"0e0b0710",
			6042 => x"020ac808",
			6043 => x"0b077104",
			6044 => x"ff215ee3",
			6045 => x"01635ee3",
			6046 => x"0601b704",
			6047 => x"016b5ee3",
			6048 => x"feff5ee3",
			6049 => x"01016404",
			6050 => x"fd845ee3",
			6051 => x"013d5ee3",
			6052 => x"0601be0c",
			6053 => x"01014708",
			6054 => x"0f0b2604",
			6055 => x"00005ee3",
			6056 => x"ff685ee3",
			6057 => x"01975ee3",
			6058 => x"fef15ee3",
			6059 => x"0706f504",
			6060 => x"fc545ee3",
			6061 => x"00039a08",
			6062 => x"0f0afc04",
			6063 => x"00d85ee3",
			6064 => x"fe7b5ee3",
			6065 => x"0a02a808",
			6066 => x"01014b04",
			6067 => x"00005ee3",
			6068 => x"01735ee3",
			6069 => x"01017904",
			6070 => x"feb05ee3",
			6071 => x"00525ee3",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1980, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(4056, initial_addr_3'length));
	end generate gen_rom_8;

	gen_rom_9: if SELECT_ROM = 9 generate
		bank <= (
			0 => x"0d05e914",
			1 => x"040df504",
			2 => x"fe7c00b5",
			3 => x"0803dc08",
			4 => x"0a02f304",
			5 => x"000000b5",
			6 => x"004d00b5",
			7 => x"02096604",
			8 => x"ff4300b5",
			9 => x"000000b5",
			10 => x"0c04cc10",
			11 => x"0f089508",
			12 => x"06016f04",
			13 => x"ff9000b5",
			14 => x"019100b5",
			15 => x"0100a104",
			16 => x"feb600b5",
			17 => x"00ab00b5",
			18 => x"0d061118",
			19 => x"040d5510",
			20 => x"0704ea04",
			21 => x"000000b5",
			22 => x"08034404",
			23 => x"000000b5",
			24 => x"0f07c704",
			25 => x"000000b5",
			26 => x"fe7800b5",
			27 => x"06017304",
			28 => x"000000b5",
			29 => x"00dd00b5",
			30 => x"0704f104",
			31 => x"018d00b5",
			32 => x"0b05450c",
			33 => x"06017408",
			34 => x"02092004",
			35 => x"011600b5",
			36 => x"fed100b5",
			37 => x"018d00b5",
			38 => x"0100c308",
			39 => x"0c050d04",
			40 => x"ffe500b5",
			41 => x"fea700b5",
			42 => x"0b063c04",
			43 => x"016f00b5",
			44 => x"001c00b5",
			45 => x"0505b114",
			46 => x"02093508",
			47 => x"0d05dc04",
			48 => x"fe770169",
			49 => x"00000169",
			50 => x"0d05a804",
			51 => x"ff7e0169",
			52 => x"0004bc04",
			53 => x"ffbc0169",
			54 => x"003d0169",
			55 => x"0d0a2b44",
			56 => x"0c04b114",
			57 => x"0704ee0c",
			58 => x"0b052008",
			59 => x"0003fb04",
			60 => x"00000169",
			61 => x"00180169",
			62 => x"ff5e0169",
			63 => x"06016704",
			64 => x"00000169",
			65 => x"01b40169",
			66 => x"0308c720",
			67 => x"0003f210",
			68 => x"0208f008",
			69 => x"03073b04",
			70 => x"ff2f0169",
			71 => x"00b10169",
			72 => x"0c04d004",
			73 => x"000b0169",
			74 => x"fe5a0169",
			75 => x"02093508",
			76 => x"03068304",
			77 => x"ffca0169",
			78 => x"00e20169",
			79 => x"06018104",
			80 => x"fecc0169",
			81 => x"003f0169",
			82 => x"0705a204",
			83 => x"01ba0169",
			84 => x"03090704",
			85 => x"feb20169",
			86 => x"0507f604",
			87 => x"00910169",
			88 => x"00110169",
			89 => x"fe6e0169",
			90 => x"01009540",
			91 => x"040d5528",
			92 => x"0c04ed1c",
			93 => x"0306b90c",
			94 => x"0c049504",
			95 => x"0000028d",
			96 => x"040d2e04",
			97 => x"ff4c028d",
			98 => x"0000028d",
			99 => x"0f086404",
			100 => x"00c5028d",
			101 => x"040bb204",
			102 => x"feed028d",
			103 => x"0f088e04",
			104 => x"004f028d",
			105 => x"0000028d",
			106 => x"0c050a08",
			107 => x"0704ee04",
			108 => x"0000028d",
			109 => x"fea1028d",
			110 => x"0000028d",
			111 => x"0803e608",
			112 => x"06016f04",
			113 => x"0000028d",
			114 => x"0105028d",
			115 => x"040eab04",
			116 => x"ff65028d",
			117 => x"0f070f04",
			118 => x"0000028d",
			119 => x"0209d404",
			120 => x"0025028d",
			121 => x"0000028d",
			122 => x"0e072514",
			123 => x"040bec0c",
			124 => x"0306e204",
			125 => x"0000028d",
			126 => x"06015204",
			127 => x"0000028d",
			128 => x"0147028d",
			129 => x"06018304",
			130 => x"ffd8028d",
			131 => x"0000028d",
			132 => x"0901130c",
			133 => x"06019108",
			134 => x"040a7b04",
			135 => x"0000028d",
			136 => x"ff2a028d",
			137 => x"0000028d",
			138 => x"09013e14",
			139 => x"0f08c608",
			140 => x"0b058304",
			141 => x"0000028d",
			142 => x"ffa8028d",
			143 => x"0e086808",
			144 => x"040aa104",
			145 => x"0000028d",
			146 => x"0132028d",
			147 => x"0000028d",
			148 => x"0f0abc10",
			149 => x"0802eb08",
			150 => x"05083e04",
			151 => x"0000028d",
			152 => x"0091028d",
			153 => x"06019e04",
			154 => x"ff2c028d",
			155 => x"0097028d",
			156 => x"030ac508",
			157 => x"0003a204",
			158 => x"0000028d",
			159 => x"00e2028d",
			160 => x"0601cc04",
			161 => x"0019028d",
			162 => x"ff67028d",
			163 => x"01009544",
			164 => x"0a02d724",
			165 => x"0c04ae08",
			166 => x"0d05e904",
			167 => x"000003b1",
			168 => x"000003b1",
			169 => x"0d061d08",
			170 => x"0704d804",
			171 => x"000003b1",
			172 => x"fef403b1",
			173 => x"0e06ce10",
			174 => x"0c04ec08",
			175 => x"07050804",
			176 => x"00a503b1",
			177 => x"000003b1",
			178 => x"02092804",
			179 => x"000003b1",
			180 => x"ff5c03b1",
			181 => x"fee003b1",
			182 => x"0803e610",
			183 => x"040d1b04",
			184 => x"000003b1",
			185 => x"0305c004",
			186 => x"000003b1",
			187 => x"0d05d104",
			188 => x"000003b1",
			189 => x"00ed03b1",
			190 => x"040eab04",
			191 => x"ff7503b1",
			192 => x"0f070f04",
			193 => x"000003b1",
			194 => x"0209d404",
			195 => x"002303b1",
			196 => x"000003b1",
			197 => x"0e072514",
			198 => x"040bec0c",
			199 => x"0306e204",
			200 => x"000003b1",
			201 => x"0002f604",
			202 => x"000003b1",
			203 => x"013a03b1",
			204 => x"0a02c704",
			205 => x"fffc03b1",
			206 => x"000003b1",
			207 => x"09010f08",
			208 => x"0f08d404",
			209 => x"000003b1",
			210 => x"ff1203b1",
			211 => x"0b07c320",
			212 => x"020af110",
			213 => x"020a5b08",
			214 => x"08034504",
			215 => x"000503b1",
			216 => x"00e103b1",
			217 => x"0901d904",
			218 => x"ff4003b1",
			219 => x"004a03b1",
			220 => x"08038d08",
			221 => x"0c062e04",
			222 => x"012403b1",
			223 => x"002e03b1",
			224 => x"0100ed04",
			225 => x"000003b1",
			226 => x"ffcc03b1",
			227 => x"0901d208",
			228 => x"00042d04",
			229 => x"001e03b1",
			230 => x"000003b1",
			231 => x"00039a04",
			232 => x"000003b1",
			233 => x"09027404",
			234 => x"feff03b1",
			235 => x"000003b1",
			236 => x"0d05e914",
			237 => x"040df504",
			238 => x"fe7f049d",
			239 => x"00051508",
			240 => x"0a02e404",
			241 => x"0000049d",
			242 => x"0048049d",
			243 => x"0a035d04",
			244 => x"ff5d049d",
			245 => x"0000049d",
			246 => x"0601cc54",
			247 => x"0f0af328",
			248 => x"0c04cc10",
			249 => x"0f089508",
			250 => x"06016f04",
			251 => x"ff97049d",
			252 => x"0185049d",
			253 => x"0b055204",
			254 => x"fec2049d",
			255 => x"009d049d",
			256 => x"0c04cd08",
			257 => x"0100a104",
			258 => x"fe33049d",
			259 => x"0043049d",
			260 => x"0507f508",
			261 => x"040a9504",
			262 => x"007f049d",
			263 => x"fffe049d",
			264 => x"0d08b304",
			265 => x"ff21049d",
			266 => x"002a049d",
			267 => x"040c5e18",
			268 => x"0101600c",
			269 => x"0802e304",
			270 => x"0000049d",
			271 => x"00039504",
			272 => x"0000049d",
			273 => x"0124049d",
			274 => x"00039604",
			275 => x"0000049d",
			276 => x"05089704",
			277 => x"0000049d",
			278 => x"ff56049d",
			279 => x"05088604",
			280 => x"fec5049d",
			281 => x"0c068c08",
			282 => x"030b1304",
			283 => x"0000049d",
			284 => x"0153049d",
			285 => x"0a02ab04",
			286 => x"0014049d",
			287 => x"ff6d049d",
			288 => x"0e0b6304",
			289 => x"0000049d",
			290 => x"0e0cf604",
			291 => x"fe38049d",
			292 => x"0601f604",
			293 => x"00c0049d",
			294 => x"ffa3049d",
			295 => x"0f082b40",
			296 => x"03063a1c",
			297 => x"040e6308",
			298 => x"0d066d04",
			299 => x"ff2b05b1",
			300 => x"000005b1",
			301 => x"0b04e304",
			302 => x"000005b1",
			303 => x"02091104",
			304 => x"000005b1",
			305 => x"0209ef08",
			306 => x"0b055404",
			307 => x"007305b1",
			308 => x"000005b1",
			309 => x"000005b1",
			310 => x"06016c18",
			311 => x"0c04cf08",
			312 => x"0900c604",
			313 => x"000005b1",
			314 => x"ff6705b1",
			315 => x"0c04d408",
			316 => x"0d060304",
			317 => x"000005b1",
			318 => x"00a805b1",
			319 => x"09012d04",
			320 => x"ffae05b1",
			321 => x"000005b1",
			322 => x"0208c904",
			323 => x"000005b1",
			324 => x"0d062b04",
			325 => x"011a05b1",
			326 => x"000005b1",
			327 => x"0306c504",
			328 => x"feed05b1",
			329 => x"08037630",
			330 => x"00043620",
			331 => x"0100e710",
			332 => x"0c050708",
			333 => x"06017404",
			334 => x"ff4a05b1",
			335 => x"005705b1",
			336 => x"040c1e04",
			337 => x"fea905b1",
			338 => x"000005b1",
			339 => x"0100ff08",
			340 => x"06015b04",
			341 => x"000005b1",
			342 => x"010e05b1",
			343 => x"0f0ac904",
			344 => x"ffe805b1",
			345 => x"004205b1",
			346 => x"00045408",
			347 => x"0c052e04",
			348 => x"014c05b1",
			349 => x"000005b1",
			350 => x"0a02bc04",
			351 => x"ffb705b1",
			352 => x"000005b1",
			353 => x"0a02db08",
			354 => x"0e06ce04",
			355 => x"000005b1",
			356 => x"fece05b1",
			357 => x"0803e60c",
			358 => x"0c051104",
			359 => x"00e505b1",
			360 => x"09020e04",
			361 => x"ff9905b1",
			362 => x"008005b1",
			363 => x"ff5905b1",
			364 => x"06015b24",
			365 => x"0100ff10",
			366 => x"0a01f70c",
			367 => x"00030204",
			368 => x"fe7106cd",
			369 => x"0e052d04",
			370 => x"000006cd",
			371 => x"022906cd",
			372 => x"fe6406cd",
			373 => x"0601520c",
			374 => x"0d083e08",
			375 => x"07064404",
			376 => x"feff06cd",
			377 => x"017c06cd",
			378 => x"039906cd",
			379 => x"0901c304",
			380 => x"fe9806cd",
			381 => x"005906cd",
			382 => x"0a03235c",
			383 => x"06019938",
			384 => x"040a5b18",
			385 => x"00035b0c",
			386 => x"0a023908",
			387 => x"01013604",
			388 => x"00af06cd",
			389 => x"05f706cd",
			390 => x"fe7e06cd",
			391 => x"0209b708",
			392 => x"0c05fa04",
			393 => x"016306cd",
			394 => x"038c06cd",
			395 => x"fec106cd",
			396 => x"0c04ea10",
			397 => x"0d05e908",
			398 => x"040dca04",
			399 => x"fe9806cd",
			400 => x"016e06cd",
			401 => x"00042804",
			402 => x"008c06cd",
			403 => x"017706cd",
			404 => x"0306e208",
			405 => x"040c8504",
			406 => x"fdfd06cd",
			407 => x"ffce06cd",
			408 => x"07052f04",
			409 => x"012706cd",
			410 => x"ffcd06cd",
			411 => x"07068814",
			412 => x"040d2e0c",
			413 => x"040ca708",
			414 => x"0100fa04",
			415 => x"00ae06cd",
			416 => x"01af06cd",
			417 => x"02df06cd",
			418 => x"0100df04",
			419 => x"011a06cd",
			420 => x"fe7506cd",
			421 => x"0a028a04",
			422 => x"fe8206cd",
			423 => x"030ab104",
			424 => x"fe3b06cd",
			425 => x"0601ab04",
			426 => x"016e06cd",
			427 => x"000006cd",
			428 => x"0c04ce04",
			429 => x"00a606cd",
			430 => x"00053e04",
			431 => x"fcf406cd",
			432 => x"00055404",
			433 => x"006306cd",
			434 => x"fe6e06cd",
			435 => x"03073b48",
			436 => x"0b055638",
			437 => x"0e06f730",
			438 => x"0d061d20",
			439 => x"0704f110",
			440 => x"0505bd08",
			441 => x"02093504",
			442 => x"ff0707f1",
			443 => x"000007f1",
			444 => x"02091104",
			445 => x"00bd07f1",
			446 => x"000007f1",
			447 => x"040c1e08",
			448 => x"0b055204",
			449 => x"feb607f1",
			450 => x"000007f1",
			451 => x"00046304",
			452 => x"001c07f1",
			453 => x"ffce07f1",
			454 => x"0601740c",
			455 => x"0900ec08",
			456 => x"02090904",
			457 => x"00fe07f1",
			458 => x"000007f1",
			459 => x"ff2b07f1",
			460 => x"017107f1",
			461 => x"03071b04",
			462 => x"fea907f1",
			463 => x"000007f1",
			464 => x"06017c08",
			465 => x"02080204",
			466 => x"000007f1",
			467 => x"fe5b07f1",
			468 => x"0d065f04",
			469 => x"004007f1",
			470 => x"ffb507f1",
			471 => x"0506a614",
			472 => x"0003aa04",
			473 => x"000007f1",
			474 => x"09010f0c",
			475 => x"0b056304",
			476 => x"008d07f1",
			477 => x"040be904",
			478 => x"ff8707f1",
			479 => x"000007f1",
			480 => x"010807f1",
			481 => x"09014b0c",
			482 => x"0308c704",
			483 => x"fe6b07f1",
			484 => x"09012d04",
			485 => x"00b507f1",
			486 => x"000007f1",
			487 => x"05077314",
			488 => x"040dca10",
			489 => x"09019608",
			490 => x"0e078e04",
			491 => x"000007f1",
			492 => x"014b07f1",
			493 => x"06018504",
			494 => x"000007f1",
			495 => x"002807f1",
			496 => x"000007f1",
			497 => x"0d07d808",
			498 => x"0901ee04",
			499 => x"fe9f07f1",
			500 => x"000007f1",
			501 => x"0d082508",
			502 => x"0e093304",
			503 => x"000007f1",
			504 => x"00b307f1",
			505 => x"030a9904",
			506 => x"ff7e07f1",
			507 => x"004d07f1",
			508 => x"06015f2c",
			509 => x"01010214",
			510 => x"08027910",
			511 => x"0506f10c",
			512 => x"08023304",
			513 => x"feb80935",
			514 => x"05055804",
			515 => x"00000935",
			516 => x"01e30935",
			517 => x"fe7a0935",
			518 => x"fe650935",
			519 => x"03096810",
			520 => x"02093a0c",
			521 => x"04094504",
			522 => x"01c90935",
			523 => x"0f093304",
			524 => x"feb60935",
			525 => x"003d0935",
			526 => x"02e70935",
			527 => x"02094d04",
			528 => x"00000935",
			529 => x"feef0935",
			530 => x"0c066c54",
			531 => x"06019a30",
			532 => x"040adc1c",
			533 => x"0c05070c",
			534 => x"06016c04",
			535 => x"feb90935",
			536 => x"0c04ed04",
			537 => x"01780935",
			538 => x"02910935",
			539 => x"0d07fd08",
			540 => x"040a1504",
			541 => x"00bb0935",
			542 => x"fe890935",
			543 => x"0d084a04",
			544 => x"01620935",
			545 => x"001b0935",
			546 => x"06016704",
			547 => x"fe6e0935",
			548 => x"0c04cc08",
			549 => x"0b04e304",
			550 => x"fe890935",
			551 => x"01520935",
			552 => x"03066904",
			553 => x"feba0935",
			554 => x"001a0935",
			555 => x"0a02e81c",
			556 => x"05084d10",
			557 => x"0901b208",
			558 => x"08036504",
			559 => x"ffa80935",
			560 => x"01830935",
			561 => x"08030204",
			562 => x"00520935",
			563 => x"01aa0935",
			564 => x"0f0bc908",
			565 => x"0c066a04",
			566 => x"feea0935",
			567 => x"01020935",
			568 => x"015b0935",
			569 => x"0601a604",
			570 => x"01430935",
			571 => x"fec40935",
			572 => x"0d09500c",
			573 => x"0100ff08",
			574 => x"0508cf04",
			575 => x"fff00935",
			576 => x"01120935",
			577 => x"fe6f0935",
			578 => x"0803b414",
			579 => x"020ae608",
			580 => x"0f0afc04",
			581 => x"ff190935",
			582 => x"05080935",
			583 => x"0d096904",
			584 => x"fe8e0935",
			585 => x"0901d204",
			586 => x"02370935",
			587 => x"00560935",
			588 => x"fe560935",
			589 => x"0505db18",
			590 => x"040c9304",
			591 => x"fe640a49",
			592 => x"0d05a804",
			593 => x"fe960a49",
			594 => x"0f080e0c",
			595 => x"06017008",
			596 => x"0c04b204",
			597 => x"005b0a49",
			598 => x"ffb60a49",
			599 => x"01790a49",
			600 => x"fedc0a49",
			601 => x"0505f61c",
			602 => x"0d060f14",
			603 => x"0b053308",
			604 => x"01007e04",
			605 => x"00000a49",
			606 => x"fea40a49",
			607 => x"06016404",
			608 => x"00000a49",
			609 => x"02090504",
			610 => x"01950a49",
			611 => x"00000a49",
			612 => x"06016304",
			613 => x"00000a49",
			614 => x"019a0a49",
			615 => x"0d061f1c",
			616 => x"040cc610",
			617 => x"0f08460c",
			618 => x"01009208",
			619 => x"00046304",
			620 => x"fdff0a49",
			621 => x"00000a49",
			622 => x"00800a49",
			623 => x"fd870a49",
			624 => x"02098108",
			625 => x"0c052804",
			626 => x"011f0a49",
			627 => x"00000a49",
			628 => x"00000a49",
			629 => x"0b05561c",
			630 => x"0f087210",
			631 => x"0003ed08",
			632 => x"05060604",
			633 => x"ffd00a49",
			634 => x"001b0a49",
			635 => x"05060804",
			636 => x"02160a49",
			637 => x"00e90a49",
			638 => x"06017904",
			639 => x"fece0a49",
			640 => x"02096604",
			641 => x"01a00a49",
			642 => x"00540a49",
			643 => x"0e06ce10",
			644 => x"00037d08",
			645 => x"0c054c04",
			646 => x"00000a49",
			647 => x"00210a49",
			648 => x"06018104",
			649 => x"fdcd0a49",
			650 => x"00000a49",
			651 => x"05062608",
			652 => x"0a029004",
			653 => x"ffed0a49",
			654 => x"016b0a49",
			655 => x"09014704",
			656 => x"ff500a49",
			657 => x"003e0a49",
			658 => x"06015b24",
			659 => x"0100ff10",
			660 => x"0a01f70c",
			661 => x"00030204",
			662 => x"fe6e0b85",
			663 => x"0e052d04",
			664 => x"00000b85",
			665 => x"025f0b85",
			666 => x"fe640b85",
			667 => x"0601520c",
			668 => x"0d083e08",
			669 => x"07064404",
			670 => x"feea0b85",
			671 => x"01b50b85",
			672 => x"04cf0b85",
			673 => x"0901c304",
			674 => x"fe8d0b85",
			675 => x"00800b85",
			676 => x"0c066c54",
			677 => x"06019930",
			678 => x"03063210",
			679 => x"06017404",
			680 => x"fe6a0b85",
			681 => x"07051808",
			682 => x"0d05ca04",
			683 => x"00540b85",
			684 => x"01e80b85",
			685 => x"fdfe0b85",
			686 => x"0c04ea10",
			687 => x"06017408",
			688 => x"0900d904",
			689 => x"017e0b85",
			690 => x"ff9c0b85",
			691 => x"0306b904",
			692 => x"00db0b85",
			693 => x"01910b85",
			694 => x"0306e208",
			695 => x"040c8504",
			696 => x"fded0b85",
			697 => x"ffdf0b85",
			698 => x"0b058304",
			699 => x"01690b85",
			700 => x"001d0b85",
			701 => x"040d2e18",
			702 => x"0b07330c",
			703 => x"0a027804",
			704 => x"00000b85",
			705 => x"09015504",
			706 => x"00680b85",
			707 => x"01c20b85",
			708 => x"09021b04",
			709 => x"fe190b85",
			710 => x"01016304",
			711 => x"024e0b85",
			712 => x"004d0b85",
			713 => x"09011b04",
			714 => x"016e0b85",
			715 => x"040d8804",
			716 => x"ffc10b85",
			717 => x"fe350b85",
			718 => x"0d094e08",
			719 => x"06017d04",
			720 => x"00270b85",
			721 => x"fe6a0b85",
			722 => x"0706e004",
			723 => x"12020b85",
			724 => x"0e0b0e10",
			725 => x"0b07b508",
			726 => x"0e0aa204",
			727 => x"00d70b85",
			728 => x"fe940b85",
			729 => x"09022e04",
			730 => x"011f0b85",
			731 => x"04cd0b85",
			732 => x"0004a708",
			733 => x"0b082804",
			734 => x"febc0b85",
			735 => x"00eb0b85",
			736 => x"fe520b85",
			737 => x"0505cc18",
			738 => x"040d6e04",
			739 => x"fe770cb9",
			740 => x"0b051110",
			741 => x"02093d04",
			742 => x"ff200cb9",
			743 => x"0209b108",
			744 => x"05050f04",
			745 => x"00000cb9",
			746 => x"00610cb9",
			747 => x"ffaf0cb9",
			748 => x"00f40cb9",
			749 => x"0f08223c",
			750 => x"0705081c",
			751 => x"0a02a60c",
			752 => x"0c04d104",
			753 => x"fe9c0cb9",
			754 => x"0c04d204",
			755 => x"01400cb9",
			756 => x"00000cb9",
			757 => x"0e059604",
			758 => x"00000cb9",
			759 => x"06016304",
			760 => x"00000cb9",
			761 => x"0c04d404",
			762 => x"01b00cb9",
			763 => x"00aa0cb9",
			764 => x"0e06e218",
			765 => x"0f080e0c",
			766 => x"0b054304",
			767 => x"00000cb9",
			768 => x"02080204",
			769 => x"00000cb9",
			770 => x"fe570cb9",
			771 => x"00048a04",
			772 => x"ffb60cb9",
			773 => x"0b058704",
			774 => x"00a50cb9",
			775 => x"00000cb9",
			776 => x"06011d04",
			777 => x"00000cb9",
			778 => x"01450cb9",
			779 => x"01009724",
			780 => x"0f086414",
			781 => x"07050808",
			782 => x"06016f04",
			783 => x"ff990cb9",
			784 => x"016d0cb9",
			785 => x"00042804",
			786 => x"fd750cb9",
			787 => x"0a02cf04",
			788 => x"ffa20cb9",
			789 => x"00000cb9",
			790 => x"0c04ef0c",
			791 => x"040bb204",
			792 => x"fdef0cb9",
			793 => x"00045b04",
			794 => x"00000cb9",
			795 => x"fec70cb9",
			796 => x"00000cb9",
			797 => x"0506150c",
			798 => x"0d063708",
			799 => x"0c04cf04",
			800 => x"00f30cb9",
			801 => x"ff620cb9",
			802 => x"01820cb9",
			803 => x"0901200c",
			804 => x"0d063f04",
			805 => x"00830cb9",
			806 => x"02097b04",
			807 => x"fe760cb9",
			808 => x"00000cb9",
			809 => x"05066c04",
			810 => x"01900cb9",
			811 => x"0d09f804",
			812 => x"fffa0cb9",
			813 => x"fe920cb9",
			814 => x"0b05110c",
			815 => x"02096c04",
			816 => x"fe680d8d",
			817 => x"00052904",
			818 => x"ff6a0d8d",
			819 => x"01300d8d",
			820 => x"0a032358",
			821 => x"0100a834",
			822 => x"0003f218",
			823 => x"07050308",
			824 => x"0003e604",
			825 => x"feea0d8d",
			826 => x"f9e90d8d",
			827 => x"0c04e708",
			828 => x"0a027204",
			829 => x"ff660d8d",
			830 => x"012e0d8d",
			831 => x"0c054804",
			832 => x"fe2e0d8d",
			833 => x"01010d8d",
			834 => x"040cc610",
			835 => x"0b056908",
			836 => x"0306b904",
			837 => x"ff560d8d",
			838 => x"008c0d8d",
			839 => x"0b057604",
			840 => x"fbb30d8d",
			841 => x"fe9e0d8d",
			842 => x"0c050d08",
			843 => x"03069604",
			844 => x"00d20d8d",
			845 => x"02080d8d",
			846 => x"fea80d8d",
			847 => x"05065104",
			848 => x"01a10d8d",
			849 => x"09014b10",
			850 => x"0705a208",
			851 => x"0a02d104",
			852 => x"fdf00d8d",
			853 => x"00000d8d",
			854 => x"040acf04",
			855 => x"01430d8d",
			856 => x"fe5a0d8d",
			857 => x"0a021d08",
			858 => x"0901a104",
			859 => x"ffa60d8d",
			860 => x"01c30d8d",
			861 => x"0f0aed04",
			862 => x"00110d8d",
			863 => x"00b50d8d",
			864 => x"0c04e904",
			865 => x"01320d8d",
			866 => x"fe1f0d8d",
			867 => x"040a5b38",
			868 => x"0b06bc18",
			869 => x"0a027814",
			870 => x"0802aa0c",
			871 => x"040a0108",
			872 => x"00034604",
			873 => x"ff1d0ed9",
			874 => x"00000ed9",
			875 => x"00bb0ed9",
			876 => x"0409b304",
			877 => x"00000ed9",
			878 => x"fee30ed9",
			879 => x"00a70ed9",
			880 => x"07065b14",
			881 => x"0901f810",
			882 => x"0100ff04",
			883 => x"00000ed9",
			884 => x"07062b04",
			885 => x"00000ed9",
			886 => x"0507f504",
			887 => x"01360ed9",
			888 => x"00000ed9",
			889 => x"00000ed9",
			890 => x"06016308",
			891 => x"06015e04",
			892 => x"ff790ed9",
			893 => x"00ad0ed9",
			894 => x"ff650ed9",
			895 => x"040b463c",
			896 => x"0100a618",
			897 => x"0003f204",
			898 => x"fe310ed9",
			899 => x"0505f90c",
			900 => x"08033704",
			901 => x"00000ed9",
			902 => x"00042004",
			903 => x"fe3b0ed9",
			904 => x"00000ed9",
			905 => x"07051804",
			906 => x"00fe0ed9",
			907 => x"00000ed9",
			908 => x"0b058304",
			909 => x"012e0ed9",
			910 => x"0003a310",
			911 => x"00039a08",
			912 => x"040adc04",
			913 => x"000c0ed9",
			914 => x"ff3e0ed9",
			915 => x"06018904",
			916 => x"00000ed9",
			917 => x"00e00ed9",
			918 => x"0901d908",
			919 => x"040ae804",
			920 => x"fff00ed9",
			921 => x"fdfd0ed9",
			922 => x"0b070e04",
			923 => x"00df0ed9",
			924 => x"ff3b0ed9",
			925 => x"06016304",
			926 => x"fed40ed9",
			927 => x"0704ef14",
			928 => x"0505bd0c",
			929 => x"0b04e304",
			930 => x"ffd40ed9",
			931 => x"040d5504",
			932 => x"00000ed9",
			933 => x"00120ed9",
			934 => x"0d060304",
			935 => x"00540ed9",
			936 => x"01700ed9",
			937 => x"0803a010",
			938 => x"040bca08",
			939 => x"08036104",
			940 => x"00430ed9",
			941 => x"fea00ed9",
			942 => x"03067804",
			943 => x"ff7a0ed9",
			944 => x"00730ed9",
			945 => x"0e059608",
			946 => x"0d05e904",
			947 => x"00000ed9",
			948 => x"00660ed9",
			949 => x"fef60ed9",
			950 => x"06015b28",
			951 => x"0100ff14",
			952 => x"0a01f710",
			953 => x"0802690c",
			954 => x"04097204",
			955 => x"fe73101d",
			956 => x"03098704",
			957 => x"002f101d",
			958 => x"0000101d",
			959 => x"01e9101d",
			960 => x"fe65101d",
			961 => x"0601520c",
			962 => x"0d083e08",
			963 => x"07064404",
			964 => x"ff0f101d",
			965 => x"0161101d",
			966 => x"030e101d",
			967 => x"0901c304",
			968 => x"fea3101d",
			969 => x"0059101d",
			970 => x"0a03236c",
			971 => x"0601993c",
			972 => x"040a5b1c",
			973 => x"0901c30c",
			974 => x"02099508",
			975 => x"0f096804",
			976 => x"0179101d",
			977 => x"febb101d",
			978 => x"034e101d",
			979 => x"0507e408",
			980 => x"0e090704",
			981 => x"fe8b101d",
			982 => x"01cc101d",
			983 => x"0d087404",
			984 => x"fe75101d",
			985 => x"01d9101d",
			986 => x"0c04ea10",
			987 => x"0d05e908",
			988 => x"040dca04",
			989 => x"fe9f101d",
			990 => x"0156101d",
			991 => x"06017404",
			992 => x"0047101d",
			993 => x"014f101d",
			994 => x"0306e208",
			995 => x"040c8504",
			996 => x"fe06101d",
			997 => x"ffd5101d",
			998 => x"05063504",
			999 => x"0133101d",
			1000 => x"ffd3101d",
			1001 => x"07068814",
			1002 => x"040d2e0c",
			1003 => x"09015504",
			1004 => x"002f101d",
			1005 => x"0802ff04",
			1006 => x"0000101d",
			1007 => x"01b5101d",
			1008 => x"0100df04",
			1009 => x"0103101d",
			1010 => x"fe83101d",
			1011 => x"0e0b7710",
			1012 => x"0d098508",
			1013 => x"05086a04",
			1014 => x"0009101d",
			1015 => x"fe9a101d",
			1016 => x"0c06c704",
			1017 => x"027d101d",
			1018 => x"0000101d",
			1019 => x"0706f504",
			1020 => x"0248101d",
			1021 => x"040d6e04",
			1022 => x"ff8b101d",
			1023 => x"0177101d",
			1024 => x"0c04ce04",
			1025 => x"008b101d",
			1026 => x"0900c408",
			1027 => x"01002304",
			1028 => x"fe97101d",
			1029 => x"007a101d",
			1030 => x"fe2e101d",
			1031 => x"0b051110",
			1032 => x"02093d04",
			1033 => x"fe941129",
			1034 => x"0209b108",
			1035 => x"0d05a804",
			1036 => x"00001129",
			1037 => x"00241129",
			1038 => x"ffb41129",
			1039 => x"0b055638",
			1040 => x"0d064430",
			1041 => x"040bb214",
			1042 => x"08036510",
			1043 => x"0306b908",
			1044 => x"0704d404",
			1045 => x"00001129",
			1046 => x"fe921129",
			1047 => x"0208f904",
			1048 => x"01741129",
			1049 => x"ffa91129",
			1050 => x"fe711129",
			1051 => x"0c04d00c",
			1052 => x"02097b08",
			1053 => x"0505cc04",
			1054 => x"006f1129",
			1055 => x"01981129",
			1056 => x"00001129",
			1057 => x"03067808",
			1058 => x"040e6304",
			1059 => x"fe851129",
			1060 => x"00831129",
			1061 => x"02096004",
			1062 => x"01031129",
			1063 => x"ffb51129",
			1064 => x"0a029204",
			1065 => x"00001129",
			1066 => x"019e1129",
			1067 => x"0c04cf0c",
			1068 => x"040b5608",
			1069 => x"06017804",
			1070 => x"00001129",
			1071 => x"00f01129",
			1072 => x"fdb81129",
			1073 => x"040b1614",
			1074 => x"08033310",
			1075 => x"0c056608",
			1076 => x"040a7b04",
			1077 => x"00001129",
			1078 => x"fe4f1129",
			1079 => x"0a025904",
			1080 => x"00001129",
			1081 => x"00f01129",
			1082 => x"01961129",
			1083 => x"030a9910",
			1084 => x"0a02a908",
			1085 => x"0003ee04",
			1086 => x"ff891129",
			1087 => x"fe1b1129",
			1088 => x"040c5204",
			1089 => x"01111129",
			1090 => x"ff281129",
			1091 => x"08037308",
			1092 => x"0802e804",
			1093 => x"ff571129",
			1094 => x"00a81129",
			1095 => x"040d6e04",
			1096 => x"fefe1129",
			1097 => x"00ea1129",
			1098 => x"09012740",
			1099 => x"07051f28",
			1100 => x"0c050720",
			1101 => x"0f08e61c",
			1102 => x"01009510",
			1103 => x"040bb208",
			1104 => x"0f084f04",
			1105 => x"00001255",
			1106 => x"fe221255",
			1107 => x"0d060f04",
			1108 => x"ffd81255",
			1109 => x"01191255",
			1110 => x"06016c04",
			1111 => x"ff621255",
			1112 => x"07050304",
			1113 => x"00001255",
			1114 => x"01871255",
			1115 => x"fea91255",
			1116 => x"0a02d404",
			1117 => x"fe1c1255",
			1118 => x"00001255",
			1119 => x"07055f08",
			1120 => x"020a2004",
			1121 => x"fe9f1255",
			1122 => x"00001255",
			1123 => x"0a02fd0c",
			1124 => x"05069b04",
			1125 => x"00001255",
			1126 => x"02088b04",
			1127 => x"00001255",
			1128 => x"00f01255",
			1129 => x"ff5d1255",
			1130 => x"05067e04",
			1131 => x"01841255",
			1132 => x"0308c718",
			1133 => x"040bde08",
			1134 => x"02091b04",
			1135 => x"00001255",
			1136 => x"fe681255",
			1137 => x"040dca0c",
			1138 => x"07057708",
			1139 => x"0209d404",
			1140 => x"00001255",
			1141 => x"01531255",
			1142 => x"00001255",
			1143 => x"ff901255",
			1144 => x"0309781c",
			1145 => x"0f096010",
			1146 => x"08025a08",
			1147 => x"0100f804",
			1148 => x"00001255",
			1149 => x"01071255",
			1150 => x"01011104",
			1151 => x"ff231255",
			1152 => x"00001255",
			1153 => x"020a8608",
			1154 => x"0901ec04",
			1155 => x"01971255",
			1156 => x"00001255",
			1157 => x"ffdf1255",
			1158 => x"0507ca10",
			1159 => x"0c05f308",
			1160 => x"01010b04",
			1161 => x"00001255",
			1162 => x"01191255",
			1163 => x"06018904",
			1164 => x"ff121255",
			1165 => x"007a1255",
			1166 => x"0c05f808",
			1167 => x"01014104",
			1168 => x"fef31255",
			1169 => x"00001255",
			1170 => x"0c061204",
			1171 => x"00cb1255",
			1172 => x"00001255",
			1173 => x"0f0ab278",
			1174 => x"0f0a7c64",
			1175 => x"0f084638",
			1176 => x"0306781c",
			1177 => x"040df510",
			1178 => x"0704ec08",
			1179 => x"0505bd04",
			1180 => x"ff1413c1",
			1181 => x"00d313c1",
			1182 => x"0b05a804",
			1183 => x"feb513c1",
			1184 => x"000013c1",
			1185 => x"0505f908",
			1186 => x"0d05ca04",
			1187 => x"000013c1",
			1188 => x"011713c1",
			1189 => x"ff7f13c1",
			1190 => x"0705080c",
			1191 => x"0d060304",
			1192 => x"000013c1",
			1193 => x"06016304",
			1194 => x"000013c1",
			1195 => x"014313c1",
			1196 => x"08037c08",
			1197 => x"01009d04",
			1198 => x"fedd13c1",
			1199 => x"000013c1",
			1200 => x"0c050704",
			1201 => x"00a613c1",
			1202 => x"000013c1",
			1203 => x"03071b14",
			1204 => x"0601810c",
			1205 => x"0b055408",
			1206 => x"040b6904",
			1207 => x"004d13c1",
			1208 => x"ff2513c1",
			1209 => x"fe5513c1",
			1210 => x"040c3204",
			1211 => x"000013c1",
			1212 => x"009413c1",
			1213 => x"0b055608",
			1214 => x"08032c04",
			1215 => x"000013c1",
			1216 => x"014f13c1",
			1217 => x"01009b08",
			1218 => x"03075404",
			1219 => x"fff713c1",
			1220 => x"014b13c1",
			1221 => x"0308c704",
			1222 => x"ff7213c1",
			1223 => x"000013c1",
			1224 => x"01012a04",
			1225 => x"fe2113c1",
			1226 => x"0b06ff04",
			1227 => x"004713c1",
			1228 => x"0b075f04",
			1229 => x"ff5413c1",
			1230 => x"040b0404",
			1231 => x"000013c1",
			1232 => x"000413c1",
			1233 => x"0a02d12c",
			1234 => x"0b071008",
			1235 => x"0f0ac304",
			1236 => x"000013c1",
			1237 => x"016113c1",
			1238 => x"040cc61c",
			1239 => x"0b07b510",
			1240 => x"040b1508",
			1241 => x"01015004",
			1242 => x"00e513c1",
			1243 => x"000013c1",
			1244 => x"01011304",
			1245 => x"000013c1",
			1246 => x"ff1513c1",
			1247 => x"08031e08",
			1248 => x"0d095b04",
			1249 => x"000013c1",
			1250 => x"00f313c1",
			1251 => x"000013c1",
			1252 => x"00043504",
			1253 => x"014113c1",
			1254 => x"000013c1",
			1255 => x"0f0d4b0c",
			1256 => x"020bbc04",
			1257 => x"000013c1",
			1258 => x"0601cc04",
			1259 => x"000013c1",
			1260 => x"fe7013c1",
			1261 => x"0a032304",
			1262 => x"011813c1",
			1263 => x"000013c1",
			1264 => x"06017060",
			1265 => x"0f09563c",
			1266 => x"06016424",
			1267 => x"0100fc10",
			1268 => x"01009304",
			1269 => x"fe511565",
			1270 => x"0900ec04",
			1271 => x"02cd1565",
			1272 => x"08026f04",
			1273 => x"fe5d1565",
			1274 => x"ffe91565",
			1275 => x"08025f04",
			1276 => x"05511565",
			1277 => x"0e08e108",
			1278 => x"0901a104",
			1279 => x"01a81565",
			1280 => x"fe621565",
			1281 => x"0d082204",
			1282 => x"059d1565",
			1283 => x"fe751565",
			1284 => x"02090014",
			1285 => x"03063a04",
			1286 => x"fe5c1565",
			1287 => x"040b7d08",
			1288 => x"0306c504",
			1289 => x"fe7d1565",
			1290 => x"042d1565",
			1291 => x"0c04ed04",
			1292 => x"0bb31565",
			1293 => x"00fe1565",
			1294 => x"fe581565",
			1295 => x"0c05f610",
			1296 => x"02096004",
			1297 => x"0a821565",
			1298 => x"0f09b108",
			1299 => x"07065504",
			1300 => x"fe711565",
			1301 => x"00d81565",
			1302 => x"05161565",
			1303 => x"040a280c",
			1304 => x"0b06dd08",
			1305 => x"08029104",
			1306 => x"04cd1565",
			1307 => x"fe7e1565",
			1308 => x"fe5d1565",
			1309 => x"040a5b04",
			1310 => x"0a271565",
			1311 => x"002d1565",
			1312 => x"0c064d48",
			1313 => x"0a026120",
			1314 => x"06018110",
			1315 => x"0901bc04",
			1316 => x"06531565",
			1317 => x"0a023004",
			1318 => x"034a1565",
			1319 => x"07064104",
			1320 => x"fe801565",
			1321 => x"ffb31565",
			1322 => x"07062e04",
			1323 => x"08e41565",
			1324 => x"06018304",
			1325 => x"05fb1565",
			1326 => x"01014504",
			1327 => x"ffae1565",
			1328 => x"04211565",
			1329 => x"040fc620",
			1330 => x"06017910",
			1331 => x"07052f08",
			1332 => x"0b051204",
			1333 => x"fe8c1565",
			1334 => x"05d51565",
			1335 => x"08030604",
			1336 => x"02861565",
			1337 => x"fe601565",
			1338 => x"07069b08",
			1339 => x"07051f04",
			1340 => x"069d1565",
			1341 => x"05b31565",
			1342 => x"020b3204",
			1343 => x"fe791565",
			1344 => x"04961565",
			1345 => x"0c04e704",
			1346 => x"03051565",
			1347 => x"fe6a1565",
			1348 => x"0c066c18",
			1349 => x"0601a610",
			1350 => x"01014d0c",
			1351 => x"0706cb08",
			1352 => x"0901ff04",
			1353 => x"fe831565",
			1354 => x"00f81565",
			1355 => x"060a1565",
			1356 => x"fe581565",
			1357 => x"01014e04",
			1358 => x"00351565",
			1359 => x"0b441565",
			1360 => x"01018e10",
			1361 => x"09026b0c",
			1362 => x"06017d04",
			1363 => x"00001565",
			1364 => x"0706b704",
			1365 => x"ff401565",
			1366 => x"fe681565",
			1367 => x"00091565",
			1368 => x"03aa1565",
			1369 => x"06017454",
			1370 => x"0505cc04",
			1371 => x"fe9916a1",
			1372 => x"0f080e24",
			1373 => x"0a02a614",
			1374 => x"0208020c",
			1375 => x"0c054c04",
			1376 => x"000016a1",
			1377 => x"0506e204",
			1378 => x"00bc16a1",
			1379 => x"000016a1",
			1380 => x"0f080504",
			1381 => x"fed116a1",
			1382 => x"000016a1",
			1383 => x"06016404",
			1384 => x"000016a1",
			1385 => x"0c04ef08",
			1386 => x"0e059604",
			1387 => x"000016a1",
			1388 => x"014c16a1",
			1389 => x"000016a1",
			1390 => x"040adc18",
			1391 => x"09011b08",
			1392 => x"040aa904",
			1393 => x"000016a1",
			1394 => x"011f16a1",
			1395 => x"0901d408",
			1396 => x"07069b04",
			1397 => x"ff4616a1",
			1398 => x"002616a1",
			1399 => x"0802aa04",
			1400 => x"00d116a1",
			1401 => x"ffb916a1",
			1402 => x"0209190c",
			1403 => x"0208e404",
			1404 => x"ff6916a1",
			1405 => x"0c04ec04",
			1406 => x"002b16a1",
			1407 => x"000016a1",
			1408 => x"0c05d504",
			1409 => x"fe6616a1",
			1410 => x"000016a1",
			1411 => x"07051818",
			1412 => x"0b055214",
			1413 => x"0f088510",
			1414 => x"0900e70c",
			1415 => x"040c5e04",
			1416 => x"fec216a1",
			1417 => x"02097004",
			1418 => x"015316a1",
			1419 => x"000016a1",
			1420 => x"016f16a1",
			1421 => x"ff1716a1",
			1422 => x"018d16a1",
			1423 => x"0c04cd08",
			1424 => x"08033104",
			1425 => x"000016a1",
			1426 => x"fe5016a1",
			1427 => x"00047d1c",
			1428 => x"0a02bf10",
			1429 => x"08036308",
			1430 => x"0c050504",
			1431 => x"011816a1",
			1432 => x"fff916a1",
			1433 => x"0f08dd04",
			1434 => x"000016a1",
			1435 => x"fd7a16a1",
			1436 => x"0c061504",
			1437 => x"019016a1",
			1438 => x"0f0c3904",
			1439 => x"fe9e16a1",
			1440 => x"00d716a1",
			1441 => x"07051f04",
			1442 => x"002916a1",
			1443 => x"0e0d3b04",
			1444 => x"fe8216a1",
			1445 => x"0c071804",
			1446 => x"002e16a1",
			1447 => x"000016a1",
			1448 => x"0e078e54",
			1449 => x"0b05562c",
			1450 => x"040ad50c",
			1451 => x"0c04d204",
			1452 => x"00001815",
			1453 => x"0d063704",
			1454 => x"fe821815",
			1455 => x"00001815",
			1456 => x"0306b910",
			1457 => x"0a02a904",
			1458 => x"fee71815",
			1459 => x"0f082b08",
			1460 => x"03063a04",
			1461 => x"ffb11815",
			1462 => x"00a81815",
			1463 => x"ff1f1815",
			1464 => x"0f088e08",
			1465 => x"0d061104",
			1466 => x"00001815",
			1467 => x"01651815",
			1468 => x"0d063f04",
			1469 => x"fed11815",
			1470 => x"00891815",
			1471 => x"0100a614",
			1472 => x"0d062d04",
			1473 => x"00001815",
			1474 => x"06018d0c",
			1475 => x"0600e804",
			1476 => x"00001815",
			1477 => x"0a02c704",
			1478 => x"fe7b1815",
			1479 => x"00001815",
			1480 => x"00001815",
			1481 => x"0b058304",
			1482 => x"00861815",
			1483 => x"06015e0c",
			1484 => x"0c056604",
			1485 => x"00001815",
			1486 => x"0d06c704",
			1487 => x"00651815",
			1488 => x"00001815",
			1489 => x"ff3c1815",
			1490 => x"0f09e134",
			1491 => x"06018c30",
			1492 => x"0f095618",
			1493 => x"02091910",
			1494 => x"0e081608",
			1495 => x"07060204",
			1496 => x"00d71815",
			1497 => x"00001815",
			1498 => x"0b06cc04",
			1499 => x"ffa91815",
			1500 => x"00001815",
			1501 => x"0b058304",
			1502 => x"00001815",
			1503 => x"fedc1815",
			1504 => x"0309780c",
			1505 => x"01013408",
			1506 => x"03091a04",
			1507 => x"00001815",
			1508 => x"00ed1815",
			1509 => x"00001815",
			1510 => x"07064204",
			1511 => x"ff761815",
			1512 => x"0409db04",
			1513 => x"00001815",
			1514 => x"00751815",
			1515 => x"01161815",
			1516 => x"0308ff04",
			1517 => x"feef1815",
			1518 => x"01011f14",
			1519 => x"0803900c",
			1520 => x"08033408",
			1521 => x"0a028b04",
			1522 => x"007c1815",
			1523 => x"ff441815",
			1524 => x"01011815",
			1525 => x"0100ed04",
			1526 => x"00001815",
			1527 => x"ffcd1815",
			1528 => x"01012a0c",
			1529 => x"0a02b608",
			1530 => x"0b06e004",
			1531 => x"00001815",
			1532 => x"fe4e1815",
			1533 => x"00001815",
			1534 => x"040c5e08",
			1535 => x"00037d04",
			1536 => x"ff9b1815",
			1537 => x"00681815",
			1538 => x"0a02e104",
			1539 => x"ff0e1815",
			1540 => x"001c1815",
			1541 => x"06016c58",
			1542 => x"09019634",
			1543 => x"06016720",
			1544 => x"0600e808",
			1545 => x"00030204",
			1546 => x"fe7f19b1",
			1547 => x"034719b1",
			1548 => x"0601630c",
			1549 => x"0e06e204",
			1550 => x"fe5d19b1",
			1551 => x"0d070804",
			1552 => x"012019b1",
			1553 => x"fe6019b1",
			1554 => x"0e060f04",
			1555 => x"fe6c19b1",
			1556 => x"0e064304",
			1557 => x"022219b1",
			1558 => x"fe9019b1",
			1559 => x"02090c10",
			1560 => x"0e05e004",
			1561 => x"fe7819b1",
			1562 => x"0a02ac08",
			1563 => x"0003fb04",
			1564 => x"00a519b1",
			1565 => x"fe7d19b1",
			1566 => x"02e319b1",
			1567 => x"fe6a19b1",
			1568 => x"0e08fd0c",
			1569 => x"0705e808",
			1570 => x"040a1504",
			1571 => x"04fc19b1",
			1572 => x"fec119b1",
			1573 => x"fe6819b1",
			1574 => x"0c05f208",
			1575 => x"0507b804",
			1576 => x"004b19b1",
			1577 => x"fe4c19b1",
			1578 => x"040a280c",
			1579 => x"0507f508",
			1580 => x"0a021d04",
			1581 => x"036919b1",
			1582 => x"ffa719b1",
			1583 => x"fe7819b1",
			1584 => x"052919b1",
			1585 => x"0b07634c",
			1586 => x"0802e820",
			1587 => x"040af51c",
			1588 => x"0901d20c",
			1589 => x"0c05f508",
			1590 => x"06017004",
			1591 => x"fe3c19b1",
			1592 => x"019019b1",
			1593 => x"047419b1",
			1594 => x"0a024908",
			1595 => x"0a023904",
			1596 => x"005219b1",
			1597 => x"fe6519b1",
			1598 => x"0b06ee04",
			1599 => x"021319b1",
			1600 => x"ff0019b1",
			1601 => x"fe4319b1",
			1602 => x"040c6014",
			1603 => x"0d05ed04",
			1604 => x"fe2a19b1",
			1605 => x"0100c208",
			1606 => x"07052f04",
			1607 => x"020a19b1",
			1608 => x"fecf19b1",
			1609 => x"00039604",
			1610 => x"003f19b1",
			1611 => x"023219b1",
			1612 => x"0c04f10c",
			1613 => x"0505a004",
			1614 => x"fe8119b1",
			1615 => x"0900b104",
			1616 => x"03e219b1",
			1617 => x"01f219b1",
			1618 => x"06018104",
			1619 => x"fe6419b1",
			1620 => x"0c054604",
			1621 => x"018319b1",
			1622 => x"ff0b19b1",
			1623 => x"09025824",
			1624 => x"0706c90c",
			1625 => x"0d092204",
			1626 => x"fe6e19b1",
			1627 => x"0e0adc04",
			1628 => x"069819b1",
			1629 => x"008419b1",
			1630 => x"0101300c",
			1631 => x"0a02ab08",
			1632 => x"0d095604",
			1633 => x"006d19b1",
			1634 => x"067f19b1",
			1635 => x"fe6119b1",
			1636 => x"0d097504",
			1637 => x"fe5f19b1",
			1638 => x"0e0b0e04",
			1639 => x"067219b1",
			1640 => x"fe7a19b1",
			1641 => x"0e0c4a04",
			1642 => x"fe8919b1",
			1643 => x"022219b1",
			1644 => x"0601673c",
			1645 => x"0100fa1c",
			1646 => x"0600e808",
			1647 => x"01009b04",
			1648 => x"fe851b25",
			1649 => x"02d61b25",
			1650 => x"0e060f04",
			1651 => x"fe5f1b25",
			1652 => x"0d07080c",
			1653 => x"0705bb08",
			1654 => x"00047004",
			1655 => x"fec51b25",
			1656 => x"01c51b25",
			1657 => x"050d1b25",
			1658 => x"fe611b25",
			1659 => x"0f096810",
			1660 => x"0e086804",
			1661 => x"01941b25",
			1662 => x"0e08fd04",
			1663 => x"fe701b25",
			1664 => x"0507ca04",
			1665 => x"016c1b25",
			1666 => x"fe961b25",
			1667 => x"05084d0c",
			1668 => x"0507f508",
			1669 => x"0507e604",
			1670 => x"00711b25",
			1671 => x"058e1b25",
			1672 => x"fe701b25",
			1673 => x"05051b25",
			1674 => x"0c066c5c",
			1675 => x"06018d38",
			1676 => x"07051f1c",
			1677 => x"0d05ed0c",
			1678 => x"040df508",
			1679 => x"0f077b04",
			1680 => x"fff71b25",
			1681 => x"fe3d1b25",
			1682 => x"02551b25",
			1683 => x"0f087208",
			1684 => x"0d061104",
			1685 => x"01941b25",
			1686 => x"027f1b25",
			1687 => x"0900ec04",
			1688 => x"fd8f1b25",
			1689 => x"01ad1b25",
			1690 => x"05079e10",
			1691 => x"040a6908",
			1692 => x"01011904",
			1693 => x"03051b25",
			1694 => x"fe881b25",
			1695 => x"07052f04",
			1696 => x"008f1b25",
			1697 => x"fe651b25",
			1698 => x"01014b08",
			1699 => x"00034b04",
			1700 => x"ffdc1b25",
			1701 => x"018b1b25",
			1702 => x"fe2e1b25",
			1703 => x"00039608",
			1704 => x"0f0a6e04",
			1705 => x"00801b25",
			1706 => x"fdfd1b25",
			1707 => x"0b072f10",
			1708 => x"040c6008",
			1709 => x"0100c304",
			1710 => x"01711b25",
			1711 => x"02211b25",
			1712 => x"0c056104",
			1713 => x"01eb1b25",
			1714 => x"fec41b25",
			1715 => x"06018e04",
			1716 => x"059d1b25",
			1717 => x"0f0b8804",
			1718 => x"fe891b25",
			1719 => x"01e21b25",
			1720 => x"01019020",
			1721 => x"0a02cc1c",
			1722 => x"01011f10",
			1723 => x"0d095608",
			1724 => x"040c6004",
			1725 => x"fe8a1b25",
			1726 => x"02fe1b25",
			1727 => x"0a029604",
			1728 => x"0ca71b25",
			1729 => x"02aa1b25",
			1730 => x"040ce108",
			1731 => x"0d097504",
			1732 => x"fe781b25",
			1733 => x"ffc31b25",
			1734 => x"02f21b25",
			1735 => x"fe5e1b25",
			1736 => x"01a11b25",
			1737 => x"0b05110c",
			1738 => x"02096c04",
			1739 => x"fe691c19",
			1740 => x"00052904",
			1741 => x"ff751c19",
			1742 => x"01141c19",
			1743 => x"0803e668",
			1744 => x"06018a34",
			1745 => x"0802aa18",
			1746 => x"0409db0c",
			1747 => x"0b06d208",
			1748 => x"0e094004",
			1749 => x"00f51c19",
			1750 => x"febe1c19",
			1751 => x"fe9f1c19",
			1752 => x"0c063008",
			1753 => x"0c05f204",
			1754 => x"00051c19",
			1755 => x"02311c19",
			1756 => x"ff3f1c19",
			1757 => x"0c04e90c",
			1758 => x"06016304",
			1759 => x"fe921c19",
			1760 => x"0f08cd04",
			1761 => x"00951c19",
			1762 => x"fe6c1c19",
			1763 => x"040ae208",
			1764 => x"08032804",
			1765 => x"00551c19",
			1766 => x"fe761c19",
			1767 => x"0901b804",
			1768 => x"ff6c1c19",
			1769 => x"fde51c19",
			1770 => x"0c052818",
			1771 => x"0c04cf08",
			1772 => x"05063204",
			1773 => x"fde11c19",
			1774 => x"00e41c19",
			1775 => x"09015a08",
			1776 => x"02096c04",
			1777 => x"00db1c19",
			1778 => x"01ed1c19",
			1779 => x"0c050c04",
			1780 => x"00001c19",
			1781 => x"01371c19",
			1782 => x"09014f0c",
			1783 => x"0100c304",
			1784 => x"fdd71c19",
			1785 => x"0100c804",
			1786 => x"01941c19",
			1787 => x"00001c19",
			1788 => x"0d086608",
			1789 => x"01011904",
			1790 => x"00381c19",
			1791 => x"01811c19",
			1792 => x"0f0aed04",
			1793 => x"ff3a1c19",
			1794 => x"008d1c19",
			1795 => x"0c04e704",
			1796 => x"01491c19",
			1797 => x"fe251c19",
			1798 => x"0601644c",
			1799 => x"09019624",
			1800 => x"0100930c",
			1801 => x"03069604",
			1802 => x"fe611dad",
			1803 => x"0306a504",
			1804 => x"01081dad",
			1805 => x"fe861dad",
			1806 => x"0900ec04",
			1807 => x"02731dad",
			1808 => x"0d07a310",
			1809 => x"0100dc08",
			1810 => x"0e070104",
			1811 => x"fe4e1dad",
			1812 => x"00031dad",
			1813 => x"0b060604",
			1814 => x"ff871dad",
			1815 => x"05891dad",
			1816 => x"fe661dad",
			1817 => x"07062b08",
			1818 => x"0d078804",
			1819 => x"01cc1dad",
			1820 => x"fe661dad",
			1821 => x"07064610",
			1822 => x"0e08cb04",
			1823 => x"fef71dad",
			1824 => x"01010204",
			1825 => x"ff411dad",
			1826 => x"08027904",
			1827 => x"05261dad",
			1828 => x"024b1dad",
			1829 => x"00032408",
			1830 => x"0b06cd04",
			1831 => x"015d1dad",
			1832 => x"fe7b1dad",
			1833 => x"0c063204",
			1834 => x"030e1dad",
			1835 => x"feac1dad",
			1836 => x"0c066c58",
			1837 => x"06019a34",
			1838 => x"0c04ea14",
			1839 => x"0b051108",
			1840 => x"040eab04",
			1841 => x"fe541dad",
			1842 => x"00c21dad",
			1843 => x"0100a808",
			1844 => x"0f088504",
			1845 => x"01971dad",
			1846 => x"001e1dad",
			1847 => x"020f1dad",
			1848 => x"08032910",
			1849 => x"0802fb08",
			1850 => x"0b06ee04",
			1851 => x"00ba1dad",
			1852 => x"ff2d1dad",
			1853 => x"06017404",
			1854 => x"ff5e1dad",
			1855 => x"01e81dad",
			1856 => x"07053108",
			1857 => x"0306e204",
			1858 => x"fee11dad",
			1859 => x"01891dad",
			1860 => x"0a02c304",
			1861 => x"fe121dad",
			1862 => x"ff951dad",
			1863 => x"0b072f14",
			1864 => x"040c7f0c",
			1865 => x"0308a904",
			1866 => x"01171dad",
			1867 => x"0a027b04",
			1868 => x"010b1dad",
			1869 => x"01f01dad",
			1870 => x"0c054604",
			1871 => x"01f91dad",
			1872 => x"fee71dad",
			1873 => x"0e0abb04",
			1874 => x"fe081dad",
			1875 => x"0c063a04",
			1876 => x"fece1dad",
			1877 => x"0601a604",
			1878 => x"feee1dad",
			1879 => x"02731dad",
			1880 => x"09026420",
			1881 => x"0a02ac1c",
			1882 => x"0d097510",
			1883 => x"0901bc08",
			1884 => x"0d092704",
			1885 => x"fef61dad",
			1886 => x"03451dad",
			1887 => x"0b07b504",
			1888 => x"fe991dad",
			1889 => x"ffa91dad",
			1890 => x"0802eb04",
			1891 => x"07821dad",
			1892 => x"0901fe04",
			1893 => x"032d1dad",
			1894 => x"fe911dad",
			1895 => x"fe651dad",
			1896 => x"0f0c3904",
			1897 => x"ff141dad",
			1898 => x"01cf1dad",
			1899 => x"040abb4c",
			1900 => x"0601793c",
			1901 => x"0c059e0c",
			1902 => x"0207a104",
			1903 => x"00001f59",
			1904 => x"0c04d104",
			1905 => x"00001f59",
			1906 => x"ff161f59",
			1907 => x"0c05f618",
			1908 => x"0e09330c",
			1909 => x"05075608",
			1910 => x"01010f04",
			1911 => x"00801f59",
			1912 => x"00001f59",
			1913 => x"ffb11f59",
			1914 => x"0507f508",
			1915 => x"0b06bc04",
			1916 => x"00001f59",
			1917 => x"009e1f59",
			1918 => x"00001f59",
			1919 => x"0e09330c",
			1920 => x"0f096004",
			1921 => x"ffed1f59",
			1922 => x"0f098b04",
			1923 => x"009b1f59",
			1924 => x"00001f59",
			1925 => x"0a021704",
			1926 => x"00001f59",
			1927 => x"01010b04",
			1928 => x"00001f59",
			1929 => x"ff4f1f59",
			1930 => x"0a024c04",
			1931 => x"00001f59",
			1932 => x"0e0a1b08",
			1933 => x"07068804",
			1934 => x"00fa1f59",
			1935 => x"00001f59",
			1936 => x"00001f59",
			1937 => x"040c1e44",
			1938 => x"06018a18",
			1939 => x"0704f10c",
			1940 => x"0d060f08",
			1941 => x"0b053304",
			1942 => x"ff8c1f59",
			1943 => x"00001f59",
			1944 => x"00cf1f59",
			1945 => x"0b075f08",
			1946 => x"0208e404",
			1947 => x"00001f59",
			1948 => x"ff3c1f59",
			1949 => x"00001f59",
			1950 => x"06018e10",
			1951 => x"0307c404",
			1952 => x"00001f59",
			1953 => x"040b2e04",
			1954 => x"00001f59",
			1955 => x"01015904",
			1956 => x"00d51f59",
			1957 => x"00001f59",
			1958 => x"0b071e10",
			1959 => x"01010208",
			1960 => x"0a02bc04",
			1961 => x"ff3a1f59",
			1962 => x"00001f59",
			1963 => x"0802f804",
			1964 => x"00001f59",
			1965 => x"01041f59",
			1966 => x"01015b08",
			1967 => x"08032804",
			1968 => x"fee21f59",
			1969 => x"00001f59",
			1970 => x"00001f59",
			1971 => x"0e08e128",
			1972 => x"01008618",
			1973 => x"0c04d10c",
			1974 => x"0505b004",
			1975 => x"00001f59",
			1976 => x"0b053504",
			1977 => x"01011f59",
			1978 => x"00001f59",
			1979 => x"040e6308",
			1980 => x"0704d404",
			1981 => x"00001f59",
			1982 => x"feee1f59",
			1983 => x"00001f59",
			1984 => x"0803e60c",
			1985 => x"06017804",
			1986 => x"00001f59",
			1987 => x"040fc604",
			1988 => x"010d1f59",
			1989 => x"00001f59",
			1990 => x"00001f59",
			1991 => x"0e0b770c",
			1992 => x"0d098508",
			1993 => x"0c061404",
			1994 => x"ffee1f59",
			1995 => x"fee21f59",
			1996 => x"00001f59",
			1997 => x"0d0a2b0c",
			1998 => x"01013b04",
			1999 => x"00001f59",
			2000 => x"01018304",
			2001 => x"00b71f59",
			2002 => x"00001f59",
			2003 => x"0c071e04",
			2004 => x"ffab1f59",
			2005 => x"00001f59",
			2006 => x"06015f28",
			2007 => x"01010214",
			2008 => x"08027910",
			2009 => x"0002f604",
			2010 => x"fe7520c5",
			2011 => x"0100e008",
			2012 => x"09006c04",
			2013 => x"000020c5",
			2014 => x"021f20c5",
			2015 => x"fef420c5",
			2016 => x"fe6520c5",
			2017 => x"03097810",
			2018 => x"0d083e0c",
			2019 => x"0901cc08",
			2020 => x"0b06ce04",
			2021 => x"fe9320c5",
			2022 => x"00a320c5",
			2023 => x"026e20c5",
			2024 => x"040320c5",
			2025 => x"fed120c5",
			2026 => x"05086a60",
			2027 => x"06018d34",
			2028 => x"040ac218",
			2029 => x"0100a108",
			2030 => x"0b055604",
			2031 => x"001220c5",
			2032 => x"fe1020c5",
			2033 => x"00037808",
			2034 => x"0a023904",
			2035 => x"013a20c5",
			2036 => x"ff7920c5",
			2037 => x"06017404",
			2038 => x"ffeb20c5",
			2039 => x"01a620c5",
			2040 => x"0b05560c",
			2041 => x"0b051104",
			2042 => x"fe6220c5",
			2043 => x"0704f104",
			2044 => x"015620c5",
			2045 => x"003620c5",
			2046 => x"08035e08",
			2047 => x"0a02b004",
			2048 => x"ff5f20c5",
			2049 => x"019c20c5",
			2050 => x"09014d04",
			2051 => x"fdef20c5",
			2052 => x"00d620c5",
			2053 => x"040c6018",
			2054 => x"00039108",
			2055 => x"0b070104",
			2056 => x"fdf920c5",
			2057 => x"01a420c5",
			2058 => x"07068608",
			2059 => x"0100c504",
			2060 => x"00ed20c5",
			2061 => x"01a220c5",
			2062 => x"0f0aed04",
			2063 => x"fe4020c5",
			2064 => x"01a420c5",
			2065 => x"0100a808",
			2066 => x"06019204",
			2067 => x"023220c5",
			2068 => x"012620c5",
			2069 => x"040dca08",
			2070 => x"0c061404",
			2071 => x"003920c5",
			2072 => x"fe4e20c5",
			2073 => x"fdda20c5",
			2074 => x"0004a02c",
			2075 => x"0d09691c",
			2076 => x"0901ce0c",
			2077 => x"0c068b08",
			2078 => x"0d092804",
			2079 => x"006120c5",
			2080 => x"01e420c5",
			2081 => x"ff0820c5",
			2082 => x"0d095008",
			2083 => x"0f0be504",
			2084 => x"fe8f20c5",
			2085 => x"016e20c5",
			2086 => x"0a026204",
			2087 => x"041b20c5",
			2088 => x"fec820c5",
			2089 => x"0003a204",
			2090 => x"033c20c5",
			2091 => x"0901d204",
			2092 => x"028420c5",
			2093 => x"0601ad04",
			2094 => x"fe8820c5",
			2095 => x"00a420c5",
			2096 => x"fe5320c5",
			2097 => x"0901db84",
			2098 => x"08033044",
			2099 => x"0a026524",
			2100 => x"0c05f810",
			2101 => x"0d08220c",
			2102 => x"0c054c04",
			2103 => x"ff6c2259",
			2104 => x"0100c004",
			2105 => x"00ed2259",
			2106 => x"ffe32259",
			2107 => x"febd2259",
			2108 => x"00035b0c",
			2109 => x"07065a04",
			2110 => x"ff7d2259",
			2111 => x"0c063004",
			2112 => x"00752259",
			2113 => x"ff9f2259",
			2114 => x"03097804",
			2115 => x"00ef2259",
			2116 => x"00002259",
			2117 => x"040aa10c",
			2118 => x"0b057408",
			2119 => x"01009f04",
			2120 => x"00002259",
			2121 => x"00d72259",
			2122 => x"ff8e2259",
			2123 => x"030a690c",
			2124 => x"0704ec04",
			2125 => x"00002259",
			2126 => x"0c04b104",
			2127 => x"00002259",
			2128 => x"fe4b2259",
			2129 => x"0e0a7604",
			2130 => x"00142259",
			2131 => x"00002259",
			2132 => x"0100c324",
			2133 => x"0c052a20",
			2134 => x"03067810",
			2135 => x"0704ef08",
			2136 => x"06017404",
			2137 => x"ffb22259",
			2138 => x"00db2259",
			2139 => x"040e6304",
			2140 => x"fecc2259",
			2141 => x"00002259",
			2142 => x"0e064308",
			2143 => x"07051a04",
			2144 => x"01392259",
			2145 => x"00002259",
			2146 => x"03071b04",
			2147 => x"ffbd2259",
			2148 => x"003c2259",
			2149 => x"fea62259",
			2150 => x"0507480c",
			2151 => x"040da908",
			2152 => x"06018d04",
			2153 => x"00002259",
			2154 => x"01942259",
			2155 => x"00002259",
			2156 => x"0507f504",
			2157 => x"fef12259",
			2158 => x"040cb604",
			2159 => x"00002259",
			2160 => x"0a02cc04",
			2161 => x"011f2259",
			2162 => x"00002259",
			2163 => x"0901fe24",
			2164 => x"0e092404",
			2165 => x"ff6c2259",
			2166 => x"040c5818",
			2167 => x"0003680c",
			2168 => x"0a023908",
			2169 => x"07065c04",
			2170 => x"00862259",
			2171 => x"00002259",
			2172 => x"ff952259",
			2173 => x"0a024c04",
			2174 => x"00002259",
			2175 => x"07066d04",
			2176 => x"014b2259",
			2177 => x"00132259",
			2178 => x"0a02a904",
			2179 => x"00002259",
			2180 => x"ff772259",
			2181 => x"0e0c7e20",
			2182 => x"0b07c31c",
			2183 => x"0101450c",
			2184 => x"0e0aee08",
			2185 => x"0d084a04",
			2186 => x"00002259",
			2187 => x"ff262259",
			2188 => x"00002259",
			2189 => x"01014908",
			2190 => x"0802dd04",
			2191 => x"00002259",
			2192 => x"01142259",
			2193 => x"0b07b504",
			2194 => x"ffcb2259",
			2195 => x"00c72259",
			2196 => x"fea72259",
			2197 => x"00bb2259",
			2198 => x"0802791c",
			2199 => x"07065b18",
			2200 => x"0c056204",
			2201 => x"000023c5",
			2202 => x"0b06df10",
			2203 => x"08021e04",
			2204 => x"000023c5",
			2205 => x"0d084c08",
			2206 => x"0507f504",
			2207 => x"00f223c5",
			2208 => x"000023c5",
			2209 => x"000023c5",
			2210 => x"000023c5",
			2211 => x"000023c5",
			2212 => x"00042850",
			2213 => x"0100a624",
			2214 => x"07051b18",
			2215 => x"0505f610",
			2216 => x"0b053508",
			2217 => x"040b7804",
			2218 => x"ff3723c5",
			2219 => x"000023c5",
			2220 => x"07050804",
			2221 => x"005523c5",
			2222 => x"000023c5",
			2223 => x"0c04b904",
			2224 => x"000023c5",
			2225 => x"fea223c5",
			2226 => x"0c04d204",
			2227 => x"005a23c5",
			2228 => x"0f083904",
			2229 => x"000023c5",
			2230 => x"ffc023c5",
			2231 => x"0d06d410",
			2232 => x"0f090d0c",
			2233 => x"0100a804",
			2234 => x"000023c5",
			2235 => x"0003b704",
			2236 => x"000023c5",
			2237 => x"012323c5",
			2238 => x"000023c5",
			2239 => x"0100e50c",
			2240 => x"0100be04",
			2241 => x"000023c5",
			2242 => x"0b05d604",
			2243 => x"000023c5",
			2244 => x"fe9f23c5",
			2245 => x"09019c08",
			2246 => x"0003d904",
			2247 => x"00ef23c5",
			2248 => x"000023c5",
			2249 => x"0a027004",
			2250 => x"ffca23c5",
			2251 => x"003223c5",
			2252 => x"0c052a28",
			2253 => x"03071b1c",
			2254 => x"0209000c",
			2255 => x"03067808",
			2256 => x"040c2c04",
			2257 => x"ff5623c5",
			2258 => x"000023c5",
			2259 => x"015323c5",
			2260 => x"00043d08",
			2261 => x"00043204",
			2262 => x"000023c5",
			2263 => x"fecf23c5",
			2264 => x"0306b904",
			2265 => x"ffd023c5",
			2266 => x"009623c5",
			2267 => x"0f09e108",
			2268 => x"08035204",
			2269 => x"000023c5",
			2270 => x"015123c5",
			2271 => x"000023c5",
			2272 => x"0004350c",
			2273 => x"0c067008",
			2274 => x"08034404",
			2275 => x"000023c5",
			2276 => x"00d823c5",
			2277 => x"000023c5",
			2278 => x"030d4e10",
			2279 => x"08036908",
			2280 => x"08036504",
			2281 => x"ffc023c5",
			2282 => x"003823c5",
			2283 => x"040ceb04",
			2284 => x"000023c5",
			2285 => x"febf23c5",
			2286 => x"08047204",
			2287 => x"008823c5",
			2288 => x"000023c5",
			2289 => x"0505af08",
			2290 => x"0804ac04",
			2291 => x"fed824d9",
			2292 => x"000024d9",
			2293 => x"0c04ca18",
			2294 => x"040bb208",
			2295 => x"0900fe04",
			2296 => x"ff2124d9",
			2297 => x"006124d9",
			2298 => x"0505b004",
			2299 => x"000024d9",
			2300 => x"06016c08",
			2301 => x"06016304",
			2302 => x"000024d9",
			2303 => x"001524d9",
			2304 => x"018a24d9",
			2305 => x"03090738",
			2306 => x"08034120",
			2307 => x"040a5b10",
			2308 => x"06017408",
			2309 => x"0c054c04",
			2310 => x"ff3724d9",
			2311 => x"002324d9",
			2312 => x"02092404",
			2313 => x"00bc24d9",
			2314 => x"000024d9",
			2315 => x"0f084608",
			2316 => x"07050804",
			2317 => x"007e24d9",
			2318 => x"ff4524d9",
			2319 => x"0c04ce04",
			2320 => x"000024d9",
			2321 => x"fe8a24d9",
			2322 => x"0c04cd0c",
			2323 => x"08035b04",
			2324 => x"000024d9",
			2325 => x"03064804",
			2326 => x"000024d9",
			2327 => x"fe7a24d9",
			2328 => x"0c052a08",
			2329 => x"03066904",
			2330 => x"ff8b24d9",
			2331 => x"005c24d9",
			2332 => x"fed024d9",
			2333 => x"05080414",
			2334 => x"0803a010",
			2335 => x"020a4608",
			2336 => x"0901fc04",
			2337 => x"009224d9",
			2338 => x"ff8e24d9",
			2339 => x"0f0a4204",
			2340 => x"000024d9",
			2341 => x"015d24d9",
			2342 => x"ffbd24d9",
			2343 => x"05083010",
			2344 => x"01014108",
			2345 => x"030a9904",
			2346 => x"fe1b24d9",
			2347 => x"000024d9",
			2348 => x"05081304",
			2349 => x"008324d9",
			2350 => x"000024d9",
			2351 => x"0c06c708",
			2352 => x"040ce104",
			2353 => x"001024d9",
			2354 => x"00f624d9",
			2355 => x"0509e304",
			2356 => x"feb624d9",
			2357 => x"000024d9",
			2358 => x"0d05b608",
			2359 => x"0209ab04",
			2360 => x"fe972605",
			2361 => x"00002605",
			2362 => x"0f083948",
			2363 => x"0306b930",
			2364 => x"040c0414",
			2365 => x"0704d808",
			2366 => x"0b053304",
			2367 => x"ffa12605",
			2368 => x"00592605",
			2369 => x"0f07eb08",
			2370 => x"0d060304",
			2371 => x"ff442605",
			2372 => x"000c2605",
			2373 => x"fe7a2605",
			2374 => x"02091b0c",
			2375 => x"06016304",
			2376 => x"00002605",
			2377 => x"0c04ef04",
			2378 => x"01862605",
			2379 => x"00002605",
			2380 => x"06018008",
			2381 => x"0704ec04",
			2382 => x"00002605",
			2383 => x"fe922605",
			2384 => x"0c04f104",
			2385 => x"01082605",
			2386 => x"ff502605",
			2387 => x"0a026210",
			2388 => x"0208090c",
			2389 => x"0705a504",
			2390 => x"00002605",
			2391 => x"0b060b04",
			2392 => x"00d02605",
			2393 => x"00002605",
			2394 => x"ff342605",
			2395 => x"040df504",
			2396 => x"01922605",
			2397 => x"00002605",
			2398 => x"0306e20c",
			2399 => x"06017c04",
			2400 => x"fdf42605",
			2401 => x"0f087204",
			2402 => x"01332605",
			2403 => x"00002605",
			2404 => x"0c064d20",
			2405 => x"0b072010",
			2406 => x"06019608",
			2407 => x"02096604",
			2408 => x"00462605",
			2409 => x"ff9c2605",
			2410 => x"040d0e04",
			2411 => x"01682605",
			2412 => x"ff502605",
			2413 => x"0d08b308",
			2414 => x"0901fa04",
			2415 => x"fc582605",
			2416 => x"00002605",
			2417 => x"0d090104",
			2418 => x"00932605",
			2419 => x"fea72605",
			2420 => x"0601af0c",
			2421 => x"040ab204",
			2422 => x"ff252605",
			2423 => x"01015004",
			2424 => x"011e2605",
			2425 => x"00292605",
			2426 => x"0e0c7e08",
			2427 => x"0b087804",
			2428 => x"fea22605",
			2429 => x"00002605",
			2430 => x"0d0a1e04",
			2431 => x"01022605",
			2432 => x"00002605",
			2433 => x"06017460",
			2434 => x"0f09b154",
			2435 => x"06016724",
			2436 => x"0901a114",
			2437 => x"0601640c",
			2438 => x"01009304",
			2439 => x"d16e27c1",
			2440 => x"0900ec04",
			2441 => x"d51f27c1",
			2442 => x"d18427c1",
			2443 => x"0306a504",
			2444 => x"d19d27c1",
			2445 => x"d32227c1",
			2446 => x"0a02170c",
			2447 => x"0b06dd08",
			2448 => x"02092e04",
			2449 => x"d34827c1",
			2450 => x"e36827c1",
			2451 => x"d19727c1",
			2452 => x"d17627c1",
			2453 => x"0c04d218",
			2454 => x"0d06030c",
			2455 => x"0505cc04",
			2456 => x"d17a27c1",
			2457 => x"01007e04",
			2458 => x"dba727c1",
			2459 => x"d1b827c1",
			2460 => x"02091b08",
			2461 => x"0306b904",
			2462 => x"e0d227c1",
			2463 => x"eb5d27c1",
			2464 => x"d1a927c1",
			2465 => x"0a022308",
			2466 => x"0c05f604",
			2467 => x"d91127c1",
			2468 => x"d1d427c1",
			2469 => x"0c061108",
			2470 => x"02083004",
			2471 => x"d3b027c1",
			2472 => x"d19527c1",
			2473 => x"03096804",
			2474 => x"d86c27c1",
			2475 => x"d19627c1",
			2476 => x"0c05f504",
			2477 => x"de1927c1",
			2478 => x"040a4904",
			2479 => x"d18427c1",
			2480 => x"d7e127c1",
			2481 => x"0c063a54",
			2482 => x"0601852c",
			2483 => x"02095d18",
			2484 => x"0c05070c",
			2485 => x"0505af04",
			2486 => x"d3b027c1",
			2487 => x"06017504",
			2488 => x"e51027c1",
			2489 => x"eb7027c1",
			2490 => x"0100a808",
			2491 => x"01009b04",
			2492 => x"d3e527c1",
			2493 => x"d1d427c1",
			2494 => x"d91127c1",
			2495 => x"0b055604",
			2496 => x"dc3f27c1",
			2497 => x"0f0a0308",
			2498 => x"040a5b04",
			2499 => x"d2f527c1",
			2500 => x"d17e27c1",
			2501 => x"0802d704",
			2502 => x"d32227c1",
			2503 => x"e5fe27c1",
			2504 => x"05083e1c",
			2505 => x"0802e30c",
			2506 => x"0b06dd04",
			2507 => x"e20427c1",
			2508 => x"0d085b04",
			2509 => x"d67b27c1",
			2510 => x"d1ac27c1",
			2511 => x"040d0e08",
			2512 => x"06018d04",
			2513 => x"e6e927c1",
			2514 => x"ecbe27c1",
			2515 => x"0c052e04",
			2516 => x"e61827c1",
			2517 => x"d2bc27c1",
			2518 => x"020b5b08",
			2519 => x"06019904",
			2520 => x"d76a27c1",
			2521 => x"d1b427c1",
			2522 => x"df8527c1",
			2523 => x"0c065210",
			2524 => x"0601a60c",
			2525 => x"06018a08",
			2526 => x"01014b04",
			2527 => x"d91127c1",
			2528 => x"d1b827c1",
			2529 => x"d18327c1",
			2530 => x"e14a27c1",
			2531 => x"09026b14",
			2532 => x"0d08b304",
			2533 => x"d7e127c1",
			2534 => x"06017d08",
			2535 => x"01014e04",
			2536 => x"d67b27c1",
			2537 => x"d1d427c1",
			2538 => x"0b076304",
			2539 => x"d2e027c1",
			2540 => x"d18227c1",
			2541 => x"030c2504",
			2542 => x"d1b827c1",
			2543 => x"de3c27c1",
			2544 => x"020ad1a0",
			2545 => x"02095140",
			2546 => x"03065914",
			2547 => x"0a02ed08",
			2548 => x"0100a104",
			2549 => x"fecf2985",
			2550 => x"00002985",
			2551 => x"0803e608",
			2552 => x"0505af04",
			2553 => x"00002985",
			2554 => x"00c92985",
			2555 => x"ff8b2985",
			2556 => x"0003ea18",
			2557 => x"0100a608",
			2558 => x"0208b904",
			2559 => x"00002985",
			2560 => x"fe612985",
			2561 => x"0506a608",
			2562 => x"0100b404",
			2563 => x"00002985",
			2564 => x"00f52985",
			2565 => x"0c05f204",
			2566 => x"ff1d2985",
			2567 => x"00302985",
			2568 => x"0e070110",
			2569 => x"02091108",
			2570 => x"0c04f104",
			2571 => x"00fc2985",
			2572 => x"fedf2985",
			2573 => x"06017c04",
			2574 => x"ff182985",
			2575 => x"00c12985",
			2576 => x"017f2985",
			2577 => x"01012838",
			2578 => x"00043f1c",
			2579 => x"040b3610",
			2580 => x"0209b108",
			2581 => x"05065d04",
			2582 => x"00002985",
			2583 => x"fefb2985",
			2584 => x"0e09e004",
			2585 => x"00a72985",
			2586 => x"ff812985",
			2587 => x"0b057404",
			2588 => x"00002985",
			2589 => x"0a02bc04",
			2590 => x"fe312985",
			2591 => x"00002985",
			2592 => x"0601830c",
			2593 => x"02096608",
			2594 => x"0c04cf04",
			2595 => x"00892985",
			2596 => x"ffc22985",
			2597 => x"fe952985",
			2598 => x"07054b08",
			2599 => x"02097004",
			2600 => x"00002985",
			2601 => x"01632985",
			2602 => x"03087504",
			2603 => x"fe9d2985",
			2604 => x"00a42985",
			2605 => x"0c05d80c",
			2606 => x"0e092404",
			2607 => x"00002985",
			2608 => x"01014704",
			2609 => x"01422985",
			2610 => x"00002985",
			2611 => x"0003920c",
			2612 => x"0e0a1b08",
			2613 => x"0802d404",
			2614 => x"ff862985",
			2615 => x"00402985",
			2616 => x"ff022985",
			2617 => x"0b071008",
			2618 => x"0802e304",
			2619 => x"00002985",
			2620 => x"011c2985",
			2621 => x"0b075f04",
			2622 => x"ff302985",
			2623 => x"00b32985",
			2624 => x"0a02d12c",
			2625 => x"0b071008",
			2626 => x"0507ab04",
			2627 => x"00002985",
			2628 => x"014c2985",
			2629 => x"040cc61c",
			2630 => x"0b07b510",
			2631 => x"05086a08",
			2632 => x"020b1f04",
			2633 => x"ffb62985",
			2634 => x"007b2985",
			2635 => x"07072204",
			2636 => x"fec62985",
			2637 => x"00002985",
			2638 => x"08031e08",
			2639 => x"030b2a04",
			2640 => x"00002985",
			2641 => x"00e72985",
			2642 => x"00002985",
			2643 => x"00043504",
			2644 => x"01332985",
			2645 => x"00002985",
			2646 => x"0a02dd04",
			2647 => x"febe2985",
			2648 => x"0c06cb10",
			2649 => x"05083e08",
			2650 => x"0b065b04",
			2651 => x"00752985",
			2652 => x"fef62985",
			2653 => x"01014704",
			2654 => x"00002985",
			2655 => x"014e2985",
			2656 => x"ff202985",
			2657 => x"03061110",
			2658 => x"06017404",
			2659 => x"fe662afb",
			2660 => x"040f0204",
			2661 => x"ff772afb",
			2662 => x"0209d404",
			2663 => x"021e2afb",
			2664 => x"ff082afb",
			2665 => x"06018a60",
			2666 => x"0c04e924",
			2667 => x"06016304",
			2668 => x"fe862afb",
			2669 => x"02091110",
			2670 => x"0208bb08",
			2671 => x"0e064304",
			2672 => x"01c92afb",
			2673 => x"fe802afb",
			2674 => x"0505cc04",
			2675 => x"ffc22afb",
			2676 => x"01ec2afb",
			2677 => x"06017908",
			2678 => x"0b054504",
			2679 => x"ffc62afb",
			2680 => x"fcce2afb",
			2681 => x"01009504",
			2682 => x"00422afb",
			2683 => x"01c12afb",
			2684 => x"040a691c",
			2685 => x"06014a0c",
			2686 => x"0900fb08",
			2687 => x"0c052804",
			2688 => x"ffcc2afb",
			2689 => x"01492afb",
			2690 => x"fe7f2afb",
			2691 => x"06016208",
			2692 => x"0c05f804",
			2693 => x"00c52afb",
			2694 => x"02622afb",
			2695 => x"00035304",
			2696 => x"ffa82afb",
			2697 => x"013b2afb",
			2698 => x"0b056310",
			2699 => x"0306c508",
			2700 => x"0f082b04",
			2701 => x"ffc02afb",
			2702 => x"fdd52afb",
			2703 => x"0f088e04",
			2704 => x"01f82afb",
			2705 => x"ffaa2afb",
			2706 => x"0e098708",
			2707 => x"0c04f104",
			2708 => x"ffa52afb",
			2709 => x"fe862afb",
			2710 => x"05081f04",
			2711 => x"00822afb",
			2712 => x"fece2afb",
			2713 => x"05080418",
			2714 => x"040d2e0c",
			2715 => x"0e089608",
			2716 => x"0b05a704",
			2717 => x"01b72afb",
			2718 => x"ff1b2afb",
			2719 => x"01a82afb",
			2720 => x"09010204",
			2721 => x"01ca2afb",
			2722 => x"040dca04",
			2723 => x"00272afb",
			2724 => x"fe102afb",
			2725 => x"0f0ad918",
			2726 => x"09022810",
			2727 => x"0f0ac908",
			2728 => x"01015804",
			2729 => x"fe232afb",
			2730 => x"00002afb",
			2731 => x"0b076304",
			2732 => x"00002afb",
			2733 => x"ff7f2afb",
			2734 => x"030aa904",
			2735 => x"02a12afb",
			2736 => x"fec32afb",
			2737 => x"0802e910",
			2738 => x"0b078208",
			2739 => x"09022d04",
			2740 => x"1d7a2afb",
			2741 => x"00002afb",
			2742 => x"030b2a04",
			2743 => x"feb82afb",
			2744 => x"067e2afb",
			2745 => x"0004a008",
			2746 => x"01015504",
			2747 => x"01162afb",
			2748 => x"ffea2afb",
			2749 => x"fe652afb",
			2750 => x"03063a20",
			2751 => x"040e6308",
			2752 => x"0d066b04",
			2753 => x"fe752bcd",
			2754 => x"00002bcd",
			2755 => x"0e050010",
			2756 => x"0209ab04",
			2757 => x"fea82bcd",
			2758 => x"0209b108",
			2759 => x"0a03bd04",
			2760 => x"00a82bcd",
			2761 => x"00002bcd",
			2762 => x"00002bcd",
			2763 => x"0505f904",
			2764 => x"011c2bcd",
			2765 => x"00002bcd",
			2766 => x"0208e428",
			2767 => x"01007d08",
			2768 => x"0e060f04",
			2769 => x"02572bcd",
			2770 => x"00002bcd",
			2771 => x"0306b90c",
			2772 => x"00042804",
			2773 => x"fe7f2bcd",
			2774 => x"03066904",
			2775 => x"fe9d2bcd",
			2776 => x"00ef2bcd",
			2777 => x"0003ea10",
			2778 => x"0100a808",
			2779 => x"0c04d204",
			2780 => x"003a2bcd",
			2781 => x"fde42bcd",
			2782 => x"04091d04",
			2783 => x"00002bcd",
			2784 => x"01772bcd",
			2785 => x"02182bcd",
			2786 => x"0505db08",
			2787 => x"02090904",
			2788 => x"003a2bcd",
			2789 => x"fe672bcd",
			2790 => x"0803e618",
			2791 => x"0505f90c",
			2792 => x"00042004",
			2793 => x"feca2bcd",
			2794 => x"06017004",
			2795 => x"00492bcd",
			2796 => x"01bf2bcd",
			2797 => x"0d061d04",
			2798 => x"fdb92bcd",
			2799 => x"040bb004",
			2800 => x"004f2bcd",
			2801 => x"ffb42bcd",
			2802 => x"fe412bcd",
			2803 => x"03063a20",
			2804 => x"06017008",
			2805 => x"01009f04",
			2806 => x"fe6c2cd1",
			2807 => x"00002cd1",
			2808 => x"0900c610",
			2809 => x"0505a004",
			2810 => x"ff622cd1",
			2811 => x"0f07b908",
			2812 => x"0005fa04",
			2813 => x"01942cd1",
			2814 => x"00002cd1",
			2815 => x"00002cd1",
			2816 => x"01008204",
			2817 => x"fdd22cd1",
			2818 => x"00002cd1",
			2819 => x"0f081620",
			2820 => x"08035310",
			2821 => x"0306a504",
			2822 => x"fe852cd1",
			2823 => x"0f07fe08",
			2824 => x"0f07d504",
			2825 => x"ff932cd1",
			2826 => x"02472cd1",
			2827 => x"ff842cd1",
			2828 => x"03065908",
			2829 => x"01007d04",
			2830 => x"01b52cd1",
			2831 => x"fe672cd1",
			2832 => x"0b055604",
			2833 => x"01f92cd1",
			2834 => x"00002cd1",
			2835 => x"0306ff20",
			2836 => x"0b055414",
			2837 => x"0f088b10",
			2838 => x"06017008",
			2839 => x"0b053304",
			2840 => x"fffc2cd1",
			2841 => x"fe782cd1",
			2842 => x"0306c504",
			2843 => x"00002cd1",
			2844 => x"01b02cd1",
			2845 => x"fdba2cd1",
			2846 => x"02091b04",
			2847 => x"fbfa2cd1",
			2848 => x"06017c04",
			2849 => x"fea02cd1",
			2850 => x"00002cd1",
			2851 => x"01009508",
			2852 => x"00046704",
			2853 => x"fd912cd1",
			2854 => x"00f22cd1",
			2855 => x"0506160c",
			2856 => x"0f08bf08",
			2857 => x"0505f904",
			2858 => x"00982cd1",
			2859 => x"01ae2cd1",
			2860 => x"00002cd1",
			2861 => x"0100f508",
			2862 => x"06018104",
			2863 => x"ff1e2cd1",
			2864 => x"004d2cd1",
			2865 => x"040b8a04",
			2866 => x"008d2cd1",
			2867 => x"ffc72cd1",
			2868 => x"07050434",
			2869 => x"0f083920",
			2870 => x"0306b91c",
			2871 => x"040c5808",
			2872 => x"03069604",
			2873 => x"fec42dcd",
			2874 => x"00002dcd",
			2875 => x"0b051408",
			2876 => x"0305b004",
			2877 => x"ff772dcd",
			2878 => x"00002dcd",
			2879 => x"0f081608",
			2880 => x"06016304",
			2881 => x"00002dcd",
			2882 => x"013c2dcd",
			2883 => x"ffbf2dcd",
			2884 => x"01412dcd",
			2885 => x"03071b10",
			2886 => x"0e06ac0c",
			2887 => x"01008608",
			2888 => x"040cc604",
			2889 => x"ff9e2dcd",
			2890 => x"00002dcd",
			2891 => x"00212dcd",
			2892 => x"fe582dcd",
			2893 => x"00fd2dcd",
			2894 => x"07050810",
			2895 => x"03066908",
			2896 => x"0c04b904",
			2897 => x"00002dcd",
			2898 => x"ff892dcd",
			2899 => x"08032004",
			2900 => x"00002dcd",
			2901 => x"015f2dcd",
			2902 => x"0d061d08",
			2903 => x"040e6304",
			2904 => x"febb2dcd",
			2905 => x"00002dcd",
			2906 => x"05061914",
			2907 => x"06017408",
			2908 => x"0c04d404",
			2909 => x"00002dcd",
			2910 => x"ff2f2dcd",
			2911 => x"00042008",
			2912 => x"0f088b04",
			2913 => x"00e22dcd",
			2914 => x"ffa72dcd",
			2915 => x"01912dcd",
			2916 => x"0c05bb10",
			2917 => x"0a02a808",
			2918 => x"040adc04",
			2919 => x"00002dcd",
			2920 => x"fe8a2dcd",
			2921 => x"07054504",
			2922 => x"00d02dcd",
			2923 => x"ffa52dcd",
			2924 => x"040bff08",
			2925 => x"0802fb04",
			2926 => x"001b2dcd",
			2927 => x"00db2dcd",
			2928 => x"0f0b2d04",
			2929 => x"ff102dcd",
			2930 => x"003d2dcd",
			2931 => x"0b05140c",
			2932 => x"040eab04",
			2933 => x"fea92e89",
			2934 => x"00053e04",
			2935 => x"00002e89",
			2936 => x"ffde2e89",
			2937 => x"0704f110",
			2938 => x"06016704",
			2939 => x"fff12e89",
			2940 => x"0704ea08",
			2941 => x"0704d704",
			2942 => x"00732e89",
			2943 => x"00002e89",
			2944 => x"01542e89",
			2945 => x"07050108",
			2946 => x"040ad504",
			2947 => x"00002e89",
			2948 => x"fe112e89",
			2949 => x"0d08661c",
			2950 => x"0e09fd10",
			2951 => x"0a02a908",
			2952 => x"040ae204",
			2953 => x"00232e89",
			2954 => x"fef32e89",
			2955 => x"0900e904",
			2956 => x"ffba2e89",
			2957 => x"00b42e89",
			2958 => x"05081208",
			2959 => x"01012504",
			2960 => x"00002e89",
			2961 => x"01532e89",
			2962 => x"00002e89",
			2963 => x"05083010",
			2964 => x"0d088d08",
			2965 => x"0e0a6d04",
			2966 => x"ff102e89",
			2967 => x"00842e89",
			2968 => x"030ac504",
			2969 => x"fd392e89",
			2970 => x"00002e89",
			2971 => x"0802ee08",
			2972 => x"07070c04",
			2973 => x"00982e89",
			2974 => x"00002e89",
			2975 => x"0b072004",
			2976 => x"00ca2e89",
			2977 => x"ffa22e89",
			2978 => x"0505cc14",
			2979 => x"040d6e08",
			2980 => x"03066904",
			2981 => x"fe6c2f9d",
			2982 => x"00002f9d",
			2983 => x"0b051108",
			2984 => x"03059904",
			2985 => x"ff572f9d",
			2986 => x"00002f9d",
			2987 => x"00e42f9d",
			2988 => x"0f082234",
			2989 => x"07050818",
			2990 => x"0a02a60c",
			2991 => x"0c04d104",
			2992 => x"fea92f9d",
			2993 => x"0c04d204",
			2994 => x"01322f9d",
			2995 => x"00002f9d",
			2996 => x"03063204",
			2997 => x"00002f9d",
			2998 => x"0c04d404",
			2999 => x"01ac2f9d",
			3000 => x"009b2f9d",
			3001 => x"0e06e214",
			3002 => x"0f07e308",
			3003 => x"00037d04",
			3004 => x"00002f9d",
			3005 => x"fe622f9d",
			3006 => x"0a02bb04",
			3007 => x"ff252f9d",
			3008 => x"0c050704",
			3009 => x"00c52f9d",
			3010 => x"00002f9d",
			3011 => x"06011d04",
			3012 => x"00002f9d",
			3013 => x"01332f9d",
			3014 => x"09011b28",
			3015 => x"0e072518",
			3016 => x"0306c508",
			3017 => x"06017d04",
			3018 => x"fe2f2f9d",
			3019 => x"00002f9d",
			3020 => x"0d065108",
			3021 => x"0f088504",
			3022 => x"00cf2f9d",
			3023 => x"ff732f9d",
			3024 => x"03073b04",
			3025 => x"fe5c2f9d",
			3026 => x"008b2f9d",
			3027 => x"03076c04",
			3028 => x"fded2f9d",
			3029 => x"0b059304",
			3030 => x"00e22f9d",
			3031 => x"06018904",
			3032 => x"00342f9d",
			3033 => x"fe922f9d",
			3034 => x"05066c08",
			3035 => x"0003c004",
			3036 => x"00002f9d",
			3037 => x"01912f9d",
			3038 => x"0307f404",
			3039 => x"fe622f9d",
			3040 => x"0d09f808",
			3041 => x"0f0aed04",
			3042 => x"ffda2f9d",
			3043 => x"00812f9d",
			3044 => x"0e0d6804",
			3045 => x"fe6a2f9d",
			3046 => x"00002f9d",
			3047 => x"0505db24",
			3048 => x"040c930c",
			3049 => x"07050804",
			3050 => x"fe5c30b9",
			3051 => x"07051804",
			3052 => x"000030b9",
			3053 => x"ff7a30b9",
			3054 => x"0d05a804",
			3055 => x"fe9e30b9",
			3056 => x"0f080e10",
			3057 => x"0601700c",
			3058 => x"0a02c408",
			3059 => x"0a02bf04",
			3060 => x"000030b9",
			3061 => x"006530b9",
			3062 => x"ffdf30b9",
			3063 => x"016f30b9",
			3064 => x"fee730b9",
			3065 => x"0505f620",
			3066 => x"0d060f14",
			3067 => x"0b053308",
			3068 => x"0900d304",
			3069 => x"000030b9",
			3070 => x"fe8330b9",
			3071 => x"07050408",
			3072 => x"06016404",
			3073 => x"000030b9",
			3074 => x"018b30b9",
			3075 => x"ffd430b9",
			3076 => x"06016304",
			3077 => x"000030b9",
			3078 => x"07051c04",
			3079 => x"01a830b9",
			3080 => x"000030b9",
			3081 => x"0d061f18",
			3082 => x"040cc610",
			3083 => x"0f08460c",
			3084 => x"07050104",
			3085 => x"002f30b9",
			3086 => x"01008004",
			3087 => x"000030b9",
			3088 => x"fe1b30b9",
			3089 => x"fdac30b9",
			3090 => x"0b055604",
			3091 => x"00c330b9",
			3092 => x"000030b9",
			3093 => x"0b055614",
			3094 => x"00043f10",
			3095 => x"0d062b08",
			3096 => x"01009004",
			3097 => x"003c30b9",
			3098 => x"fe6530b9",
			3099 => x"0b055404",
			3100 => x"002d30b9",
			3101 => x"01c230b9",
			3102 => x"01de30b9",
			3103 => x"0e06ce10",
			3104 => x"00037d08",
			3105 => x"07059104",
			3106 => x"000030b9",
			3107 => x"002230b9",
			3108 => x"06018104",
			3109 => x"fde230b9",
			3110 => x"000030b9",
			3111 => x"07051f08",
			3112 => x"0100a304",
			3113 => x"000030b9",
			3114 => x"018b30b9",
			3115 => x"09014b04",
			3116 => x"ff0430b9",
			3117 => x"003530b9",
			3118 => x"00042834",
			3119 => x"01009308",
			3120 => x"040b7604",
			3121 => x"fe7031dd",
			3122 => x"000031dd",
			3123 => x"00042428",
			3124 => x"0c04d108",
			3125 => x"06017004",
			3126 => x"000031dd",
			3127 => x"012931dd",
			3128 => x"0705a410",
			3129 => x"0208f008",
			3130 => x"040ac204",
			3131 => x"000031dd",
			3132 => x"008631dd",
			3133 => x"06019604",
			3134 => x"ff0031dd",
			3135 => x"000031dd",
			3136 => x"08033408",
			3137 => x"0d087204",
			3138 => x"003031dd",
			3139 => x"ffb731dd",
			3140 => x"0c065004",
			3141 => x"012a31dd",
			3142 => x"000031dd",
			3143 => x"feed31dd",
			3144 => x"0c052a3c",
			3145 => x"0601741c",
			3146 => x"02090010",
			3147 => x"0e05e908",
			3148 => x"0e05ce04",
			3149 => x"ff7931dd",
			3150 => x"000031dd",
			3151 => x"0a02a504",
			3152 => x"000031dd",
			3153 => x"014431dd",
			3154 => x"040d5508",
			3155 => x"0704d504",
			3156 => x"000031dd",
			3157 => x"feb531dd",
			3158 => x"000031dd",
			3159 => x"0a032118",
			3160 => x"06018510",
			3161 => x"02095d08",
			3162 => x"040b8504",
			3163 => x"000031dd",
			3164 => x"00bb31dd",
			3165 => x"0f089504",
			3166 => x"000031dd",
			3167 => x"ff6c31dd",
			3168 => x"00043204",
			3169 => x"000031dd",
			3170 => x"017031dd",
			3171 => x"0a035404",
			3172 => x"ff5a31dd",
			3173 => x"000031dd",
			3174 => x"0004350c",
			3175 => x"0c067008",
			3176 => x"06019a04",
			3177 => x"000031dd",
			3178 => x"00c731dd",
			3179 => x"000031dd",
			3180 => x"0e0c7e10",
			3181 => x"040d2e0c",
			3182 => x"08038208",
			3183 => x"08036904",
			3184 => x"000031dd",
			3185 => x"ff0e31dd",
			3186 => x"002731dd",
			3187 => x"fea031dd",
			3188 => x"07075204",
			3189 => x"00b431dd",
			3190 => x"fffa31dd",
			3191 => x"03063a14",
			3192 => x"06017008",
			3193 => x"01009f04",
			3194 => x"fe6d32b1",
			3195 => x"000032b1",
			3196 => x"07051808",
			3197 => x"0b050404",
			3198 => x"ff5832b1",
			3199 => x"016d32b1",
			3200 => x"fdb632b1",
			3201 => x"00050854",
			3202 => x"00042524",
			3203 => x"0306b908",
			3204 => x"00041c04",
			3205 => x"fe6532b1",
			3206 => x"fbba32b1",
			3207 => x"0f082b0c",
			3208 => x"0003fb08",
			3209 => x"0705a504",
			3210 => x"ffb832b1",
			3211 => x"017132b1",
			3212 => x"025432b1",
			3213 => x"0100a608",
			3214 => x"0f089504",
			3215 => x"ffd332b1",
			3216 => x"fd3532b1",
			3217 => x"05065104",
			3218 => x"017232b1",
			3219 => x"001232b1",
			3220 => x"00046c10",
			3221 => x"0a02a504",
			3222 => x"fecf32b1",
			3223 => x"0c068b08",
			3224 => x"06017c04",
			3225 => x"008732b1",
			3226 => x"015c32b1",
			3227 => x"fef032b1",
			3228 => x"0a02db10",
			3229 => x"08038808",
			3230 => x"0a02c304",
			3231 => x"fea332b1",
			3232 => x"00ed32b1",
			3233 => x"0f086404",
			3234 => x"fffd32b1",
			3235 => x"fdf532b1",
			3236 => x"0c054608",
			3237 => x"0004dd04",
			3238 => x"016532b1",
			3239 => x"000032b1",
			3240 => x"0b07d604",
			3241 => x"fe7f32b1",
			3242 => x"013032b1",
			3243 => x"fe3032b1",
			3244 => x"0705043c",
			3245 => x"0f083924",
			3246 => x"0306b920",
			3247 => x"040c5808",
			3248 => x"03069604",
			3249 => x"fed133f5",
			3250 => x"000033f5",
			3251 => x"0b05140c",
			3252 => x"02093d08",
			3253 => x"0704f104",
			3254 => x"ff5933f5",
			3255 => x"000033f5",
			3256 => x"000033f5",
			3257 => x"0f081608",
			3258 => x"06016304",
			3259 => x"000033f5",
			3260 => x"012e33f5",
			3261 => x"ffc433f5",
			3262 => x"013633f5",
			3263 => x"03071b14",
			3264 => x"01009310",
			3265 => x"0704f10c",
			3266 => x"040be904",
			3267 => x"007333f5",
			3268 => x"040c7904",
			3269 => x"ffc033f5",
			3270 => x"000033f5",
			3271 => x"ff2a33f5",
			3272 => x"fe6d33f5",
			3273 => x"00f433f5",
			3274 => x"07050818",
			3275 => x"0004580c",
			3276 => x"06016304",
			3277 => x"000033f5",
			3278 => x"0b056504",
			3279 => x"017e33f5",
			3280 => x"000033f5",
			3281 => x"0505cc08",
			3282 => x"0505bd04",
			3283 => x"000033f5",
			3284 => x"ffc533f5",
			3285 => x"000033f5",
			3286 => x"0306e21c",
			3287 => x"0a02cf0c",
			3288 => x"07059108",
			3289 => x"0b054304",
			3290 => x"000033f5",
			3291 => x"fe8933f5",
			3292 => x"000033f5",
			3293 => x"03063a08",
			3294 => x"0d05f704",
			3295 => x"000033f5",
			3296 => x"ffc733f5",
			3297 => x"07051c04",
			3298 => x"00d633f5",
			3299 => x"000033f5",
			3300 => x"05063514",
			3301 => x"0004200c",
			3302 => x"01009904",
			3303 => x"ff2633f5",
			3304 => x"06017404",
			3305 => x"ffb533f5",
			3306 => x"012d33f5",
			3307 => x"040c5204",
			3308 => x"019133f5",
			3309 => x"000033f5",
			3310 => x"0b05d610",
			3311 => x"06019208",
			3312 => x"0b058304",
			3313 => x"000033f5",
			3314 => x"feaa33f5",
			3315 => x"0b05a704",
			3316 => x"007433f5",
			3317 => x"000033f5",
			3318 => x"0003f308",
			3319 => x"05080104",
			3320 => x"006733f5",
			3321 => x"fff933f5",
			3322 => x"0a02a104",
			3323 => x"fe8a33f5",
			3324 => x"000033f5",
			3325 => x"0601855c",
			3326 => x"07065b54",
			3327 => x"0100b438",
			3328 => x"05060620",
			3329 => x"0d061110",
			3330 => x"0c04b908",
			3331 => x"0505b004",
			3332 => x"ff5f3519",
			3333 => x"00853519",
			3334 => x"08037e04",
			3335 => x"fef23519",
			3336 => x"00003519",
			3337 => x"0c04ce08",
			3338 => x"07050104",
			3339 => x"fef63519",
			3340 => x"004c3519",
			3341 => x"07051f04",
			3342 => x"01073519",
			3343 => x"ffff3519",
			3344 => x"0c04cf0c",
			3345 => x"0a02ab08",
			3346 => x"0900fb04",
			3347 => x"009d3519",
			3348 => x"00003519",
			3349 => x"ff713519",
			3350 => x"06018108",
			3351 => x"0100a804",
			3352 => x"fe963519",
			3353 => x"00003519",
			3354 => x"00003519",
			3355 => x"0e098714",
			3356 => x"0c05fc0c",
			3357 => x"0e06e204",
			3358 => x"00003519",
			3359 => x"0901f804",
			3360 => x"00c43519",
			3361 => x"00003519",
			3362 => x"0507b804",
			3363 => x"00003519",
			3364 => x"ff9d3519",
			3365 => x"0a025404",
			3366 => x"ff253519",
			3367 => x"00843519",
			3368 => x"0706cb04",
			3369 => x"fe5e3519",
			3370 => x"00003519",
			3371 => x"05067e0c",
			3372 => x"0c04b504",
			3373 => x"00003519",
			3374 => x"02092e04",
			3375 => x"00003519",
			3376 => x"01453519",
			3377 => x"09014b0c",
			3378 => x"0308c704",
			3379 => x"fe7e3519",
			3380 => x"0100b404",
			3381 => x"00a73519",
			3382 => x"00003519",
			3383 => x"05074808",
			3384 => x"0c050c04",
			3385 => x"00003519",
			3386 => x"01283519",
			3387 => x"0e09e008",
			3388 => x"0901db04",
			3389 => x"fecd3519",
			3390 => x"00003519",
			3391 => x"0003ed08",
			3392 => x"0a025704",
			3393 => x"00003519",
			3394 => x"007c3519",
			3395 => x"0a029b04",
			3396 => x"feee3519",
			3397 => x"001c3519",
			3398 => x"06016c50",
			3399 => x"09019630",
			3400 => x"06016314",
			3401 => x"01009704",
			3402 => x"fe583665",
			3403 => x"0002f604",
			3404 => x"fe673665",
			3405 => x"0f090d08",
			3406 => x"0c056604",
			3407 => x"ffa63665",
			3408 => x"0a783665",
			3409 => x"fe623665",
			3410 => x"03063a04",
			3411 => x"fe5f3665",
			3412 => x"0f07fe0c",
			3413 => x"0c04ea08",
			3414 => x"00043504",
			3415 => x"01973665",
			3416 => x"06353665",
			3417 => x"00473665",
			3418 => x"09017a08",
			3419 => x"0208f704",
			3420 => x"003f3665",
			3421 => x"fe5e3665",
			3422 => x"06433665",
			3423 => x"0209b71c",
			3424 => x"0a01f204",
			3425 => x"04a13665",
			3426 => x"0e08e108",
			3427 => x"0f08dd04",
			3428 => x"011e3665",
			3429 => x"fe633665",
			3430 => x"0d082508",
			3431 => x"01012804",
			3432 => x"04a93665",
			3433 => x"feb83665",
			3434 => x"0c05f504",
			3435 => x"00103665",
			3436 => x"fe613665",
			3437 => x"03ec3665",
			3438 => x"0c065234",
			3439 => x"0a026718",
			3440 => x"01010f04",
			3441 => x"049d3665",
			3442 => x"0d07fd08",
			3443 => x"0e095104",
			3444 => x"fe603665",
			3445 => x"004a3665",
			3446 => x"00035304",
			3447 => x"fe5f3665",
			3448 => x"040a3a04",
			3449 => x"096c3665",
			3450 => x"00ff3665",
			3451 => x"040fc614",
			3452 => x"0505bd08",
			3453 => x"040d8804",
			3454 => x"fe623665",
			3455 => x"01d23665",
			3456 => x"00039604",
			3457 => x"ff853665",
			3458 => x"05086a04",
			3459 => x"02d23665",
			3460 => x"00893665",
			3461 => x"06018104",
			3462 => x"fe703665",
			3463 => x"01c83665",
			3464 => x"0902641c",
			3465 => x"05086a08",
			3466 => x"05083e04",
			3467 => x"fe883665",
			3468 => x"02f83665",
			3469 => x"06017d04",
			3470 => x"01593665",
			3471 => x"0d094e08",
			3472 => x"0100ff04",
			3473 => x"fff53665",
			3474 => x"fe603665",
			3475 => x"0a02ab04",
			3476 => x"001d3665",
			3477 => x"fe5b3665",
			3478 => x"030c6c04",
			3479 => x"fe8b3665",
			3480 => x"040b3665",
			3481 => x"03063a18",
			3482 => x"0a02ed08",
			3483 => x"01009f04",
			3484 => x"fe743751",
			3485 => x"00003751",
			3486 => x"0705180c",
			3487 => x"0b050408",
			3488 => x"0b04ce04",
			3489 => x"fec93751",
			3490 => x"00003751",
			3491 => x"01533751",
			3492 => x"fe883751",
			3493 => x"0005085c",
			3494 => x"0d094e3c",
			3495 => x"0508041c",
			3496 => x"07065810",
			3497 => x"00042508",
			3498 => x"0306b904",
			3499 => x"fdc73751",
			3500 => x"00113751",
			3501 => x"00045b04",
			3502 => x"00ff3751",
			3503 => x"000c3751",
			3504 => x"0f097104",
			3505 => x"fede3751",
			3506 => x"0b06e004",
			3507 => x"018c3751",
			3508 => x"004f3751",
			3509 => x"030a8110",
			3510 => x"05084d08",
			3511 => x"07066d04",
			3512 => x"ffc73751",
			3513 => x"fe303751",
			3514 => x"01011704",
			3515 => x"00a23751",
			3516 => x"fed43751",
			3517 => x"0e0a4808",
			3518 => x"040ac204",
			3519 => x"00003751",
			3520 => x"01e13751",
			3521 => x"030a9904",
			3522 => x"fe093751",
			3523 => x"00003751",
			3524 => x"0706f508",
			3525 => x"0706e304",
			3526 => x"01a13751",
			3527 => x"04fe3751",
			3528 => x"0901d20c",
			3529 => x"0508f804",
			3530 => x"00003751",
			3531 => x"00042d04",
			3532 => x"017c3751",
			3533 => x"00003751",
			3534 => x"0b082408",
			3535 => x"0c068d04",
			3536 => x"006b3751",
			3537 => x"fea13751",
			3538 => x"01073751",
			3539 => x"fe3c3751",
			3540 => x"0802791c",
			3541 => x"07065b18",
			3542 => x"07059104",
			3543 => x"0000382d",
			3544 => x"0b06df10",
			3545 => x"08021e04",
			3546 => x"0000382d",
			3547 => x"0d084c08",
			3548 => x"0507f504",
			3549 => x"00e0382d",
			3550 => x"0000382d",
			3551 => x"0000382d",
			3552 => x"0000382d",
			3553 => x"0000382d",
			3554 => x"06015b04",
			3555 => x"feeb382d",
			3556 => x"0b052414",
			3557 => x"0d05ed10",
			3558 => x"0704ec08",
			3559 => x"0704c004",
			3560 => x"0000382d",
			3561 => x"0000382d",
			3562 => x"07050304",
			3563 => x"ffe8382d",
			3564 => x"0000382d",
			3565 => x"010d382d",
			3566 => x"03073b1c",
			3567 => x"040b6b0c",
			3568 => x"01009304",
			3569 => x"fe78382d",
			3570 => x"040ad504",
			3571 => x"fefd382d",
			3572 => x"003a382d",
			3573 => x"03067808",
			3574 => x"02094d04",
			3575 => x"ff0e382d",
			3576 => x"0000382d",
			3577 => x"02090c04",
			3578 => x"012c382d",
			3579 => x"0000382d",
			3580 => x"0f08d410",
			3581 => x"0b058308",
			3582 => x"0e075804",
			3583 => x"0156382d",
			3584 => x"0000382d",
			3585 => x"0705a204",
			3586 => x"0000382d",
			3587 => x"0060382d",
			3588 => x"08036608",
			3589 => x"040cd804",
			3590 => x"fff8382d",
			3591 => x"00e7382d",
			3592 => x"0e0c7e04",
			3593 => x"ff6d382d",
			3594 => x"005d382d",
			3595 => x"030a997c",
			3596 => x"0d08725c",
			3597 => x"0309c03c",
			3598 => x"0208e41c",
			3599 => x"0208ab10",
			3600 => x"0e06f708",
			3601 => x"0600e804",
			3602 => x"00003979",
			3603 => x"ff153979",
			3604 => x"0b061b04",
			3605 => x"00423979",
			3606 => x"00003979",
			3607 => x"0c049404",
			3608 => x"00003979",
			3609 => x"0c04d204",
			3610 => x"01113979",
			3611 => x"00013979",
			3612 => x"00042810",
			3613 => x"0705d108",
			3614 => x"0c04ed04",
			3615 => x"ffdd3979",
			3616 => x"feac3979",
			3617 => x"0802be04",
			3618 => x"ffcd3979",
			3619 => x"006f3979",
			3620 => x"00042e08",
			3621 => x"0a02a504",
			3622 => x"00003979",
			3623 => x"013d3979",
			3624 => x"0308a904",
			3625 => x"ffbe3979",
			3626 => x"004e3979",
			3627 => x"00037d10",
			3628 => x"030a120c",
			3629 => x"040a3a04",
			3630 => x"00003979",
			3631 => x"0c061304",
			3632 => x"00513979",
			3633 => x"00003979",
			3634 => x"ffbb3979",
			3635 => x"0902190c",
			3636 => x"0601bb08",
			3637 => x"0b06fe04",
			3638 => x"012e3979",
			3639 => x"00003979",
			3640 => x"00003979",
			3641 => x"00003979",
			3642 => x"020a8314",
			3643 => x"0b072008",
			3644 => x"0c063004",
			3645 => x"ff243979",
			3646 => x"00003979",
			3647 => x"0c065008",
			3648 => x"00033e04",
			3649 => x"00003979",
			3650 => x"00e23979",
			3651 => x"00003979",
			3652 => x"0901d704",
			3653 => x"00003979",
			3654 => x"0d087f04",
			3655 => x"00003979",
			3656 => x"fe5d3979",
			3657 => x"0d0a1e24",
			3658 => x"0f0aed0c",
			3659 => x"00037804",
			3660 => x"00003979",
			3661 => x"030aa104",
			3662 => x"00003979",
			3663 => x"ff6f3979",
			3664 => x"07065704",
			3665 => x"00003979",
			3666 => x"0a025f04",
			3667 => x"00003979",
			3668 => x"0901ee08",
			3669 => x"0601af04",
			3670 => x"003b3979",
			3671 => x"00003979",
			3672 => x"06018a04",
			3673 => x"00003979",
			3674 => x"00c33979",
			3675 => x"0c071e04",
			3676 => x"ff1a3979",
			3677 => x"00003979",
			3678 => x"01014570",
			3679 => x"0208e430",
			3680 => x"0208ab10",
			3681 => x"0e06f708",
			3682 => x"0600e804",
			3683 => x"00003abd",
			3684 => x"ff213abd",
			3685 => x"0b061b04",
			3686 => x"003c3abd",
			3687 => x"00003abd",
			3688 => x"0c049404",
			3689 => x"00003abd",
			3690 => x"0c04d20c",
			3691 => x"06016304",
			3692 => x"00003abd",
			3693 => x"0b051204",
			3694 => x"00003abd",
			3695 => x"011e3abd",
			3696 => x"0c04ed08",
			3697 => x"0d063804",
			3698 => x"ff5e3abd",
			3699 => x"00003abd",
			3700 => x"09014b04",
			3701 => x"00aa3abd",
			3702 => x"00003abd",
			3703 => x"0d09222c",
			3704 => x"0d08721c",
			3705 => x"0d075510",
			3706 => x"07051f08",
			3707 => x"040b6304",
			3708 => x"ff683abd",
			3709 => x"00263abd",
			3710 => x"06019604",
			3711 => x"fede3abd",
			3712 => x"00003abd",
			3713 => x"0100d204",
			3714 => x"00f43abd",
			3715 => x"040c6004",
			3716 => x"000e3abd",
			3717 => x"ff303abd",
			3718 => x"09019c08",
			3719 => x"0100fa04",
			3720 => x"00003abd",
			3721 => x"00233abd",
			3722 => x"0e0aee04",
			3723 => x"fed53abd",
			3724 => x"00003abd",
			3725 => x"0d0a5f10",
			3726 => x"0601af0c",
			3727 => x"0100f504",
			3728 => x"00003abd",
			3729 => x"0508b304",
			3730 => x"00003abd",
			3731 => x"00e73abd",
			3732 => x"00003abd",
			3733 => x"00003abd",
			3734 => x"0c06cb30",
			3735 => x"0101490c",
			3736 => x"0706a108",
			3737 => x"0e0a4804",
			3738 => x"01173abd",
			3739 => x"00003abd",
			3740 => x"00003abd",
			3741 => x"01015e14",
			3742 => x"08034c10",
			3743 => x"0f0aed08",
			3744 => x"07067004",
			3745 => x"00003abd",
			3746 => x"ff863abd",
			3747 => x"0706f504",
			3748 => x"00c73abd",
			3749 => x"ffeb3abd",
			3750 => x"ff703abd",
			3751 => x"0f0afc04",
			3752 => x"00003abd",
			3753 => x"0e0adc04",
			3754 => x"00003abd",
			3755 => x"06018e04",
			3756 => x"00003abd",
			3757 => x"00e63abd",
			3758 => x"ff363abd",
			3759 => x"0505af08",
			3760 => x"0804ac04",
			3761 => x"fecf3bb1",
			3762 => x"00003bb1",
			3763 => x"0c04ca14",
			3764 => x"040bb208",
			3765 => x"0900fe04",
			3766 => x"ff143bb1",
			3767 => x"006d3bb1",
			3768 => x"0505b004",
			3769 => x"00003bb1",
			3770 => x"06016404",
			3771 => x"00003bb1",
			3772 => x"01693bb1",
			3773 => x"040a5b2c",
			3774 => x"0b06bc14",
			3775 => x"0a027810",
			3776 => x"0c05fa08",
			3777 => x"0e05ac04",
			3778 => x"00003bb1",
			3779 => x"ff3b3bb1",
			3780 => x"00034604",
			3781 => x"00003bb1",
			3782 => x"00413bb1",
			3783 => x"00af3bb1",
			3784 => x"0507bb08",
			3785 => x"01010f04",
			3786 => x"00003bb1",
			3787 => x"018b3bb1",
			3788 => x"0a021d08",
			3789 => x"09019c04",
			3790 => x"ff8a3bb1",
			3791 => x"00d73bb1",
			3792 => x"040a0104",
			3793 => x"ff293bb1",
			3794 => x"00003bb1",
			3795 => x"0601851c",
			3796 => x"0c060f10",
			3797 => x"0003f208",
			3798 => x"040bd604",
			3799 => x"fe833bb1",
			3800 => x"00183bb1",
			3801 => x"0704ef04",
			3802 => x"00cd3bb1",
			3803 => x"ff933bb1",
			3804 => x"01011b04",
			3805 => x"00d93bb1",
			3806 => x"0802d404",
			3807 => x"ff7f3bb1",
			3808 => x"002d3bb1",
			3809 => x"0b057408",
			3810 => x"01008204",
			3811 => x"00003bb1",
			3812 => x"015d3bb1",
			3813 => x"0c06c708",
			3814 => x"09011b04",
			3815 => x"ff003bb1",
			3816 => x"002c3bb1",
			3817 => x"0509e304",
			3818 => x"feab3bb1",
			3819 => x"00003bb1",
			3820 => x"0b051408",
			3821 => x"02093d04",
			3822 => x"feaf3cbd",
			3823 => x"00003cbd",
			3824 => x"00043a40",
			3825 => x"08035e34",
			3826 => x"0a02a820",
			3827 => x"040b8310",
			3828 => x"01012608",
			3829 => x"01012404",
			3830 => x"fff63cbd",
			3831 => x"fd623cbd",
			3832 => x"00039204",
			3833 => x"00123cbd",
			3834 => x"00b93cbd",
			3835 => x"020b0f08",
			3836 => x"0003ee04",
			3837 => x"ffc63cbd",
			3838 => x"fdd83cbd",
			3839 => x"040c3204",
			3840 => x"00813cbd",
			3841 => x"ff863cbd",
			3842 => x"0004200c",
			3843 => x"0100bc04",
			3844 => x"ff7d3cbd",
			3845 => x"05084d04",
			3846 => x"01033cbd",
			3847 => x"fff93cbd",
			3848 => x"0601ba04",
			3849 => x"01743cbd",
			3850 => x"00003cbd",
			3851 => x"0100d004",
			3852 => x"fe933cbd",
			3853 => x"01014704",
			3854 => x"00003cbd",
			3855 => x"ff503cbd",
			3856 => x"020bd730",
			3857 => x"00045814",
			3858 => x"040bbf08",
			3859 => x"06018004",
			3860 => x"fe633cbd",
			3861 => x"00163cbd",
			3862 => x"0900cb04",
			3863 => x"00003cbd",
			3864 => x"0a02a904",
			3865 => x"00003cbd",
			3866 => x"01a83cbd",
			3867 => x"0a02bf0c",
			3868 => x"0208c708",
			3869 => x"040c5e04",
			3870 => x"00003cbd",
			3871 => x"003f3cbd",
			3872 => x"fec93cbd",
			3873 => x"08038808",
			3874 => x"06017004",
			3875 => x"00003cbd",
			3876 => x"01463cbd",
			3877 => x"0a02db04",
			3878 => x"ff3c3cbd",
			3879 => x"00423cbd",
			3880 => x"0e0cbb08",
			3881 => x"0601c404",
			3882 => x"00003cbd",
			3883 => x"fe683cbd",
			3884 => x"0601ec04",
			3885 => x"01053cbd",
			3886 => x"fffa3cbd",
			3887 => x"040ae244",
			3888 => x"0409db18",
			3889 => x"03097814",
			3890 => x"0a021d10",
			3891 => x"0b06cd0c",
			3892 => x"01010f04",
			3893 => x"00003e29",
			3894 => x"0b06bc04",
			3895 => x"00003e29",
			3896 => x"00e93e29",
			3897 => x"00003e29",
			3898 => x"00003e29",
			3899 => x"ff9a3e29",
			3900 => x"030a121c",
			3901 => x"0c056210",
			3902 => x"0c04ec08",
			3903 => x"0306ff04",
			3904 => x"00003e29",
			3905 => x"00bb3e29",
			3906 => x"0c050504",
			3907 => x"00003e29",
			3908 => x"ff843e29",
			3909 => x"0c061408",
			3910 => x"09021504",
			3911 => x"00e63e29",
			3912 => x"00003e29",
			3913 => x"00003e29",
			3914 => x"0c062e08",
			3915 => x"020a5b04",
			3916 => x"ff353e29",
			3917 => x"00003e29",
			3918 => x"0c065004",
			3919 => x"00a63e29",
			3920 => x"00003e29",
			3921 => x"040aef0c",
			3922 => x"06018e08",
			3923 => x"0003f704",
			3924 => x"febe3e29",
			3925 => x"00003e29",
			3926 => x"00003e29",
			3927 => x"020ab738",
			3928 => x"0b05631c",
			3929 => x"0306c510",
			3930 => x"01007d08",
			3931 => x"0b051104",
			3932 => x"ffe83e29",
			3933 => x"00903e29",
			3934 => x"0b052404",
			3935 => x"00003e29",
			3936 => x"ff573e29",
			3937 => x"0f087204",
			3938 => x"01433e29",
			3939 => x"06017804",
			3940 => x"ff753e29",
			3941 => x"00273e29",
			3942 => x"040b360c",
			3943 => x"06018804",
			3944 => x"00003e29",
			3945 => x"0a026704",
			3946 => x"00003e29",
			3947 => x"00793e29",
			3948 => x"0a02bf08",
			3949 => x"0901db04",
			3950 => x"fed03e29",
			3951 => x"00003e29",
			3952 => x"0b05bf04",
			3953 => x"00803e29",
			3954 => x"ff613e29",
			3955 => x"0601c018",
			3956 => x"040b460c",
			3957 => x"030b2a08",
			3958 => x"0b072f04",
			3959 => x"00003e29",
			3960 => x"ffa83e29",
			3961 => x"00003e29",
			3962 => x"0a02fd08",
			3963 => x"0e0bef04",
			3964 => x"00983e29",
			3965 => x"00003e29",
			3966 => x"00003e29",
			3967 => x"0e0c7e10",
			3968 => x"020bbc08",
			3969 => x"01014704",
			3970 => x"00003e29",
			3971 => x"00043e29",
			3972 => x"08036804",
			3973 => x"00003e29",
			3974 => x"feb03e29",
			3975 => x"0d09f804",
			3976 => x"00543e29",
			3977 => x"00003e29",
			3978 => x"0003ee5c",
			3979 => x"07059110",
			3980 => x"0c04ec08",
			3981 => x"06017004",
			3982 => x"00003fbd",
			3983 => x"001a3fbd",
			3984 => x"07050804",
			3985 => x"00003fbd",
			3986 => x"ff293fbd",
			3987 => x"0d087224",
			3988 => x"00036814",
			3989 => x"0a02390c",
			3990 => x"0507f508",
			3991 => x"0c061404",
			3992 => x"006f3fbd",
			3993 => x"00003fbd",
			3994 => x"00003fbd",
			3995 => x"0802c304",
			3996 => x"ff6e3fbd",
			3997 => x"00003fbd",
			3998 => x"0902120c",
			3999 => x"0c056304",
			4000 => x"00003fbd",
			4001 => x"0a024104",
			4002 => x"00003fbd",
			4003 => x"00e93fbd",
			4004 => x"00003fbd",
			4005 => x"0c062e0c",
			4006 => x"0003af08",
			4007 => x"030a1204",
			4008 => x"00003fbd",
			4009 => x"fee73fbd",
			4010 => x"00003fbd",
			4011 => x"0601930c",
			4012 => x"0d08b304",
			4013 => x"00003fbd",
			4014 => x"05090a04",
			4015 => x"00943fbd",
			4016 => x"00003fbd",
			4017 => x"08031a08",
			4018 => x"0d08b304",
			4019 => x"00003fbd",
			4020 => x"ff913fbd",
			4021 => x"0e0aaa04",
			4022 => x"00003fbd",
			4023 => x"004f3fbd",
			4024 => x"05061528",
			4025 => x"0d062b20",
			4026 => x"07050814",
			4027 => x"0f088b10",
			4028 => x"0d061108",
			4029 => x"0c04b904",
			4030 => x"004f3fbd",
			4031 => x"ffbd3fbd",
			4032 => x"03068304",
			4033 => x"00003fbd",
			4034 => x"00eb3fbd",
			4035 => x"ff343fbd",
			4036 => x"0306c508",
			4037 => x"02098104",
			4038 => x"ff133fbd",
			4039 => x"00003fbd",
			4040 => x"00003fbd",
			4041 => x"0306a504",
			4042 => x"00003fbd",
			4043 => x"01093fbd",
			4044 => x"020ab724",
			4045 => x"0a029e08",
			4046 => x"0e06ce04",
			4047 => x"00003fbd",
			4048 => x"feb53fbd",
			4049 => x"07054510",
			4050 => x"0c04d208",
			4051 => x"0d064704",
			4052 => x"00253fbd",
			4053 => x"ff423fbd",
			4054 => x"06017404",
			4055 => x"00003fbd",
			4056 => x"00f73fbd",
			4057 => x"0e08fd08",
			4058 => x"0b057604",
			4059 => x"00003fbd",
			4060 => x"fee93fbd",
			4061 => x"001c3fbd",
			4062 => x"0601cc18",
			4063 => x"020b8b0c",
			4064 => x"0c061204",
			4065 => x"003b3fbd",
			4066 => x"0e0abb04",
			4067 => x"ff4a3fbd",
			4068 => x"00003fbd",
			4069 => x"0706f908",
			4070 => x"08038d04",
			4071 => x"00f73fbd",
			4072 => x"00003fbd",
			4073 => x"00003fbd",
			4074 => x"020bd704",
			4075 => x"00263fbd",
			4076 => x"0e0cf604",
			4077 => x"fec93fbd",
			4078 => x"00003fbd",
			4079 => x"03065938",
			4080 => x"03063228",
			4081 => x"0305e118",
			4082 => x"0305a004",
			4083 => x"fe554139",
			4084 => x"02093d0c",
			4085 => x"0208d404",
			4086 => x"fe554139",
			4087 => x"0208d604",
			4088 => x"004c4139",
			4089 => x"fe864139",
			4090 => x"0209b104",
			4091 => x"017c4139",
			4092 => x"fec94139",
			4093 => x"0a02f308",
			4094 => x"0b059504",
			4095 => x"fe554139",
			4096 => x"026f4139",
			4097 => x"07050804",
			4098 => x"04c44139",
			4099 => x"fe794139",
			4100 => x"00047c04",
			4101 => x"fe564139",
			4102 => x"07051c08",
			4103 => x"0f082b04",
			4104 => x"06554139",
			4105 => x"fe824139",
			4106 => x"fe6b4139",
			4107 => x"0c065268",
			4108 => x"0a025934",
			4109 => x"0f095618",
			4110 => x"03078c0c",
			4111 => x"0705a504",
			4112 => x"fe654139",
			4113 => x"0f071704",
			4114 => x"fec04139",
			4115 => x"0af34139",
			4116 => x"0100fc04",
			4117 => x"fe574139",
			4118 => x"08025f04",
			4119 => x"03dd4139",
			4120 => x"fec74139",
			4121 => x"0507f510",
			4122 => x"0901b808",
			4123 => x"0c05f404",
			4124 => x"03124139",
			4125 => x"08424139",
			4126 => x"0d07fd04",
			4127 => x"fed84139",
			4128 => x"01be4139",
			4129 => x"0d08b304",
			4130 => x"fe5a4139",
			4131 => x"01014504",
			4132 => x"06d74139",
			4133 => x"fec24139",
			4134 => x"0306c51c",
			4135 => x"0c04ea10",
			4136 => x"0a02a608",
			4137 => x"0d061d04",
			4138 => x"fe6e4139",
			4139 => x"00de4139",
			4140 => x"0d05ed04",
			4141 => x"fe664139",
			4142 => x"04724139",
			4143 => x"07051808",
			4144 => x"0f082204",
			4145 => x"03834139",
			4146 => x"fe3b4139",
			4147 => x"fe5c4139",
			4148 => x"05086a10",
			4149 => x"0e098708",
			4150 => x"0c052704",
			4151 => x"04374139",
			4152 => x"ffc54139",
			4153 => x"00039604",
			4154 => x"023e4139",
			4155 => x"04624139",
			4156 => x"00040304",
			4157 => x"fe604139",
			4158 => x"04e44139",
			4159 => x"09026b18",
			4160 => x"0d08b304",
			4161 => x"02444139",
			4162 => x"0b076308",
			4163 => x"0c066c04",
			4164 => x"03a14139",
			4165 => x"fe774139",
			4166 => x"05088604",
			4167 => x"00324139",
			4168 => x"0706b704",
			4169 => x"fff74139",
			4170 => x"fe704139",
			4171 => x"00042904",
			4172 => x"fe9a4139",
			4173 => x"04724139",
			4174 => x"01014588",
			4175 => x"02095140",
			4176 => x"03073b24",
			4177 => x"0a02920c",
			4178 => x"05060604",
			4179 => x"0000429d",
			4180 => x"040a4904",
			4181 => x"0000429d",
			4182 => x"fe9d429d",
			4183 => x"0705180c",
			4184 => x"09010208",
			4185 => x"07050104",
			4186 => x"0000429d",
			4187 => x"00d1429d",
			4188 => x"ff82429d",
			4189 => x"0306ff08",
			4190 => x"01007804",
			4191 => x"0000429d",
			4192 => x"ff2b429d",
			4193 => x"0000429d",
			4194 => x"0307c408",
			4195 => x"06011d04",
			4196 => x"0000429d",
			4197 => x"010a429d",
			4198 => x"02094d10",
			4199 => x"0c062e08",
			4200 => x"0c05d704",
			4201 => x"0000429d",
			4202 => x"ff6c429d",
			4203 => x"0c063004",
			4204 => x"0020429d",
			4205 => x"0000429d",
			4206 => x"0035429d",
			4207 => x"06019630",
			4208 => x"0c05bc18",
			4209 => x"0a02b00c",
			4210 => x"0901d708",
			4211 => x"040a9504",
			4212 => x"0000429d",
			4213 => x"fe9a429d",
			4214 => x"0000429d",
			4215 => x"08036304",
			4216 => x"0122429d",
			4217 => x"0f087204",
			4218 => x"0000429d",
			4219 => x"ff1f429d",
			4220 => x"0101170c",
			4221 => x"06019008",
			4222 => x"06016004",
			4223 => x"ffe7429d",
			4224 => x"00d6429d",
			4225 => x"ffc7429d",
			4226 => x"07066d08",
			4227 => x"07065804",
			4228 => x"ffcf429d",
			4229 => x"0053429d",
			4230 => x"fe8d429d",
			4231 => x"0c054c08",
			4232 => x"0a031804",
			4233 => x"00f4429d",
			4234 => x"0000429d",
			4235 => x"0803630c",
			4236 => x"07068604",
			4237 => x"00f5429d",
			4238 => x"020b7704",
			4239 => x"feed429d",
			4240 => x"00b6429d",
			4241 => x"fee6429d",
			4242 => x"0c06cb28",
			4243 => x"01014908",
			4244 => x"0706a104",
			4245 => x"00f7429d",
			4246 => x"0000429d",
			4247 => x"01015f18",
			4248 => x"030b3a10",
			4249 => x"0f0aed08",
			4250 => x"07067004",
			4251 => x"0000429d",
			4252 => x"ff90429d",
			4253 => x"0706f504",
			4254 => x"00c5429d",
			4255 => x"0000429d",
			4256 => x"01015b04",
			4257 => x"ff5c429d",
			4258 => x"0000429d",
			4259 => x"030b2a04",
			4260 => x"0000429d",
			4261 => x"00d9429d",
			4262 => x"ff41429d",
			4263 => x"040b304c",
			4264 => x"00040244",
			4265 => x"0c05f81c",
			4266 => x"0a02a118",
			4267 => x"0003ee10",
			4268 => x"040a7b08",
			4269 => x"00034b04",
			4270 => x"ffd843e9",
			4271 => x"002443e9",
			4272 => x"0901d704",
			4273 => x"ff0d43e9",
			4274 => x"000043e9",
			4275 => x"0306c504",
			4276 => x"000043e9",
			4277 => x"00c543e9",
			4278 => x"fef843e9",
			4279 => x"0c065014",
			4280 => x"0100e804",
			4281 => x"000043e9",
			4282 => x"09020a08",
			4283 => x"020aa604",
			4284 => x"00a443e9",
			4285 => x"000043e9",
			4286 => x"040acf04",
			4287 => x"002c43e9",
			4288 => x"000043e9",
			4289 => x"0f0aed08",
			4290 => x"0508dd04",
			4291 => x"ff9943e9",
			4292 => x"000043e9",
			4293 => x"0802e304",
			4294 => x"000043e9",
			4295 => x"00039604",
			4296 => x"004843e9",
			4297 => x"000043e9",
			4298 => x"0306b904",
			4299 => x"000043e9",
			4300 => x"011d43e9",
			4301 => x"040b4610",
			4302 => x"0a026404",
			4303 => x"000043e9",
			4304 => x"0c04ea04",
			4305 => x"000043e9",
			4306 => x"040b3604",
			4307 => x"000043e9",
			4308 => x"fe7643e9",
			4309 => x"0003ed14",
			4310 => x"0309b004",
			4311 => x"000043e9",
			4312 => x"0902300c",
			4313 => x"0a02a008",
			4314 => x"0802e604",
			4315 => x"000043e9",
			4316 => x"00c043e9",
			4317 => x"000043e9",
			4318 => x"000043e9",
			4319 => x"0a02a618",
			4320 => x"020b160c",
			4321 => x"0e0aa408",
			4322 => x"0003ee04",
			4323 => x"000043e9",
			4324 => x"fe8e43e9",
			4325 => x"000043e9",
			4326 => x"01014e08",
			4327 => x"0e0b9404",
			4328 => x"008743e9",
			4329 => x"000043e9",
			4330 => x"000043e9",
			4331 => x"02096010",
			4332 => x"0306e208",
			4333 => x"02091904",
			4334 => x"006e43e9",
			4335 => x"ff8343e9",
			4336 => x"0a02bc04",
			4337 => x"015043e9",
			4338 => x"000043e9",
			4339 => x"00043a08",
			4340 => x"0e090704",
			4341 => x"ff0f43e9",
			4342 => x"000043e9",
			4343 => x"00047904",
			4344 => x"005643e9",
			4345 => x"ff9643e9",
			4346 => x"03063214",
			4347 => x"01009d10",
			4348 => x"0305a004",
			4349 => x"fe56451d",
			4350 => x"0803be04",
			4351 => x"fe56451d",
			4352 => x"07050804",
			4353 => x"0440451d",
			4354 => x"fe73451d",
			4355 => x"01d8451d",
			4356 => x"0c065264",
			4357 => x"0802d228",
			4358 => x"0003020c",
			4359 => x"01010608",
			4360 => x"08026f04",
			4361 => x"fe63451d",
			4362 => x"00df451d",
			4363 => x"031a451d",
			4364 => x"0409a00c",
			4365 => x"0d082408",
			4366 => x"0c059f04",
			4367 => x"feae451d",
			4368 => x"054d451d",
			4369 => x"fe6b451d",
			4370 => x"03092208",
			4371 => x"0c05f804",
			4372 => x"fe5d451d",
			4373 => x"0021451d",
			4374 => x"00037804",
			4375 => x"ffca451d",
			4376 => x"05f3451d",
			4377 => x"0306c520",
			4378 => x"040c0410",
			4379 => x"0306a508",
			4380 => x"03069604",
			4381 => x"fe55451d",
			4382 => x"ff9a451d",
			4383 => x"0208f704",
			4384 => x"0328451d",
			4385 => x"fe37451d",
			4386 => x"0f082b08",
			4387 => x"07051c04",
			4388 => x"04b5451d",
			4389 => x"fe6a451d",
			4390 => x"0306b904",
			4391 => x"fe5a451d",
			4392 => x"0116451d",
			4393 => x"040c6c10",
			4394 => x"0802f808",
			4395 => x"040ac904",
			4396 => x"0423451d",
			4397 => x"ffcc451d",
			4398 => x"0706a104",
			4399 => x"0376451d",
			4400 => x"fe78451d",
			4401 => x"0c04f104",
			4402 => x"03e1451d",
			4403 => x"0f09a304",
			4404 => x"fe56451d",
			4405 => x"018e451d",
			4406 => x"0902641c",
			4407 => x"05086a08",
			4408 => x"0e09c104",
			4409 => x"fe78451d",
			4410 => x"03de451d",
			4411 => x"08034510",
			4412 => x"040cb608",
			4413 => x"01010604",
			4414 => x"0bff451d",
			4415 => x"fe89451d",
			4416 => x"08034204",
			4417 => x"2162451d",
			4418 => x"0573451d",
			4419 => x"fe58451d",
			4420 => x"030c6c04",
			4421 => x"fe82451d",
			4422 => x"05a0451d",
			4423 => x"0b05110c",
			4424 => x"0a035d04",
			4425 => x"fe6a4609",
			4426 => x"0006a004",
			4427 => x"01004609",
			4428 => x"00004609",
			4429 => x"0a032364",
			4430 => x"0802aa28",
			4431 => x"0409db14",
			4432 => x"03097810",
			4433 => x"0f095608",
			4434 => x"0507b804",
			4435 => x"00db4609",
			4436 => x"ff234609",
			4437 => x"0b06dc04",
			4438 => x"02d54609",
			4439 => x"ffd04609",
			4440 => x"fe834609",
			4441 => x"0c063010",
			4442 => x"0c05f208",
			4443 => x"0c05d604",
			4444 => x"00904609",
			4445 => x"ffad4609",
			4446 => x"0c061204",
			4447 => x"03074609",
			4448 => x"01604609",
			4449 => x"ff214609",
			4450 => x"040cbf20",
			4451 => x"0306b910",
			4452 => x"040bb708",
			4453 => x"0f082204",
			4454 => x"fe4a4609",
			4455 => x"fcd94609",
			4456 => x"0c04b204",
			4457 => x"01b24609",
			4458 => x"ff874609",
			4459 => x"0f083908",
			4460 => x"07051804",
			4461 => x"023c4609",
			4462 => x"00004609",
			4463 => x"03071b04",
			4464 => x"ff3d4609",
			4465 => x"00404609",
			4466 => x"0b05450c",
			4467 => x"0505af04",
			4468 => x"00004609",
			4469 => x"0c04ec04",
			4470 => x"01d64609",
			4471 => x"00874609",
			4472 => x"03069608",
			4473 => x"03067804",
			4474 => x"fdbf4609",
			4475 => x"ffc54609",
			4476 => x"040ceb04",
			4477 => x"01cb4609",
			4478 => x"004a4609",
			4479 => x"0c04e904",
			4480 => x"01534609",
			4481 => x"fe1d4609",
			4482 => x"06016c60",
			4483 => x"09019638",
			4484 => x"0601631c",
			4485 => x"01009704",
			4486 => x"fe5a4795",
			4487 => x"0002f60c",
			4488 => x"0d070808",
			4489 => x"0b05f804",
			4490 => x"fe6f4795",
			4491 => x"041a4795",
			4492 => x"fe5e4795",
			4493 => x"0f090d08",
			4494 => x"07059104",
			4495 => x"fe884795",
			4496 => x"061b4795",
			4497 => x"fe684795",
			4498 => x"03063a04",
			4499 => x"fe614795",
			4500 => x"0f07fe0c",
			4501 => x"0c04ea08",
			4502 => x"03065904",
			4503 => x"023d4795",
			4504 => x"05764795",
			4505 => x"003b4795",
			4506 => x"09017a08",
			4507 => x"0208f704",
			4508 => x"00364795",
			4509 => x"fe624795",
			4510 => x"04904795",
			4511 => x"02099518",
			4512 => x"0a01f204",
			4513 => x"03644795",
			4514 => x"0c05f610",
			4515 => x"03092e08",
			4516 => x"02090004",
			4517 => x"001a4795",
			4518 => x"fe6b4795",
			4519 => x"0d081804",
			4520 => x"05344795",
			4521 => x"ffd24795",
			4522 => x"fe664795",
			4523 => x"06016a0c",
			4524 => x"0c061004",
			4525 => x"06c94795",
			4526 => x"06015f04",
			4527 => x"fec84795",
			4528 => x"01224795",
			4529 => x"fe9a4795",
			4530 => x"0c065244",
			4531 => x"0a02671c",
			4532 => x"01010f04",
			4533 => x"034f4795",
			4534 => x"0e092408",
			4535 => x"0a023004",
			4536 => x"01b24795",
			4537 => x"fe624795",
			4538 => x"0b06ee08",
			4539 => x"01012304",
			4540 => x"08054795",
			4541 => x"01034795",
			4542 => x"0d08b304",
			4543 => x"fe164795",
			4544 => x"010f4795",
			4545 => x"00055420",
			4546 => x"06017910",
			4547 => x"07052f08",
			4548 => x"0505bd04",
			4549 => x"fe6f4795",
			4550 => x"026e4795",
			4551 => x"020a5b04",
			4552 => x"fe4d4795",
			4553 => x"00fe4795",
			4554 => x"0706a108",
			4555 => x"00039604",
			4556 => x"ffa74795",
			4557 => x"02854795",
			4558 => x"030b4104",
			4559 => x"fe5c4795",
			4560 => x"02984795",
			4561 => x"06018104",
			4562 => x"fe774795",
			4563 => x"00004795",
			4564 => x"0902641c",
			4565 => x"05086a08",
			4566 => x"0f0aad04",
			4567 => x"fe7b4795",
			4568 => x"02a94795",
			4569 => x"06017d04",
			4570 => x"012c4795",
			4571 => x"0d094e08",
			4572 => x"0706c904",
			4573 => x"ff754795",
			4574 => x"fe5c4795",
			4575 => x"0a02ab04",
			4576 => x"00344795",
			4577 => x"fe5d4795",
			4578 => x"030c6c04",
			4579 => x"fe964795",
			4580 => x"03394795",
			4581 => x"09012754",
			4582 => x"0b055628",
			4583 => x"06016304",
			4584 => x"febb48d1",
			4585 => x"0c050920",
			4586 => x"02092810",
			4587 => x"0306a508",
			4588 => x"040c5804",
			4589 => x"ff7848d1",
			4590 => x"00e948d1",
			4591 => x"0e072504",
			4592 => x"016448d1",
			4593 => x"000048d1",
			4594 => x"02093d08",
			4595 => x"0704ef04",
			4596 => x"000048d1",
			4597 => x"febf48d1",
			4598 => x"0d060f04",
			4599 => x"ff4148d1",
			4600 => x"009948d1",
			4601 => x"fe1a48d1",
			4602 => x"06019124",
			4603 => x"040b5618",
			4604 => x"0c04e908",
			4605 => x"06017004",
			4606 => x"000048d1",
			4607 => x"00fe48d1",
			4608 => x"0c054c08",
			4609 => x"05062604",
			4610 => x"000048d1",
			4611 => x"febb48d1",
			4612 => x"06010304",
			4613 => x"000048d1",
			4614 => x"00aa48d1",
			4615 => x"0505f904",
			4616 => x"000048d1",
			4617 => x"03077c04",
			4618 => x"fe4448d1",
			4619 => x"ffcd48d1",
			4620 => x"09011304",
			4621 => x"00e648d1",
			4622 => x"000048d1",
			4623 => x"05067e04",
			4624 => x"017748d1",
			4625 => x"0308c714",
			4626 => x"00043a08",
			4627 => x"02091b04",
			4628 => x"000048d1",
			4629 => x"fe7148d1",
			4630 => x"040dca08",
			4631 => x"07058b04",
			4632 => x"013548d1",
			4633 => x"000048d1",
			4634 => x"ff9c48d1",
			4635 => x"0d082520",
			4636 => x"0c05f610",
			4637 => x"0f096008",
			4638 => x"08028704",
			4639 => x"000048d1",
			4640 => x"ff7e48d1",
			4641 => x"0f0abc04",
			4642 => x"014548d1",
			4643 => x"000048d1",
			4644 => x"0c05f908",
			4645 => x"0507c904",
			4646 => x"fecb48d1",
			4647 => x"000048d1",
			4648 => x"0c061404",
			4649 => x"00cc48d1",
			4650 => x"000048d1",
			4651 => x"0c05d404",
			4652 => x"feac48d1",
			4653 => x"06016208",
			4654 => x"09019604",
			4655 => x"ffaa48d1",
			4656 => x"00d148d1",
			4657 => x"030a2804",
			4658 => x"ff5948d1",
			4659 => x"002748d1",
			4660 => x"0e078e60",
			4661 => x"0b055638",
			4662 => x"040ad50c",
			4663 => x"0c04d204",
			4664 => x"00004aad",
			4665 => x"0d063704",
			4666 => x"fe944aad",
			4667 => x"00004aad",
			4668 => x"0306a51c",
			4669 => x"040c9310",
			4670 => x"0b053108",
			4671 => x"06017004",
			4672 => x"ff6f4aad",
			4673 => x"00a64aad",
			4674 => x"0704ea04",
			4675 => x"00004aad",
			4676 => x"fee34aad",
			4677 => x"0505a004",
			4678 => x"ffd64aad",
			4679 => x"07051b04",
			4680 => x"00c44aad",
			4681 => x"ffe24aad",
			4682 => x"0f088e08",
			4683 => x"0d061104",
			4684 => x"00004aad",
			4685 => x"015b4aad",
			4686 => x"0d063f04",
			4687 => x"fedb4aad",
			4688 => x"00804aad",
			4689 => x"0208e214",
			4690 => x"040abb0c",
			4691 => x"0f07a604",
			4692 => x"00004aad",
			4693 => x"0003b804",
			4694 => x"ffbf4aad",
			4695 => x"00004aad",
			4696 => x"00040304",
			4697 => x"00a14aad",
			4698 => x"00004aad",
			4699 => x"06018d0c",
			4700 => x"0c04cc04",
			4701 => x"00004aad",
			4702 => x"09012004",
			4703 => x"fe714aad",
			4704 => x"00004aad",
			4705 => x"05063304",
			4706 => x"00464aad",
			4707 => x"00004aad",
			4708 => x"0507f63c",
			4709 => x"06018c2c",
			4710 => x"0c059910",
			4711 => x"040c4c0c",
			4712 => x"0b058304",
			4713 => x"00004aad",
			4714 => x"0705d104",
			4715 => x"fea54aad",
			4716 => x"00004aad",
			4717 => x"004c4aad",
			4718 => x"0901c30c",
			4719 => x"0d084c08",
			4720 => x"00030204",
			4721 => x"00004aad",
			4722 => x"00e14aad",
			4723 => x"00004aad",
			4724 => x"040a0108",
			4725 => x"0b06be04",
			4726 => x"00004aad",
			4727 => x"ff3a4aad",
			4728 => x"040aa904",
			4729 => x"005b4aad",
			4730 => x"fff74aad",
			4731 => x"00042e08",
			4732 => x"09013804",
			4733 => x"00004aad",
			4734 => x"015a4aad",
			4735 => x"0c054604",
			4736 => x"00df4aad",
			4737 => x"ff314aad",
			4738 => x"05083e20",
			4739 => x"07066e10",
			4740 => x"0802e808",
			4741 => x"0c063004",
			4742 => x"ff844aad",
			4743 => x"00004aad",
			4744 => x"040c0404",
			4745 => x"00f04aad",
			4746 => x"fff44aad",
			4747 => x"030a8a0c",
			4748 => x"0b06ee04",
			4749 => x"00004aad",
			4750 => x"0d086d04",
			4751 => x"00004aad",
			4752 => x"fe504aad",
			4753 => x"00004aad",
			4754 => x"0e0a4814",
			4755 => x"0d089a04",
			4756 => x"00004aad",
			4757 => x"0c065008",
			4758 => x"00033504",
			4759 => x"00004aad",
			4760 => x"01234aad",
			4761 => x"030a8104",
			4762 => x"00004aad",
			4763 => x"000a4aad",
			4764 => x"0508a310",
			4765 => x"0e0abb08",
			4766 => x"030a8104",
			4767 => x"00004aad",
			4768 => x"feee4aad",
			4769 => x"05088604",
			4770 => x"00634aad",
			4771 => x"ff834aad",
			4772 => x"0706f508",
			4773 => x"0d093504",
			4774 => x"00004aad",
			4775 => x"00cf4aad",
			4776 => x"0901ff04",
			4777 => x"006e4aad",
			4778 => x"ff964aad",
			4779 => x"0505a00c",
			4780 => x"00067104",
			4781 => x"fea14bf9",
			4782 => x"04140204",
			4783 => x"00004bf9",
			4784 => x"fff04bf9",
			4785 => x"0f083948",
			4786 => x"06016314",
			4787 => x"0e06e208",
			4788 => x"0600e804",
			4789 => x"00004bf9",
			4790 => x"feba4bf9",
			4791 => x"0100b704",
			4792 => x"00004bf9",
			4793 => x"08021e04",
			4794 => x"00004bf9",
			4795 => x"01234bf9",
			4796 => x"02091b1c",
			4797 => x"040c0410",
			4798 => x"0b053508",
			4799 => x"0a029b04",
			4800 => x"00004bf9",
			4801 => x"fef44bf9",
			4802 => x"00044a04",
			4803 => x"00f94bf9",
			4804 => x"ffc94bf9",
			4805 => x"0c04ef08",
			4806 => x"0b051104",
			4807 => x"00004bf9",
			4808 => x"01724bf9",
			4809 => x"00004bf9",
			4810 => x"06018010",
			4811 => x"01007808",
			4812 => x"02093a04",
			4813 => x"000b4bf9",
			4814 => x"00004bf9",
			4815 => x"0900dc04",
			4816 => x"feb64bf9",
			4817 => x"00004bf9",
			4818 => x"0c04f104",
			4819 => x"01034bf9",
			4820 => x"ff6e4bf9",
			4821 => x"040b1628",
			4822 => x"06018e18",
			4823 => x"0100a608",
			4824 => x"040aed04",
			4825 => x"febb4bf9",
			4826 => x"00564bf9",
			4827 => x"05065108",
			4828 => x"0003c404",
			4829 => x"00004bf9",
			4830 => x"01684bf9",
			4831 => x"0c059c04",
			4832 => x"fe834bf9",
			4833 => x"002c4bf9",
			4834 => x"00037d04",
			4835 => x"00004bf9",
			4836 => x"0c068a08",
			4837 => x"01016004",
			4838 => x"01674bf9",
			4839 => x"00004bf9",
			4840 => x"00004bf9",
			4841 => x"06018d18",
			4842 => x"0b05560c",
			4843 => x"0d062d08",
			4844 => x"040bb204",
			4845 => x"fed74bf9",
			4846 => x"00244bf9",
			4847 => x"016d4bf9",
			4848 => x"0c04ef04",
			4849 => x"fe084bf9",
			4850 => x"01010b04",
			4851 => x"00654bf9",
			4852 => x"fdf44bf9",
			4853 => x"0b05b404",
			4854 => x"01824bf9",
			4855 => x"020ab708",
			4856 => x"06019a04",
			4857 => x"fe4f4bf9",
			4858 => x"00b04bf9",
			4859 => x"0003ee04",
			4860 => x"00a34bf9",
			4861 => x"ffcd4bf9",
			4862 => x"0306110c",
			4863 => x"06017404",
			4864 => x"fe674d3d",
			4865 => x"0704ef04",
			4866 => x"01494d3d",
			4867 => x"fe904d3d",
			4868 => x"06018a4c",
			4869 => x"07052f24",
			4870 => x"06016304",
			4871 => x"fe7f4d3d",
			4872 => x"02091110",
			4873 => x"0306a508",
			4874 => x"040c9304",
			4875 => x"ff414d3d",
			4876 => x"02624d3d",
			4877 => x"0208bb04",
			4878 => x"fffc4d3d",
			4879 => x"01bf4d3d",
			4880 => x"06017408",
			4881 => x"0900be04",
			4882 => x"01934d3d",
			4883 => x"fe5c4d3d",
			4884 => x"0f086404",
			4885 => x"01844d3d",
			4886 => x"001a4d3d",
			4887 => x"0a027b1c",
			4888 => x"0b06ee10",
			4889 => x"0e091508",
			4890 => x"0802ae04",
			4891 => x"00284d3d",
			4892 => x"ff054d3d",
			4893 => x"0a021704",
			4894 => x"03084d3d",
			4895 => x"00964d3d",
			4896 => x"0901ce08",
			4897 => x"0f0a0304",
			4898 => x"fe904d3d",
			4899 => x"014b4d3d",
			4900 => x"fe3c4d3d",
			4901 => x"0a027f04",
			4902 => x"fb904d3d",
			4903 => x"0a028004",
			4904 => x"01564d3d",
			4905 => x"fe204d3d",
			4906 => x"0508041c",
			4907 => x"040d2e10",
			4908 => x"0e089608",
			4909 => x"07054904",
			4910 => x"01b04d3d",
			4911 => x"ff2d4d3d",
			4912 => x"0802eb04",
			4913 => x"00534d3d",
			4914 => x"01aa4d3d",
			4915 => x"09010204",
			4916 => x"01bb4d3d",
			4917 => x"040dca04",
			4918 => x"00254d3d",
			4919 => x"fe284d3d",
			4920 => x"0f0ad914",
			4921 => x"07066d04",
			4922 => x"00d44d3d",
			4923 => x"0802db08",
			4924 => x"06018e04",
			4925 => x"ffb24d3d",
			4926 => x"02354d3d",
			4927 => x"0f0acb04",
			4928 => x"fe194d3d",
			4929 => x"ff554d3d",
			4930 => x"030b4110",
			4931 => x"0802e908",
			4932 => x"030b1b04",
			4933 => x"00154d3d",
			4934 => x"06444d3d",
			4935 => x"00044e04",
			4936 => x"010b4d3d",
			4937 => x"fe724d3d",
			4938 => x"0004a008",
			4939 => x"0e0b7704",
			4940 => x"feb94d3d",
			4941 => x"00c04d3d",
			4942 => x"fe674d3d",
			4943 => x"06016434",
			4944 => x"00034b24",
			4945 => x"0002dd04",
			4946 => x"fe6a4ed9",
			4947 => x"0b06cd10",
			4948 => x"0c06110c",
			4949 => x"0c056204",
			4950 => x"feb24ed9",
			4951 => x"0d078804",
			4952 => x"032e4ed9",
			4953 => x"00544ed9",
			4954 => x"05bd4ed9",
			4955 => x"02099508",
			4956 => x"0d082504",
			4957 => x"00004ed9",
			4958 => x"fe6e4ed9",
			4959 => x"0b073304",
			4960 => x"032c4ed9",
			4961 => x"fe944ed9",
			4962 => x"03069604",
			4963 => x"fe624ed9",
			4964 => x"0f082208",
			4965 => x"0f07f204",
			4966 => x"fe1e4ed9",
			4967 => x"01564ed9",
			4968 => x"fe624ed9",
			4969 => x"0c066d74",
			4970 => x"06018140",
			4971 => x"02093520",
			4972 => x"0b055610",
			4973 => x"03065908",
			4974 => x"040c9304",
			4975 => x"fe304ed9",
			4976 => x"01a44ed9",
			4977 => x"0d05f704",
			4978 => x"ff604ed9",
			4979 => x"01f34ed9",
			4980 => x"040a8808",
			4981 => x"06017404",
			4982 => x"fe914ed9",
			4983 => x"023d4ed9",
			4984 => x"0003f104",
			4985 => x"fc864ed9",
			4986 => x"ffe04ed9",
			4987 => x"03091a10",
			4988 => x"0c04ea08",
			4989 => x"02097804",
			4990 => x"00b54ed9",
			4991 => x"fdf94ed9",
			4992 => x"0f07b904",
			4993 => x"00004ed9",
			4994 => x"fe244ed9",
			4995 => x"0f097108",
			4996 => x"0e090704",
			4997 => x"009f4ed9",
			4998 => x"04954ed9",
			4999 => x"00033e04",
			5000 => x"fe594ed9",
			5001 => x"00544ed9",
			5002 => x"0802fb18",
			5003 => x"07066d0c",
			5004 => x"040b0908",
			5005 => x"00036804",
			5006 => x"fef44ed9",
			5007 => x"01f34ed9",
			5008 => x"ff914ed9",
			5009 => x"05080404",
			5010 => x"013c4ed9",
			5011 => x"0b074404",
			5012 => x"fdf64ed9",
			5013 => x"001e4ed9",
			5014 => x"0e0a3910",
			5015 => x"07054508",
			5016 => x"0d060f04",
			5017 => x"00c84ed9",
			5018 => x"02084ed9",
			5019 => x"03088d04",
			5020 => x"ff274ed9",
			5021 => x"01094ed9",
			5022 => x"06019104",
			5023 => x"04254ed9",
			5024 => x"0b072f04",
			5025 => x"01d64ed9",
			5026 => x"00b64ed9",
			5027 => x"0d095010",
			5028 => x"0c06c408",
			5029 => x"06017d04",
			5030 => x"00004ed9",
			5031 => x"fe674ed9",
			5032 => x"030af104",
			5033 => x"039d4ed9",
			5034 => x"ff6a4ed9",
			5035 => x"00039d08",
			5036 => x"0e0ac404",
			5037 => x"ff4b4ed9",
			5038 => x"11824ed9",
			5039 => x"0004a70c",
			5040 => x"040be404",
			5041 => x"fe734ed9",
			5042 => x"0a029604",
			5043 => x"03684ed9",
			5044 => x"00754ed9",
			5045 => x"fe624ed9",
			5046 => x"0601643c",
			5047 => x"0901a120",
			5048 => x"0100a10c",
			5049 => x"03069604",
			5050 => x"fe635075",
			5051 => x"0306a504",
			5052 => x"00915075",
			5053 => x"fe7d5075",
			5054 => x"0705ff10",
			5055 => x"0c056204",
			5056 => x"fe895075",
			5057 => x"0002f604",
			5058 => x"febe5075",
			5059 => x"0003d804",
			5060 => x"03165075",
			5061 => x"ff905075",
			5062 => x"fe5d5075",
			5063 => x"0a020808",
			5064 => x"0b06cd04",
			5065 => x"049f5075",
			5066 => x"ff875075",
			5067 => x"0b06bc04",
			5068 => x"fe895075",
			5069 => x"01011b0c",
			5070 => x"07064604",
			5071 => x"01845075",
			5072 => x"01010604",
			5073 => x"00f35075",
			5074 => x"fe7b5075",
			5075 => x"02b55075",
			5076 => x"0b077168",
			5077 => x"06018138",
			5078 => x"0b055618",
			5079 => x"0f088b10",
			5080 => x"0306c508",
			5081 => x"0f082b04",
			5082 => x"01035075",
			5083 => x"fe245075",
			5084 => x"040ad504",
			5085 => x"017a5075",
			5086 => x"02425075",
			5087 => x"03073b04",
			5088 => x"fdc05075",
			5089 => x"00c15075",
			5090 => x"040a9510",
			5091 => x"0a025408",
			5092 => x"0f097d04",
			5093 => x"014e5075",
			5094 => x"ff4f5075",
			5095 => x"0100b704",
			5096 => x"01065075",
			5097 => x"03535075",
			5098 => x"0b068d08",
			5099 => x"0003ee04",
			5100 => x"fd825075",
			5101 => x"ff3f5075",
			5102 => x"01011f04",
			5103 => x"016b5075",
			5104 => x"fece5075",
			5105 => x"0e0a9a20",
			5106 => x"05080410",
			5107 => x"0e09e008",
			5108 => x"07054504",
			5109 => x"01c15075",
			5110 => x"00525075",
			5111 => x"09021d04",
			5112 => x"01d05075",
			5113 => x"00c45075",
			5114 => x"07066d08",
			5115 => x"040ab204",
			5116 => x"00215075",
			5117 => x"018c5075",
			5118 => x"030a6904",
			5119 => x"fe445075",
			5120 => x"00125075",
			5121 => x"06019204",
			5122 => x"07965075",
			5123 => x"05089408",
			5124 => x"0c063a04",
			5125 => x"01d15075",
			5126 => x"00545075",
			5127 => x"fe9c5075",
			5128 => x"0004a028",
			5129 => x"0901fe14",
			5130 => x"0601af0c",
			5131 => x"0901e808",
			5132 => x"0508dd04",
			5133 => x"00005075",
			5134 => x"025a5075",
			5135 => x"04cf5075",
			5136 => x"01011f04",
			5137 => x"01595075",
			5138 => x"feb45075",
			5139 => x"040d0010",
			5140 => x"0b07b808",
			5141 => x"0c06ac04",
			5142 => x"fe645075",
			5143 => x"00735075",
			5144 => x"00039a04",
			5145 => x"05725075",
			5146 => x"fe745075",
			5147 => x"018c5075",
			5148 => x"fe645075",
			5149 => x"040a5b40",
			5150 => x"0c05f824",
			5151 => x"07063f18",
			5152 => x"0100b404",
			5153 => x"00005209",
			5154 => x"0101130c",
			5155 => x"08021e04",
			5156 => x"00005209",
			5157 => x"0c05f704",
			5158 => x"00b05209",
			5159 => x"00005209",
			5160 => x"0e092404",
			5161 => x"ffd75209",
			5162 => x"00005209",
			5163 => x"0209b704",
			5164 => x"ff3b5209",
			5165 => x"0802b704",
			5166 => x"003d5209",
			5167 => x"00005209",
			5168 => x"07067018",
			5169 => x"0802aa10",
			5170 => x"04091d04",
			5171 => x"00005209",
			5172 => x"0b06de08",
			5173 => x"0002dd04",
			5174 => x"00005209",
			5175 => x"00e55209",
			5176 => x"00005209",
			5177 => x"0802c304",
			5178 => x"ffe55209",
			5179 => x"00115209",
			5180 => x"00005209",
			5181 => x"00043a3c",
			5182 => x"08036338",
			5183 => x"030a691c",
			5184 => x"0c050710",
			5185 => x"01009508",
			5186 => x"0b055404",
			5187 => x"00005209",
			5188 => x"fec15209",
			5189 => x"00042d04",
			5190 => x"00bd5209",
			5191 => x"ffc05209",
			5192 => x"0100e704",
			5193 => x"fe985209",
			5194 => x"07066d04",
			5195 => x"00165209",
			5196 => x"ff225209",
			5197 => x"01013f0c",
			5198 => x"0c05f504",
			5199 => x"00005209",
			5200 => x"0a02a804",
			5201 => x"00c05209",
			5202 => x"00005209",
			5203 => x"0a026c08",
			5204 => x"0c068d04",
			5205 => x"008f5209",
			5206 => x"00005209",
			5207 => x"0c063a04",
			5208 => x"00005209",
			5209 => x"ff3a5209",
			5210 => x"feee5209",
			5211 => x"00045b20",
			5212 => x"0508fb1c",
			5213 => x"040bbf10",
			5214 => x"00044708",
			5215 => x"08035e04",
			5216 => x"00005209",
			5217 => x"00545209",
			5218 => x"00045404",
			5219 => x"ff735209",
			5220 => x"00005209",
			5221 => x"0900cd04",
			5222 => x"00005209",
			5223 => x"0c061404",
			5224 => x"01625209",
			5225 => x"00005209",
			5226 => x"ff7d5209",
			5227 => x"0a02db14",
			5228 => x"0100800c",
			5229 => x"0505cc04",
			5230 => x"ffbf5209",
			5231 => x"02092004",
			5232 => x"00ad5209",
			5233 => x"00005209",
			5234 => x"040be404",
			5235 => x"00005209",
			5236 => x"fefa5209",
			5237 => x"0803e610",
			5238 => x"0c051108",
			5239 => x"01007e04",
			5240 => x"00005209",
			5241 => x"01105209",
			5242 => x"030bfd04",
			5243 => x"ff8b5209",
			5244 => x"00835209",
			5245 => x"040f0204",
			5246 => x"ff035209",
			5247 => x"05058404",
			5248 => x"00005209",
			5249 => x"00345209",
			5250 => x"06016334",
			5251 => x"0100fa14",
			5252 => x"0600e808",
			5253 => x"00030204",
			5254 => x"ffcb53df",
			5255 => x"005953df",
			5256 => x"04085208",
			5257 => x"08021e04",
			5258 => x"ff2653df",
			5259 => x"00b453df",
			5260 => x"fe6a53df",
			5261 => x"03097818",
			5262 => x"0c060f10",
			5263 => x"04098704",
			5264 => x"fec353df",
			5265 => x"0a021704",
			5266 => x"01cc53df",
			5267 => x"0e087804",
			5268 => x"006653df",
			5269 => x"ff2e53df",
			5270 => x"0901a904",
			5271 => x"ffe653df",
			5272 => x"02ae53df",
			5273 => x"0100fc04",
			5274 => x"006353df",
			5275 => x"fe6353df",
			5276 => x"06018d70",
			5277 => x"0f08723c",
			5278 => x"0306691c",
			5279 => x"0c04b20c",
			5280 => x"0704d404",
			5281 => x"feb053df",
			5282 => x"040c2c04",
			5283 => x"ffb253df",
			5284 => x"022053df",
			5285 => x"0e05ce08",
			5286 => x"0d05e904",
			5287 => x"fe9653df",
			5288 => x"008b53df",
			5289 => x"0e060f04",
			5290 => x"fda153df",
			5291 => x"ff5553df",
			5292 => x"00042010",
			5293 => x"0306b908",
			5294 => x"00040304",
			5295 => x"fec353df",
			5296 => x"fce953df",
			5297 => x"0c04d204",
			5298 => x"022d53df",
			5299 => x"ffd953df",
			5300 => x"07050808",
			5301 => x"0f07fe04",
			5302 => x"02b553df",
			5303 => x"018d53df",
			5304 => x"06017404",
			5305 => x"feda53df",
			5306 => x"018953df",
			5307 => x"040b3c14",
			5308 => x"00040310",
			5309 => x"0100aa08",
			5310 => x"0e075804",
			5311 => x"fb6553df",
			5312 => x"fe5753df",
			5313 => x"05065104",
			5314 => x"019553df",
			5315 => x"ffe153df",
			5316 => x"01a953df",
			5317 => x"040bb210",
			5318 => x"06018908",
			5319 => x"00042004",
			5320 => x"fda753df",
			5321 => x"fff653df",
			5322 => x"0f0afc04",
			5323 => x"fb6a53df",
			5324 => x"ff9f53df",
			5325 => x"06017808",
			5326 => x"0003ed04",
			5327 => x"003f53df",
			5328 => x"fe2c53df",
			5329 => x"0900ef04",
			5330 => x"fee953df",
			5331 => x"009c53df",
			5332 => x"0d087f20",
			5333 => x"08034c0c",
			5334 => x"00039504",
			5335 => x"ff3d53df",
			5336 => x"040c0404",
			5337 => x"01a853df",
			5338 => x"000053df",
			5339 => x"07054b08",
			5340 => x"09014d04",
			5341 => x"01d753df",
			5342 => x"007853df",
			5343 => x"09015804",
			5344 => x"fd5b53df",
			5345 => x"0705ea04",
			5346 => x"01a653df",
			5347 => x"ff3f53df",
			5348 => x"0f0adf0c",
			5349 => x"0f0a9208",
			5350 => x"0f0a8a04",
			5351 => x"ffb953df",
			5352 => x"007553df",
			5353 => x"fe5253df",
			5354 => x"00039d0c",
			5355 => x"0f0aed04",
			5356 => x"ffa753df",
			5357 => x"07070c04",
			5358 => x"02b153df",
			5359 => x"004153df",
			5360 => x"030ae108",
			5361 => x"030aa904",
			5362 => x"ff3453df",
			5363 => x"01c353df",
			5364 => x"0d090104",
			5365 => x"011c53df",
			5366 => x"ff4553df",
			5367 => x"03063a24",
			5368 => x"0a02ed08",
			5369 => x"0b059904",
			5370 => x"fe7054c1",
			5371 => x"000054c1",
			5372 => x"0a03230c",
			5373 => x"0505af04",
			5374 => x"ff7c54c1",
			5375 => x"06017804",
			5376 => x"000054c1",
			5377 => x"013754c1",
			5378 => x"0209ab04",
			5379 => x"fe8254c1",
			5380 => x"0209c908",
			5381 => x"0e03a604",
			5382 => x"000054c1",
			5383 => x"00b154c1",
			5384 => x"000054c1",
			5385 => x"0f07eb18",
			5386 => x"0900cf08",
			5387 => x"08036e04",
			5388 => x"000054c1",
			5389 => x"022354c1",
			5390 => x"03065904",
			5391 => x"feac54c1",
			5392 => x"00028d04",
			5393 => x"000054c1",
			5394 => x"0704ed04",
			5395 => x"000054c1",
			5396 => x"017554c1",
			5397 => x"0505db10",
			5398 => x"0f08220c",
			5399 => x"03067808",
			5400 => x"0e061e04",
			5401 => x"fe9454c1",
			5402 => x"000054c1",
			5403 => x"013054c1",
			5404 => x"fe2d54c1",
			5405 => x"0704f10c",
			5406 => x"0003f204",
			5407 => x"fedf54c1",
			5408 => x"0d060f04",
			5409 => x"000054c1",
			5410 => x"01ef54c1",
			5411 => x"0d061d10",
			5412 => x"00045808",
			5413 => x"0208e904",
			5414 => x"000054c1",
			5415 => x"fd2b54c1",
			5416 => x"0a02c604",
			5417 => x"ff3754c1",
			5418 => x"006254c1",
			5419 => x"0803e608",
			5420 => x"05061504",
			5421 => x"00bb54c1",
			5422 => x"001154c1",
			5423 => x"fe4e54c1",
			5424 => x"03063a24",
			5425 => x"040e6308",
			5426 => x"0d066b04",
			5427 => x"fe8255c5",
			5428 => x"000055c5",
			5429 => x"0305a010",
			5430 => x"0209ab04",
			5431 => x"febf55c5",
			5432 => x"0209b108",
			5433 => x"0b060904",
			5434 => x"005355c5",
			5435 => x"000055c5",
			5436 => x"000055c5",
			5437 => x"04116208",
			5438 => x"07051a04",
			5439 => x"011055c5",
			5440 => x"000055c5",
			5441 => x"000055c5",
			5442 => x"0f07eb1c",
			5443 => x"01007d08",
			5444 => x"08036e04",
			5445 => x"000055c5",
			5446 => x"021855c5",
			5447 => x"0d060f04",
			5448 => x"fed155c5",
			5449 => x"0f078104",
			5450 => x"000055c5",
			5451 => x"0c04d104",
			5452 => x"000055c5",
			5453 => x"0e061e04",
			5454 => x"000855c5",
			5455 => x"019555c5",
			5456 => x"0d060f10",
			5457 => x"0f082208",
			5458 => x"06017004",
			5459 => x"fea255c5",
			5460 => x"008955c5",
			5461 => x"0306b904",
			5462 => x"fddc55c5",
			5463 => x"ffae55c5",
			5464 => x"0f084618",
			5465 => x"07050808",
			5466 => x"0306a504",
			5467 => x"007055c5",
			5468 => x"021855c5",
			5469 => x"0306ff08",
			5470 => x"08037c04",
			5471 => x"fe9e55c5",
			5472 => x"00f255c5",
			5473 => x"06015b04",
			5474 => x"000055c5",
			5475 => x"016c55c5",
			5476 => x"0100a810",
			5477 => x"0003f308",
			5478 => x"0d064504",
			5479 => x"fd6055c5",
			5480 => x"ff0555c5",
			5481 => x"0f08e604",
			5482 => x"004855c5",
			5483 => x"fe2055c5",
			5484 => x"0b058304",
			5485 => x"018d55c5",
			5486 => x"0100ef04",
			5487 => x"ff5155c5",
			5488 => x"004355c5",
			5489 => x"07050434",
			5490 => x"0e06ac28",
			5491 => x"0306b920",
			5492 => x"040c5808",
			5493 => x"0d061104",
			5494 => x"fedd56c9",
			5495 => x"000056c9",
			5496 => x"02091910",
			5497 => x"0b051408",
			5498 => x"02091104",
			5499 => x"ffbb56c9",
			5500 => x"000056c9",
			5501 => x"0c04d404",
			5502 => x"014856c9",
			5503 => x"000056c9",
			5504 => x"06017c04",
			5505 => x"fefa56c9",
			5506 => x"000056c9",
			5507 => x"0900e704",
			5508 => x"000056c9",
			5509 => x"015d56c9",
			5510 => x"03071b08",
			5511 => x"06017804",
			5512 => x"000056c9",
			5513 => x"fe3456c9",
			5514 => x"00f756c9",
			5515 => x"07050814",
			5516 => x"0c04e70c",
			5517 => x"06016304",
			5518 => x"000056c9",
			5519 => x"0d05e904",
			5520 => x"000056c9",
			5521 => x"018d56c9",
			5522 => x"07050604",
			5523 => x"ff7656c9",
			5524 => x"008656c9",
			5525 => x"0d061d08",
			5526 => x"040e6304",
			5527 => x"feac56c9",
			5528 => x"000056c9",
			5529 => x"0b058318",
			5530 => x"06017408",
			5531 => x"0900d904",
			5532 => x"000056c9",
			5533 => x"fe9356c9",
			5534 => x"00042008",
			5535 => x"01009d04",
			5536 => x"ff9756c9",
			5537 => x"012d56c9",
			5538 => x"07054504",
			5539 => x"01a856c9",
			5540 => x"000056c9",
			5541 => x"07055f0c",
			5542 => x"06019208",
			5543 => x"07051f04",
			5544 => x"000056c9",
			5545 => x"fe6b56c9",
			5546 => x"002d56c9",
			5547 => x"0003f308",
			5548 => x"03097804",
			5549 => x"008c56c9",
			5550 => x"000e56c9",
			5551 => x"0a02a104",
			5552 => x"fe6856c9",
			5553 => x"000056c9",
			5554 => x"03063a18",
			5555 => x"0a02ed08",
			5556 => x"01009f04",
			5557 => x"fe6d5795",
			5558 => x"00005795",
			5559 => x"0705180c",
			5560 => x"0b050408",
			5561 => x"0b04ce04",
			5562 => x"feae5795",
			5563 => x"00005795",
			5564 => x"016a5795",
			5565 => x"fe575795",
			5566 => x"0005084c",
			5567 => x"0004251c",
			5568 => x"0306b908",
			5569 => x"00041c04",
			5570 => x"fe5f5795",
			5571 => x"fb455795",
			5572 => x"0505f604",
			5573 => x"025e5795",
			5574 => x"0100a608",
			5575 => x"0100a304",
			5576 => x"ffb45795",
			5577 => x"fbdd5795",
			5578 => x"05065104",
			5579 => x"017d5795",
			5580 => x"001c5795",
			5581 => x"00046c10",
			5582 => x"0a02a504",
			5583 => x"fec55795",
			5584 => x"0c068b08",
			5585 => x"0900f304",
			5586 => x"009c5795",
			5587 => x"01695795",
			5588 => x"fedf5795",
			5589 => x"0a02db10",
			5590 => x"0f087208",
			5591 => x"0a02c304",
			5592 => x"fe9d5795",
			5593 => x"00b65795",
			5594 => x"00047904",
			5595 => x"000d5795",
			5596 => x"fe405795",
			5597 => x"0c054608",
			5598 => x"040e6304",
			5599 => x"016e5795",
			5600 => x"ffc95795",
			5601 => x"0b07d604",
			5602 => x"fe715795",
			5603 => x"014a5795",
			5604 => x"fe165795",
			5605 => x"03063a1c",
			5606 => x"06017008",
			5607 => x"01009f04",
			5608 => x"fe7958a9",
			5609 => x"000058a9",
			5610 => x"0e05ac10",
			5611 => x"0305c008",
			5612 => x"02093d04",
			5613 => x"fef258a9",
			5614 => x"000058a9",
			5615 => x"0b053304",
			5616 => x"014a58a9",
			5617 => x"000058a9",
			5618 => x"fe3f58a9",
			5619 => x"0f084634",
			5620 => x"0705081c",
			5621 => x"0d05f70c",
			5622 => x"0f07d508",
			5623 => x"040adc04",
			5624 => x"000058a9",
			5625 => x"00fc58a9",
			5626 => x"fef158a9",
			5627 => x"0208ad04",
			5628 => x"ff4358a9",
			5629 => x"0e05e904",
			5630 => x"001958a9",
			5631 => x"06016304",
			5632 => x"000058a9",
			5633 => x"019658a9",
			5634 => x"0306a508",
			5635 => x"040ceb04",
			5636 => x"fe9b58a9",
			5637 => x"000058a9",
			5638 => x"0506f10c",
			5639 => x"0f083908",
			5640 => x"0f078104",
			5641 => x"000058a9",
			5642 => x"011e58a9",
			5643 => x"000058a9",
			5644 => x"ff0d58a9",
			5645 => x"03076c20",
			5646 => x"0e073b1c",
			5647 => x"0705040c",
			5648 => x"03071b08",
			5649 => x"040bb204",
			5650 => x"fddd58a9",
			5651 => x"ff7c58a9",
			5652 => x"012558a9",
			5653 => x"0c04ec08",
			5654 => x"06017404",
			5655 => x"ffbd58a9",
			5656 => x"01a358a9",
			5657 => x"06018104",
			5658 => x"ff0558a9",
			5659 => x"010958a9",
			5660 => x"fdcf58a9",
			5661 => x"0d0a2b18",
			5662 => x"0b058308",
			5663 => x"06018004",
			5664 => x"000058a9",
			5665 => x"019258a9",
			5666 => x"03087508",
			5667 => x"05065104",
			5668 => x"002c58a9",
			5669 => x"fece58a9",
			5670 => x"0705a104",
			5671 => x"01d458a9",
			5672 => x"004258a9",
			5673 => x"fe6258a9",
			5674 => x"06015f2c",
			5675 => x"01010214",
			5676 => x"08027910",
			5677 => x"0506f10c",
			5678 => x"07059104",
			5679 => x"fec559a5",
			5680 => x"0801e404",
			5681 => x"000059a5",
			5682 => x"01d659a5",
			5683 => x"fe7e59a5",
			5684 => x"fe6659a5",
			5685 => x"03097814",
			5686 => x"02094d10",
			5687 => x"0101210c",
			5688 => x"0a020004",
			5689 => x"010659a5",
			5690 => x"0d081704",
			5691 => x"004259a5",
			5692 => x"feb259a5",
			5693 => x"01e659a5",
			5694 => x"033859a5",
			5695 => x"fef459a5",
			5696 => x"0a033e4c",
			5697 => x"06019a2c",
			5698 => x"040a8818",
			5699 => x"0c06140c",
			5700 => x"09010f04",
			5701 => x"fede59a5",
			5702 => x"0901b804",
			5703 => x"01dc59a5",
			5704 => x"00a259a5",
			5705 => x"08029e08",
			5706 => x"02098104",
			5707 => x"ffe959a5",
			5708 => x"01eb59a5",
			5709 => x"fe6e59a5",
			5710 => x"06016704",
			5711 => x"fe5b59a5",
			5712 => x"0f082b08",
			5713 => x"07051f04",
			5714 => x"010c59a5",
			5715 => x"fdef59a5",
			5716 => x"0306c504",
			5717 => x"fe6259a5",
			5718 => x"001959a5",
			5719 => x"07068810",
			5720 => x"040d2e0c",
			5721 => x"09015804",
			5722 => x"003459a5",
			5723 => x"08030804",
			5724 => x"007459a5",
			5725 => x"019e59a5",
			5726 => x"000059a5",
			5727 => x"0e0c7e0c",
			5728 => x"09023b08",
			5729 => x"0f0b4404",
			5730 => x"ff2259a5",
			5731 => x"010159a5",
			5732 => x"fe3559a5",
			5733 => x"017959a5",
			5734 => x"0505f604",
			5735 => x"006c59a5",
			5736 => x"fe4559a5",
			5737 => x"0705052c",
			5738 => x"06017920",
			5739 => x"0e06ac18",
			5740 => x"0d05f704",
			5741 => x"ff535ad9",
			5742 => x"0c04cf08",
			5743 => x"06017404",
			5744 => x"ff9d5ad9",
			5745 => x"00005ad9",
			5746 => x"02092408",
			5747 => x"06016304",
			5748 => x"00005ad9",
			5749 => x"00d45ad9",
			5750 => x"00005ad9",
			5751 => x"08033704",
			5752 => x"00005ad9",
			5753 => x"fec35ad9",
			5754 => x"0d061f08",
			5755 => x"0704ee04",
			5756 => x"002f5ad9",
			5757 => x"ff8a5ad9",
			5758 => x"00bb5ad9",
			5759 => x"02096028",
			5760 => x"06017018",
			5761 => x"0c056208",
			5762 => x"0b053304",
			5763 => x"00005ad9",
			5764 => x"ff5d5ad9",
			5765 => x"0b06d20c",
			5766 => x"0e06e204",
			5767 => x"00005ad9",
			5768 => x"01013004",
			5769 => x"00795ad9",
			5770 => x"00005ad9",
			5771 => x"00005ad9",
			5772 => x"0a024904",
			5773 => x"00005ad9",
			5774 => x"0d060304",
			5775 => x"00005ad9",
			5776 => x"0e065a04",
			5777 => x"00005ad9",
			5778 => x"010b5ad9",
			5779 => x"0b073324",
			5780 => x"0803901c",
			5781 => x"020ad910",
			5782 => x"00043108",
			5783 => x"0100e704",
			5784 => x"ff3c5ad9",
			5785 => x"001c5ad9",
			5786 => x"07057704",
			5787 => x"00e05ad9",
			5788 => x"ffe95ad9",
			5789 => x"0f0b9808",
			5790 => x"0c063304",
			5791 => x"012a5ad9",
			5792 => x"00005ad9",
			5793 => x"00005ad9",
			5794 => x"0100b404",
			5795 => x"00005ad9",
			5796 => x"ff205ad9",
			5797 => x"0e0cac1c",
			5798 => x"01012e0c",
			5799 => x"0706b404",
			5800 => x"ffe25ad9",
			5801 => x"0e09fd04",
			5802 => x"00005ad9",
			5803 => x"00615ad9",
			5804 => x"06018e08",
			5805 => x"00039a04",
			5806 => x"00005ad9",
			5807 => x"002e5ad9",
			5808 => x"00039504",
			5809 => x"00005ad9",
			5810 => x"ff075ad9",
			5811 => x"0601ec04",
			5812 => x"00c45ad9",
			5813 => x"00005ad9",
			5814 => x"0505db24",
			5815 => x"040c930c",
			5816 => x"07050804",
			5817 => x"fe5f5c0d",
			5818 => x"07051804",
			5819 => x"00005c0d",
			5820 => x"ff815c0d",
			5821 => x"0d05a804",
			5822 => x"fea85c0d",
			5823 => x"0c04b208",
			5824 => x"06016704",
			5825 => x"00005c0d",
			5826 => x"01775c0d",
			5827 => x"06017808",
			5828 => x"040d2e04",
			5829 => x"fed55c0d",
			5830 => x"00005c0d",
			5831 => x"01165c0d",
			5832 => x"0505f620",
			5833 => x"0d060f14",
			5834 => x"00042404",
			5835 => x"feb35c0d",
			5836 => x"02091908",
			5837 => x"06016404",
			5838 => x"00005c0d",
			5839 => x"01785c0d",
			5840 => x"0900d604",
			5841 => x"00005c0d",
			5842 => x"ff155c0d",
			5843 => x"06016304",
			5844 => x"00005c0d",
			5845 => x"07051c04",
			5846 => x"01985c0d",
			5847 => x"00005c0d",
			5848 => x"0d061f1c",
			5849 => x"040cc610",
			5850 => x"0704f104",
			5851 => x"ff455c0d",
			5852 => x"01008004",
			5853 => x"00005c0d",
			5854 => x"00041c04",
			5855 => x"00005c0d",
			5856 => x"fdb65c0d",
			5857 => x"02098108",
			5858 => x"0c052804",
			5859 => x"010e5c0d",
			5860 => x"00005c0d",
			5861 => x"00005c0d",
			5862 => x"0209111c",
			5863 => x"0a029010",
			5864 => x"03073b08",
			5865 => x"040a5b04",
			5866 => x"00005c0d",
			5867 => x"fee65c0d",
			5868 => x"0100b404",
			5869 => x"fffe5c0d",
			5870 => x"01125c0d",
			5871 => x"0c050708",
			5872 => x"05061904",
			5873 => x"01dc5c0d",
			5874 => x"00005c0d",
			5875 => x"ffa65c0d",
			5876 => x"0e06ce10",
			5877 => x"06017908",
			5878 => x"0e061e04",
			5879 => x"00005c0d",
			5880 => x"fdab5c0d",
			5881 => x"0d065d04",
			5882 => x"018f5c0d",
			5883 => x"fed95c0d",
			5884 => x"0d0a1e08",
			5885 => x"030a9904",
			5886 => x"00015c0d",
			5887 => x"00995c0d",
			5888 => x"0c071e04",
			5889 => x"fe425c0d",
			5890 => x"00005c0d",
			5891 => x"03073b54",
			5892 => x"0a029220",
			5893 => x"0f082b14",
			5894 => x"0e068d08",
			5895 => x"0600e804",
			5896 => x"00005d69",
			5897 => x"ff365d69",
			5898 => x"01009b04",
			5899 => x"00005d69",
			5900 => x"0801e404",
			5901 => x"00005d69",
			5902 => x"00645d69",
			5903 => x"0c04b904",
			5904 => x"00005d69",
			5905 => x"0d065204",
			5906 => x"fe145d69",
			5907 => x"00005d69",
			5908 => x"040b2908",
			5909 => x"0306b904",
			5910 => x"00005d69",
			5911 => x"011b5d69",
			5912 => x"040b9d10",
			5913 => x"0704d704",
			5914 => x"00005d69",
			5915 => x"01009708",
			5916 => x"0c04b104",
			5917 => x"00005d69",
			5918 => x"febe5d69",
			5919 => x"00005d69",
			5920 => x"06017410",
			5921 => x"0208fe08",
			5922 => x"03063a04",
			5923 => x"ff5e5d69",
			5924 => x"00fc5d69",
			5925 => x"0704d504",
			5926 => x"00005d69",
			5927 => x"fea35d69",
			5928 => x"0d065208",
			5929 => x"0209ce04",
			5930 => x"00e45d69",
			5931 => x"ffda5d69",
			5932 => x"ff095d69",
			5933 => x"0f091520",
			5934 => x"0d080b1c",
			5935 => x"040bbd14",
			5936 => x"0100a308",
			5937 => x"0c04ed04",
			5938 => x"00005d69",
			5939 => x"fff15d69",
			5940 => x"0901b208",
			5941 => x"08021e04",
			5942 => x"00005d69",
			5943 => x"00ff5d69",
			5944 => x"00005d69",
			5945 => x"07053404",
			5946 => x"00075d69",
			5947 => x"ffee5d69",
			5948 => x"00005d69",
			5949 => x"09014b10",
			5950 => x"020a6b08",
			5951 => x"0d069e04",
			5952 => x"00005d69",
			5953 => x"fe7f5d69",
			5954 => x"00049c04",
			5955 => x"00ce5d69",
			5956 => x"00005d69",
			5957 => x"0d07960c",
			5958 => x"0c050c04",
			5959 => x"00005d69",
			5960 => x"0209ef04",
			5961 => x"00005d69",
			5962 => x"01415d69",
			5963 => x"01012510",
			5964 => x"0f0aed08",
			5965 => x"06018304",
			5966 => x"00005d69",
			5967 => x"fe4e5d69",
			5968 => x"00043504",
			5969 => x"00745d69",
			5970 => x"00005d69",
			5971 => x"040b8a08",
			5972 => x"0a025704",
			5973 => x"00005d69",
			5974 => x"008c5d69",
			5975 => x"0f0b2604",
			5976 => x"ff045d69",
			5977 => x"00155d69",
			5978 => x"0306ff40",
			5979 => x"0b055634",
			5980 => x"00042414",
			5981 => x"0d061f0c",
			5982 => x"08032604",
			5983 => x"00005e9d",
			5984 => x"040b8004",
			5985 => x"fe985e9d",
			5986 => x"00005e9d",
			5987 => x"040af504",
			5988 => x"00005e9d",
			5989 => x"00605e9d",
			5990 => x"0f088b1c",
			5991 => x"03067810",
			5992 => x"040c5e08",
			5993 => x"03065904",
			5994 => x"fecb5e9d",
			5995 => x"00005e9d",
			5996 => x"0b053304",
			5997 => x"00745e9d",
			5998 => x"ffc35e9d",
			5999 => x"02092404",
			6000 => x"01735e9d",
			6001 => x"0306c504",
			6002 => x"ffbb5e9d",
			6003 => x"00fc5e9d",
			6004 => x"feca5e9d",
			6005 => x"0f082204",
			6006 => x"00005e9d",
			6007 => x"02098e04",
			6008 => x"fdef5e9d",
			6009 => x"00005e9d",
			6010 => x"0506260c",
			6011 => x"01009504",
			6012 => x"ff425e9d",
			6013 => x"0003d104",
			6014 => x"00005e9d",
			6015 => x"01795e9d",
			6016 => x"0b05c71c",
			6017 => x"06018d14",
			6018 => x"07051a08",
			6019 => x"0b056504",
			6020 => x"fff45e9d",
			6021 => x"00005e9d",
			6022 => x"00044608",
			6023 => x"0100d204",
			6024 => x"fe835e9d",
			6025 => x"00005e9d",
			6026 => x"00005e9d",
			6027 => x"0b05b404",
			6028 => x"01035e9d",
			6029 => x"ff605e9d",
			6030 => x"0b060b14",
			6031 => x"07057508",
			6032 => x"020a6304",
			6033 => x"ffca5e9d",
			6034 => x"00105e9d",
			6035 => x"03075404",
			6036 => x"00005e9d",
			6037 => x"040da904",
			6038 => x"01705e9d",
			6039 => x"00005e9d",
			6040 => x"0003ee10",
			6041 => x"0f095608",
			6042 => x"0506f104",
			6043 => x"00005e9d",
			6044 => x"ff795e9d",
			6045 => x"07062a04",
			6046 => x"00005e9d",
			6047 => x"006b5e9d",
			6048 => x"08032b08",
			6049 => x"030a9904",
			6050 => x"fe465e9d",
			6051 => x"00005e9d",
			6052 => x"020cab04",
			6053 => x"ffe75e9d",
			6054 => x"00cf5e9d",
			6055 => x"0b051418",
			6056 => x"02093d10",
			6057 => x"0505bd04",
			6058 => x"fe695f99",
			6059 => x"0b051204",
			6060 => x"ff435f99",
			6061 => x"0505bf04",
			6062 => x"00035f99",
			6063 => x"00005f99",
			6064 => x"0803e604",
			6065 => x"fee65f99",
			6066 => x"016f5f99",
			6067 => x"0a033e60",
			6068 => x"06018d38",
			6069 => x"0c04cc18",
			6070 => x"0601700c",
			6071 => x"0f07eb08",
			6072 => x"0a02a604",
			6073 => x"feeb5f99",
			6074 => x"01c85f99",
			6075 => x"fe455f99",
			6076 => x"02093504",
			6077 => x"01d85f99",
			6078 => x"0d061f04",
			6079 => x"feda5f99",
			6080 => x"01a45f99",
			6081 => x"03066910",
			6082 => x"0b052408",
			6083 => x"06016b04",
			6084 => x"fef35f99",
			6085 => x"01205f99",
			6086 => x"0803c704",
			6087 => x"fe1a5f99",
			6088 => x"003a5f99",
			6089 => x"0e064308",
			6090 => x"0b055604",
			6091 => x"01fa5f99",
			6092 => x"fee95f99",
			6093 => x"0306b904",
			6094 => x"fe795f99",
			6095 => x"ffea5f99",
			6096 => x"0d086510",
			6097 => x"08034c04",
			6098 => x"01a05f99",
			6099 => x"0b05b404",
			6100 => x"01b85f99",
			6101 => x"0100ca04",
			6102 => x"fe445f99",
			6103 => x"00b45f99",
			6104 => x"0f0adf0c",
			6105 => x"0b06ff04",
			6106 => x"00795f99",
			6107 => x"0e0a1b04",
			6108 => x"00005f99",
			6109 => x"fe695f99",
			6110 => x"0c05f004",
			6111 => x"feaf5f99",
			6112 => x"0b073304",
			6113 => x"01725f99",
			6114 => x"00245f99",
			6115 => x"0c04ea04",
			6116 => x"00005f99",
			6117 => x"fe5e5f99",
			6118 => x"0d05e914",
			6119 => x"040df504",
			6120 => x"fe7860b5",
			6121 => x"00051508",
			6122 => x"0a02e404",
			6123 => x"000060b5",
			6124 => x"005460b5",
			6125 => x"02098e04",
			6126 => x"ff3560b5",
			6127 => x"000060b5",
			6128 => x"040b8330",
			6129 => x"0100920c",
			6130 => x"040b4a04",
			6131 => x"fe2d60b5",
			6132 => x"0505ea04",
			6133 => x"000060b5",
			6134 => x"002960b5",
			6135 => x"0c04d008",
			6136 => x"0306ff04",
			6137 => x"000060b5",
			6138 => x"019260b5",
			6139 => x"0c05f80c",
			6140 => x"0704f104",
			6141 => x"01a560b5",
			6142 => x"05080104",
			6143 => x"001460b5",
			6144 => x"fec160b5",
			6145 => x"0901a908",
			6146 => x"0706ca04",
			6147 => x"fee360b5",
			6148 => x"006660b5",
			6149 => x"09020a04",
			6150 => x"010a60b5",
			6151 => x"004760b5",
			6152 => x"07058d18",
			6153 => x"0a02a904",
			6154 => x"fe6760b5",
			6155 => x"03087510",
			6156 => x"02096008",
			6157 => x"0306e204",
			6158 => x"004b60b5",
			6159 => x"01d860b5",
			6160 => x"0a02db04",
			6161 => x"ff3560b5",
			6162 => x"005260b5",
			6163 => x"01b760b5",
			6164 => x"020adf14",
			6165 => x"0a02bc0c",
			6166 => x"040c4404",
			6167 => x"fddd60b5",
			6168 => x"0a027a04",
			6169 => x"002460b5",
			6170 => x"000060b5",
			6171 => x"040d0e04",
			6172 => x"004460b5",
			6173 => x"ffbf60b5",
			6174 => x"08037310",
			6175 => x"0c065208",
			6176 => x"0a029204",
			6177 => x"000060b5",
			6178 => x"013860b5",
			6179 => x"0508f804",
			6180 => x"fef960b5",
			6181 => x"009b60b5",
			6182 => x"0e0cbb08",
			6183 => x"020bbc04",
			6184 => x"ffc760b5",
			6185 => x"fe1860b5",
			6186 => x"0d0a1104",
			6187 => x"00ff60b5",
			6188 => x"ff8760b5",
			6189 => x"0b051418",
			6190 => x"02093d10",
			6191 => x"0505bd04",
			6192 => x"fe6761b9",
			6193 => x"0b051204",
			6194 => x"ff3a61b9",
			6195 => x"0505bf04",
			6196 => x"000361b9",
			6197 => x"000061b9",
			6198 => x"0803e604",
			6199 => x"fedc61b9",
			6200 => x"018e61b9",
			6201 => x"0a033e64",
			6202 => x"06018d34",
			6203 => x"0c04cc18",
			6204 => x"040bb20c",
			6205 => x"01009708",
			6206 => x"0f084604",
			6207 => x"ffc161b9",
			6208 => x"fcca61b9",
			6209 => x"018361b9",
			6210 => x"0505cc08",
			6211 => x"0f07b204",
			6212 => x"019b61b9",
			6213 => x"fe8a61b9",
			6214 => x"01da61b9",
			6215 => x"0d060f0c",
			6216 => x"0c04cd04",
			6217 => x"fc3061b9",
			6218 => x"040cc604",
			6219 => x"feef61b9",
			6220 => x"008761b9",
			6221 => x"0b054508",
			6222 => x"06016c04",
			6223 => x"000061b9",
			6224 => x"019261b9",
			6225 => x"040b3604",
			6226 => x"fff561b9",
			6227 => x"ff0e61b9",
			6228 => x"0d086514",
			6229 => x"08034c04",
			6230 => x"01a461b9",
			6231 => x"0c054508",
			6232 => x"08035604",
			6233 => x"ff3661b9",
			6234 => x"019061b9",
			6235 => x"0100fc04",
			6236 => x"fdbe61b9",
			6237 => x"00b961b9",
			6238 => x"0f0adf0c",
			6239 => x"0b06ff04",
			6240 => x"008461b9",
			6241 => x"0e0a1b04",
			6242 => x"000061b9",
			6243 => x"fe5c61b9",
			6244 => x"00039d08",
			6245 => x"0f0aed04",
			6246 => x"ffc461b9",
			6247 => x"01eb61b9",
			6248 => x"0a027404",
			6249 => x"fec061b9",
			6250 => x"006261b9",
			6251 => x"0505f904",
			6252 => x"000061b9",
			6253 => x"fe5761b9",
			6254 => x"040ae248",
			6255 => x"0409db18",
			6256 => x"03097814",
			6257 => x"0a021d10",
			6258 => x"0b06cd0c",
			6259 => x"01010f04",
			6260 => x"0000630d",
			6261 => x"0b06bc04",
			6262 => x"0000630d",
			6263 => x"00d9630d",
			6264 => x"0000630d",
			6265 => x"0000630d",
			6266 => x"ffa0630d",
			6267 => x"030a1220",
			6268 => x"07059110",
			6269 => x"0c05050c",
			6270 => x"0306e204",
			6271 => x"0000630d",
			6272 => x"07052f04",
			6273 => x"00d0630d",
			6274 => x"0000630d",
			6275 => x"ff81630d",
			6276 => x"0c06140c",
			6277 => x"09021208",
			6278 => x"0901d904",
			6279 => x"0122630d",
			6280 => x"005e630d",
			6281 => x"0000630d",
			6282 => x"0000630d",
			6283 => x"0c062e08",
			6284 => x"020a5b04",
			6285 => x"ff43630d",
			6286 => x"0000630d",
			6287 => x"0c065004",
			6288 => x"0098630d",
			6289 => x"0000630d",
			6290 => x"040aef0c",
			6291 => x"01013208",
			6292 => x"0003f704",
			6293 => x"fecf630d",
			6294 => x"0000630d",
			6295 => x"0000630d",
			6296 => x"0f0ad13c",
			6297 => x"07052f1c",
			6298 => x"0306b910",
			6299 => x"0b053508",
			6300 => x"040c0404",
			6301 => x"ff5f630d",
			6302 => x"007f630d",
			6303 => x"0208c704",
			6304 => x"0000630d",
			6305 => x"ff15630d",
			6306 => x"0a029204",
			6307 => x"ff7f630d",
			6308 => x"02093504",
			6309 => x"0110630d",
			6310 => x"0000630d",
			6311 => x"0a02db10",
			6312 => x"0901db08",
			6313 => x"0a025f04",
			6314 => x"0000630d",
			6315 => x"fee6630d",
			6316 => x"0b071e04",
			6317 => x"0022630d",
			6318 => x"0000630d",
			6319 => x"0a02fd08",
			6320 => x"0e06e204",
			6321 => x"0000630d",
			6322 => x"009b630d",
			6323 => x"07053104",
			6324 => x"0000630d",
			6325 => x"ffc6630d",
			6326 => x"0a02d110",
			6327 => x"00039204",
			6328 => x"0000630d",
			6329 => x"07069b04",
			6330 => x"00f0630d",
			6331 => x"0706b704",
			6332 => x"0000630d",
			6333 => x"0051630d",
			6334 => x"0e0cbb08",
			6335 => x"020bbc04",
			6336 => x"0000630d",
			6337 => x"fee4630d",
			6338 => x"0000630d",
			6339 => x"06017448",
			6340 => x"0505cc04",
			6341 => x"fe9f6439",
			6342 => x"0f080e1c",
			6343 => x"0601640c",
			6344 => x"0207b508",
			6345 => x"00028d04",
			6346 => x"00006439",
			6347 => x"00836439",
			6348 => x"fee26439",
			6349 => x"040bb704",
			6350 => x"00006439",
			6351 => x"03063204",
			6352 => x"00006439",
			6353 => x"0c050704",
			6354 => x"01586439",
			6355 => x"00006439",
			6356 => x"040adc14",
			6357 => x"09011b08",
			6358 => x"040aa904",
			6359 => x"00006439",
			6360 => x"010b6439",
			6361 => x"09019604",
			6362 => x"fec96439",
			6363 => x"0c061304",
			6364 => x"00036439",
			6365 => x"ff046439",
			6366 => x"0209190c",
			6367 => x"0208e404",
			6368 => x"ff7c6439",
			6369 => x"0c04ec04",
			6370 => x"002d6439",
			6371 => x"00006439",
			6372 => x"0c05d504",
			6373 => x"fe6c6439",
			6374 => x"00006439",
			6375 => x"0705181c",
			6376 => x"0b055218",
			6377 => x"0f088514",
			6378 => x"0c04ea10",
			6379 => x"0d05e908",
			6380 => x"02091104",
			6381 => x"ffd56439",
			6382 => x"00206439",
			6383 => x"0900cd04",
			6384 => x"00006439",
			6385 => x"017d6439",
			6386 => x"ffa36439",
			6387 => x"ff256439",
			6388 => x"01846439",
			6389 => x"0c04cd08",
			6390 => x"08033104",
			6391 => x"00006439",
			6392 => x"fe6a6439",
			6393 => x"00047d1c",
			6394 => x"0a02bf10",
			6395 => x"08036308",
			6396 => x"08034104",
			6397 => x"ffed6439",
			6398 => x"00c36439",
			6399 => x"0f08dd04",
			6400 => x"00006439",
			6401 => x"fdae6439",
			6402 => x"0c061504",
			6403 => x"01866439",
			6404 => x"0f0c3904",
			6405 => x"feaa6439",
			6406 => x"00cc6439",
			6407 => x"07051f04",
			6408 => x"001b6439",
			6409 => x"030d4e04",
			6410 => x"fe956439",
			6411 => x"0a038804",
			6412 => x"002b6439",
			6413 => x"00006439",
			6414 => x"03061114",
			6415 => x"06017404",
			6416 => x"fe67657d",
			6417 => x"0b051104",
			6418 => x"ff74657d",
			6419 => x"02093a04",
			6420 => x"01c3657d",
			6421 => x"0a035404",
			6422 => x"ff9f657d",
			6423 => x"0000657d",
			6424 => x"06018a44",
			6425 => x"0b06ee30",
			6426 => x"06014a10",
			6427 => x"0900fb0c",
			6428 => x"01009704",
			6429 => x"fedc657d",
			6430 => x"0001fa04",
			6431 => x"0000657d",
			6432 => x"0125657d",
			6433 => x"fe89657d",
			6434 => x"040a5b10",
			6435 => x"0901df08",
			6436 => x"09010f04",
			6437 => x"feb3657d",
			6438 => x"013b657d",
			6439 => x"0a024c04",
			6440 => x"fef3657d",
			6441 => x"01e8657d",
			6442 => x"0f082b08",
			6443 => x"040c9304",
			6444 => x"0039657d",
			6445 => x"01ce657d",
			6446 => x"0d061d04",
			6447 => x"fe0b657d",
			6448 => x"000a657d",
			6449 => x"0101190c",
			6450 => x"0f0a0304",
			6451 => x"fe9b657d",
			6452 => x"0100fa04",
			6453 => x"0000657d",
			6454 => x"01ad657d",
			6455 => x"0802ed04",
			6456 => x"fe65657d",
			6457 => x"fc3c657d",
			6458 => x"0508041c",
			6459 => x"040d2e10",
			6460 => x"0e089608",
			6461 => x"0b05a704",
			6462 => x"01ab657d",
			6463 => x"ff3b657d",
			6464 => x"0802eb04",
			6465 => x"003f657d",
			6466 => x"01a7657d",
			6467 => x"09010204",
			6468 => x"01ae657d",
			6469 => x"0601a604",
			6470 => x"fe3d657d",
			6471 => x"002b657d",
			6472 => x"0f0ad914",
			6473 => x"0902280c",
			6474 => x"0d086604",
			6475 => x"0000657d",
			6476 => x"0f0acb04",
			6477 => x"fe2f657d",
			6478 => x"ffec657d",
			6479 => x"0f0a9204",
			6480 => x"0219657d",
			6481 => x"fee3657d",
			6482 => x"040c4410",
			6483 => x"01016008",
			6484 => x"0f0aed04",
			6485 => x"ff98657d",
			6486 => x"01da657d",
			6487 => x"0d090104",
			6488 => x"004f657d",
			6489 => x"fe8d657d",
			6490 => x"0004a008",
			6491 => x"040cd804",
			6492 => x"ff18657d",
			6493 => x"00ad657d",
			6494 => x"fe6b657d",
			6495 => x"0b051408",
			6496 => x"02093d04",
			6497 => x"febe6671",
			6498 => x"00006671",
			6499 => x"0c04b914",
			6500 => x"040b7008",
			6501 => x"03071b04",
			6502 => x"fec46671",
			6503 => x"008c6671",
			6504 => x"0505b104",
			6505 => x"00006671",
			6506 => x"06016704",
			6507 => x"00006671",
			6508 => x"01756671",
			6509 => x"040ae224",
			6510 => x"05061508",
			6511 => x"06016804",
			6512 => x"00006671",
			6513 => x"01646671",
			6514 => x"03076c0c",
			6515 => x"0f07a308",
			6516 => x"0c054c04",
			6517 => x"00006671",
			6518 => x"00356671",
			6519 => x"fe886671",
			6520 => x"00037008",
			6521 => x"0209e804",
			6522 => x"00196671",
			6523 => x"fefe6671",
			6524 => x"0507ea04",
			6525 => x"00f76671",
			6526 => x"00006671",
			6527 => x"0601851c",
			6528 => x"0b05430c",
			6529 => x"0d05ed04",
			6530 => x"ff3c6671",
			6531 => x"02094304",
			6532 => x"01056671",
			6533 => x"ffbb6671",
			6534 => x"040b4a08",
			6535 => x"00040204",
			6536 => x"fe3f6671",
			6537 => x"ffec6671",
			6538 => x"03075404",
			6539 => x"ff226671",
			6540 => x"00f86671",
			6541 => x"0c054310",
			6542 => x"00042e08",
			6543 => x"05065e04",
			6544 => x"007e6671",
			6545 => x"ffb16671",
			6546 => x"0b054304",
			6547 => x"00006671",
			6548 => x"01516671",
			6549 => x"0e09fd08",
			6550 => x"040b8304",
			6551 => x"007b6671",
			6552 => x"fe5e6671",
			6553 => x"0d087f04",
			6554 => x"00f96671",
			6555 => x"ffd56671",
			6556 => x"0507f688",
			6557 => x"0705e64c",
			6558 => x"08034218",
			6559 => x"0c04d008",
			6560 => x"06017004",
			6561 => x"0000681d",
			6562 => x"000f681d",
			6563 => x"0f082b04",
			6564 => x"0000681d",
			6565 => x"0208b904",
			6566 => x"0000681d",
			6567 => x"06019604",
			6568 => x"fef1681d",
			6569 => x"0000681d",
			6570 => x"0306e21c",
			6571 => x"0f082210",
			6572 => x"03063a08",
			6573 => x"0f07b904",
			6574 => x"0000681d",
			6575 => x"ff40681d",
			6576 => x"01008a04",
			6577 => x"00af681d",
			6578 => x"fff6681d",
			6579 => x"0704f104",
			6580 => x"0000681d",
			6581 => x"06018004",
			6582 => x"fec7681d",
			6583 => x"0000681d",
			6584 => x"02094d08",
			6585 => x"00043604",
			6586 => x"0110681d",
			6587 => x"0000681d",
			6588 => x"0a02bf08",
			6589 => x"0c04ea04",
			6590 => x"0000681d",
			6591 => x"ff53681d",
			6592 => x"0803dc04",
			6593 => x"00b2681d",
			6594 => x"ffaf681d",
			6595 => x"0f096018",
			6596 => x"0c05d710",
			6597 => x"0a02330c",
			6598 => x"07062c08",
			6599 => x"01012404",
			6600 => x"0070681d",
			6601 => x"0000681d",
			6602 => x"0000681d",
			6603 => x"0000681d",
			6604 => x"07066d04",
			6605 => x"ff46681d",
			6606 => x"0000681d",
			6607 => x"07065518",
			6608 => x"07062e0c",
			6609 => x"0c05f608",
			6610 => x"0c059f04",
			6611 => x"0000681d",
			6612 => x"00bd681d",
			6613 => x"0000681d",
			6614 => x"0f097104",
			6615 => x"0000681d",
			6616 => x"07064104",
			6617 => x"ff6a681d",
			6618 => x"0000681d",
			6619 => x"0c05d504",
			6620 => x"0000681d",
			6621 => x"0d080a04",
			6622 => x"0000681d",
			6623 => x"00ea681d",
			6624 => x"030a9918",
			6625 => x"0101450c",
			6626 => x"0706ca08",
			6627 => x"09020804",
			6628 => x"fec2681d",
			6629 => x"0000681d",
			6630 => x"0000681d",
			6631 => x"07066d04",
			6632 => x"004e681d",
			6633 => x"07068804",
			6634 => x"ffb6681d",
			6635 => x"0000681d",
			6636 => x"0d08b30c",
			6637 => x"0c05f504",
			6638 => x"0000681d",
			6639 => x"0f0b0904",
			6640 => x"0000681d",
			6641 => x"00b8681d",
			6642 => x"0e0b7718",
			6643 => x"0601900c",
			6644 => x"0c068404",
			6645 => x"0000681d",
			6646 => x"0706de04",
			6647 => x"0000681d",
			6648 => x"006c681d",
			6649 => x"0a026404",
			6650 => x"0000681d",
			6651 => x"05091b04",
			6652 => x"feec681d",
			6653 => x"0000681d",
			6654 => x"0d0a2b0c",
			6655 => x"01013b04",
			6656 => x"0000681d",
			6657 => x"020bbc04",
			6658 => x"0000681d",
			6659 => x"00bb681d",
			6660 => x"0c071e04",
			6661 => x"ffa5681d",
			6662 => x"0000681d",
			6663 => x"0505b114",
			6664 => x"02093504",
			6665 => x"fe786909",
			6666 => x"040df504",
			6667 => x"ff3a6909",
			6668 => x"0209b108",
			6669 => x"0004d204",
			6670 => x"00006909",
			6671 => x"00bf6909",
			6672 => x"ff836909",
			6673 => x"0d0a2b60",
			6674 => x"040b9d3c",
			6675 => x"0100f81c",
			6676 => x"02093510",
			6677 => x"0003f208",
			6678 => x"0100a804",
			6679 => x"fe836909",
			6680 => x"003a6909",
			6681 => x"0c050704",
			6682 => x"00b96909",
			6683 => x"fdf16909",
			6684 => x"08036808",
			6685 => x"0a02a804",
			6686 => x"fe926909",
			6687 => x"00836909",
			6688 => x"fd726909",
			6689 => x"0507f510",
			6690 => x"0c05f808",
			6691 => x"0209b704",
			6692 => x"ffff6909",
			6693 => x"00f46909",
			6694 => x"0b06dd04",
			6695 => x"01776909",
			6696 => x"000f6909",
			6697 => x"01014508",
			6698 => x"0100ff04",
			6699 => x"01296909",
			6700 => x"ff116909",
			6701 => x"0706f504",
			6702 => x"00cf6909",
			6703 => x"ff926909",
			6704 => x"0c04b208",
			6705 => x"06016704",
			6706 => x"00006909",
			6707 => x"01cb6909",
			6708 => x"0e06000c",
			6709 => x"07051808",
			6710 => x"040cc604",
			6711 => x"ff046909",
			6712 => x"011f6909",
			6713 => x"fe356909",
			6714 => x"0c052a08",
			6715 => x"0505db04",
			6716 => x"ff586909",
			6717 => x"011d6909",
			6718 => x"020ad604",
			6719 => x"fecc6909",
			6720 => x"00736909",
			6721 => x"fe546909",
			6722 => x"09010f50",
			6723 => x"0704f120",
			6724 => x"06016404",
			6725 => x"fec46a7d",
			6726 => x"03063a10",
			6727 => x"0704eb0c",
			6728 => x"0b04e304",
			6729 => x"00006a7d",
			6730 => x"06017404",
			6731 => x"00006a7d",
			6732 => x"01016a7d",
			6733 => x"ff5c6a7d",
			6734 => x"02095d08",
			6735 => x"0704ea04",
			6736 => x"00006a7d",
			6737 => x"017c6a7d",
			6738 => x"00006a7d",
			6739 => x"040e6320",
			6740 => x"0f08cd18",
			6741 => x"06018510",
			6742 => x"02092e08",
			6743 => x"0c050704",
			6744 => x"00026a7d",
			6745 => x"fe856a7d",
			6746 => x"0d062b04",
			6747 => x"fe8d6a7d",
			6748 => x"ffd56a7d",
			6749 => x"06018a04",
			6750 => x"01296a7d",
			6751 => x"00006a7d",
			6752 => x"06019404",
			6753 => x"fe096a7d",
			6754 => x"00006a7d",
			6755 => x"0c050d0c",
			6756 => x"06017804",
			6757 => x"00006a7d",
			6758 => x"04118b04",
			6759 => x"01236a7d",
			6760 => x"00006a7d",
			6761 => x"00006a7d",
			6762 => x"0f09e130",
			6763 => x"0b06e02c",
			6764 => x"0b06bc18",
			6765 => x"0802d70c",
			6766 => x"03071b04",
			6767 => x"00006a7d",
			6768 => x"0f09b104",
			6769 => x"feb26a7d",
			6770 => x"00006a7d",
			6771 => x"0f09b108",
			6772 => x"05065104",
			6773 => x"00e26a7d",
			6774 => x"ffd06a7d",
			6775 => x"017b6a7d",
			6776 => x"07062b04",
			6777 => x"ffde6a7d",
			6778 => x"07063d08",
			6779 => x"0209a404",
			6780 => x"02396a7d",
			6781 => x"00006a7d",
			6782 => x"07064304",
			6783 => x"00006a7d",
			6784 => x"00e36a7d",
			6785 => x"ff2c6a7d",
			6786 => x"0901870c",
			6787 => x"07058d04",
			6788 => x"00006a7d",
			6789 => x"00040704",
			6790 => x"00006a7d",
			6791 => x"fe646a7d",
			6792 => x"0507d810",
			6793 => x"00037804",
			6794 => x"00006a7d",
			6795 => x"0f0ad108",
			6796 => x"0901fe04",
			6797 => x"01636a7d",
			6798 => x"00006a7d",
			6799 => x"00006a7d",
			6800 => x"05083e10",
			6801 => x"030a9908",
			6802 => x"040bc404",
			6803 => x"ff8d6a7d",
			6804 => x"fe2c6a7d",
			6805 => x"0f0b9804",
			6806 => x"01056a7d",
			6807 => x"00006a7d",
			6808 => x"0b073308",
			6809 => x"0b071e04",
			6810 => x"00006a7d",
			6811 => x"01586a7d",
			6812 => x"0c063304",
			6813 => x"fee66a7d",
			6814 => x"003c6a7d",
			6815 => x"06016c58",
			6816 => x"0100fa30",
			6817 => x"0601671c",
			6818 => x"0600e808",
			6819 => x"0c052e04",
			6820 => x"fe7a6c19",
			6821 => x"044e6c19",
			6822 => x"03069604",
			6823 => x"fe5c6c19",
			6824 => x"0e064308",
			6825 => x"06015f04",
			6826 => x"fef06c19",
			6827 => x"04346c19",
			6828 => x"0d070804",
			6829 => x"ff416c19",
			6830 => x"fe5e6c19",
			6831 => x"02090c10",
			6832 => x"0e05e004",
			6833 => x"fe736c19",
			6834 => x"0a02ac08",
			6835 => x"0003fb04",
			6836 => x"00c66c19",
			6837 => x"fe766c19",
			6838 => x"03596c19",
			6839 => x"fe676c19",
			6840 => x"03092e08",
			6841 => x"0100ff04",
			6842 => x"00ee6c19",
			6843 => x"fe666c19",
			6844 => x"00032410",
			6845 => x"07063f04",
			6846 => x"02c96c19",
			6847 => x"01011d08",
			6848 => x"0b06cd04",
			6849 => x"00c16c19",
			6850 => x"fe706c19",
			6851 => x"01ab6c19",
			6852 => x"0a02390c",
			6853 => x"01011304",
			6854 => x"08316c19",
			6855 => x"0d083104",
			6856 => x"03f56c19",
			6857 => x"ffef6c19",
			6858 => x"fe456c19",
			6859 => x"0b07634c",
			6860 => x"0802e824",
			6861 => x"040adc1c",
			6862 => x"00038110",
			6863 => x"0507ca08",
			6864 => x"0e096204",
			6865 => x"00376c19",
			6866 => x"04c06c19",
			6867 => x"020a4604",
			6868 => x"fee36c19",
			6869 => x"01186c19",
			6870 => x"00038c08",
			6871 => x"0e098704",
			6872 => x"001a6c19",
			6873 => x"046d6c19",
			6874 => x"01506c19",
			6875 => x"05086a04",
			6876 => x"fe3d6c19",
			6877 => x"00696c19",
			6878 => x"040c6010",
			6879 => x"0d05ed04",
			6880 => x"fe216c19",
			6881 => x"0706ca08",
			6882 => x"00039604",
			6883 => x"00496c19",
			6884 => x"02416c19",
			6885 => x"078c6c19",
			6886 => x"0c04f10c",
			6887 => x"0505a004",
			6888 => x"fe766c19",
			6889 => x"0411a304",
			6890 => x"028a6c19",
			6891 => x"ff506c19",
			6892 => x"06018104",
			6893 => x"fe616c19",
			6894 => x"07058d04",
			6895 => x"01b66c19",
			6896 => x"fef96c19",
			6897 => x"01017f24",
			6898 => x"0706ca0c",
			6899 => x"020ba008",
			6900 => x"0b077104",
			6901 => x"01c46c19",
			6902 => x"fe666c19",
			6903 => x"02db6c19",
			6904 => x"0101300c",
			6905 => x"0a02ab08",
			6906 => x"0d098504",
			6907 => x"01716c19",
			6908 => x"10056c19",
			6909 => x"fe5f6c19",
			6910 => x"0d097504",
			6911 => x"fe5d6c19",
			6912 => x"0508fd04",
			6913 => x"07a66c19",
			6914 => x"fe726c19",
			6915 => x"020cab04",
			6916 => x"fe716c19",
			6917 => x"02b36c19",
			6918 => x"0e078e6c",
			6919 => x"0b056348",
			6920 => x"0d062a30",
			6921 => x"040b9d14",
			6922 => x"0208b408",
			6923 => x"0306a504",
			6924 => x"ffb46ddd",
			6925 => x"00756ddd",
			6926 => x"08032604",
			6927 => x"00006ddd",
			6928 => x"00042804",
			6929 => x"fe8b6ddd",
			6930 => x"00006ddd",
			6931 => x"03063a0c",
			6932 => x"0a02ed04",
			6933 => x"fee86ddd",
			6934 => x"0b050404",
			6935 => x"00006ddd",
			6936 => x"009c6ddd",
			6937 => x"0c04d408",
			6938 => x"0d05ed04",
			6939 => x"00006ddd",
			6940 => x"00f96ddd",
			6941 => x"08039904",
			6942 => x"ff426ddd",
			6943 => x"000f6ddd",
			6944 => x"00043208",
			6945 => x"06016804",
			6946 => x"00006ddd",
			6947 => x"01686ddd",
			6948 => x"0e06ac08",
			6949 => x"0306a504",
			6950 => x"00006ddd",
			6951 => x"01256ddd",
			6952 => x"06018904",
			6953 => x"fefc6ddd",
			6954 => x"00466ddd",
			6955 => x"00042810",
			6956 => x"0c04ce04",
			6957 => x"00006ddd",
			6958 => x"03076c08",
			6959 => x"040a4904",
			6960 => x"00006ddd",
			6961 => x"fdf46ddd",
			6962 => x"00006ddd",
			6963 => x"0d065208",
			6964 => x"0306ff04",
			6965 => x"00006ddd",
			6966 => x"01186ddd",
			6967 => x"0a02c704",
			6968 => x"fedd6ddd",
			6969 => x"03079c04",
			6970 => x"00006ddd",
			6971 => x"ffc76ddd",
			6972 => x"040b8540",
			6973 => x"06018a20",
			6974 => x"0c058308",
			6975 => x"05065104",
			6976 => x"00006ddd",
			6977 => x"fec36ddd",
			6978 => x"09020a0c",
			6979 => x"0802dd08",
			6980 => x"0901a904",
			6981 => x"00966ddd",
			6982 => x"00036ddd",
			6983 => x"01366ddd",
			6984 => x"040a9504",
			6985 => x"00006ddd",
			6986 => x"09020e04",
			6987 => x"00006ddd",
			6988 => x"ff366ddd",
			6989 => x"0d086504",
			6990 => x"016e6ddd",
			6991 => x"0f0aed0c",
			6992 => x"020a5b04",
			6993 => x"004c6ddd",
			6994 => x"0b070e04",
			6995 => x"00006ddd",
			6996 => x"ff156ddd",
			6997 => x"0b079308",
			6998 => x"09022b04",
			6999 => x"01326ddd",
			7000 => x"00006ddd",
			7001 => x"09022e04",
			7002 => x"ffdb6ddd",
			7003 => x"004c6ddd",
			7004 => x"0803341c",
			7005 => x"030a8a0c",
			7006 => x"06018804",
			7007 => x"00006ddd",
			7008 => x"0e0aa404",
			7009 => x"fe456ddd",
			7010 => x"00006ddd",
			7011 => x"05088608",
			7012 => x"0003d804",
			7013 => x"00006ddd",
			7014 => x"00d36ddd",
			7015 => x"0901c304",
			7016 => x"00006ddd",
			7017 => x"ffdc6ddd",
			7018 => x"0c050a04",
			7019 => x"ff426ddd",
			7020 => x"0c058508",
			7021 => x"040baa04",
			7022 => x"00006ddd",
			7023 => x"01386ddd",
			7024 => x"0e0c7e08",
			7025 => x"08035504",
			7026 => x"00836ddd",
			7027 => x"ff516ddd",
			7028 => x"0004bc04",
			7029 => x"01086ddd",
			7030 => x"00006ddd",
			7031 => x"0b051114",
			7032 => x"02093d04",
			7033 => x"fe846f11",
			7034 => x"0209b10c",
			7035 => x"0900ac08",
			7036 => x"09005d04",
			7037 => x"00006f11",
			7038 => x"00446f11",
			7039 => x"00006f11",
			7040 => x"ff9d6f11",
			7041 => x"0704f124",
			7042 => x"0f081614",
			7043 => x"0208ab04",
			7044 => x"ff246f11",
			7045 => x"0c04ec0c",
			7046 => x"0b051204",
			7047 => x"00006f11",
			7048 => x"0a029504",
			7049 => x"00006f11",
			7050 => x"01886f11",
			7051 => x"00006f11",
			7052 => x"02095d0c",
			7053 => x"0306b904",
			7054 => x"ff586f11",
			7055 => x"0003fb04",
			7056 => x"fffa6f11",
			7057 => x"01566f11",
			7058 => x"febb6f11",
			7059 => x"09012040",
			7060 => x"0208c720",
			7061 => x"0208a410",
			7062 => x"09010f08",
			7063 => x"0a01fa04",
			7064 => x"00006f11",
			7065 => x"ff236f11",
			7066 => x"05066c04",
			7067 => x"000f6f11",
			7068 => x"00006f11",
			7069 => x"07050808",
			7070 => x"03063204",
			7071 => x"00006f11",
			7072 => x"01696f11",
			7073 => x"05069904",
			7074 => x"ff326f11",
			7075 => x"00ff6f11",
			7076 => x"05062610",
			7077 => x"0d062b08",
			7078 => x"040c1e04",
			7079 => x"feab6f11",
			7080 => x"ffe26f11",
			7081 => x"00040204",
			7082 => x"fed56f11",
			7083 => x"00b26f11",
			7084 => x"02097b08",
			7085 => x"0d064504",
			7086 => x"00006f11",
			7087 => x"fdf46f11",
			7088 => x"0c050504",
			7089 => x"00b96f11",
			7090 => x"ff2a6f11",
			7091 => x"05067908",
			7092 => x"0e083c04",
			7093 => x"01b76f11",
			7094 => x"ff736f11",
			7095 => x"0308750c",
			7096 => x"0207cf08",
			7097 => x"0f071f04",
			7098 => x"00006f11",
			7099 => x"00ad6f11",
			7100 => x"fe656f11",
			7101 => x"07058d08",
			7102 => x"00041404",
			7103 => x"00006f11",
			7104 => x"01bb6f11",
			7105 => x"0705d104",
			7106 => x"fe4d6f11",
			7107 => x"00046f11",
			7108 => x"06017450",
			7109 => x"0505cc04",
			7110 => x"fe95706d",
			7111 => x"01007d10",
			7112 => x"0f08050c",
			7113 => x"08036e04",
			7114 => x"0000706d",
			7115 => x"03063204",
			7116 => x"0000706d",
			7117 => x"018e706d",
			7118 => x"ffa0706d",
			7119 => x"0802aa1c",
			7120 => x"040a0110",
			7121 => x"0d082208",
			7122 => x"00033504",
			7123 => x"008b706d",
			7124 => x"ff17706d",
			7125 => x"0d085904",
			7126 => x"fea2706d",
			7127 => x"0000706d",
			7128 => x"06016004",
			7129 => x"0000706d",
			7130 => x"03096804",
			7131 => x"0000706d",
			7132 => x"0192706d",
			7133 => x"0f084610",
			7134 => x"0e068d08",
			7135 => x"0900d904",
			7136 => x"0000706d",
			7137 => x"ff25706d",
			7138 => x"040aa104",
			7139 => x"0000706d",
			7140 => x"00d2706d",
			7141 => x"0c05da08",
			7142 => x"0c04ce04",
			7143 => x"fff7706d",
			7144 => x"fe7b706d",
			7145 => x"0d083f04",
			7146 => x"ff28706d",
			7147 => x"0076706d",
			7148 => x"0d064730",
			7149 => x"0b055224",
			7150 => x"0d062a1c",
			7151 => x"0b053510",
			7152 => x"0900d308",
			7153 => x"0b04f304",
			7154 => x"0000706d",
			7155 => x"0153706d",
			7156 => x"00045304",
			7157 => x"003a706d",
			7158 => x"fed9706d",
			7159 => x"0d061d08",
			7160 => x"0505f604",
			7161 => x"ff98706d",
			7162 => x"fe54706d",
			7163 => x"0000706d",
			7164 => x"00040b04",
			7165 => x"0000706d",
			7166 => x"0171706d",
			7167 => x"0003f104",
			7168 => x"0000706d",
			7169 => x"0f080e04",
			7170 => x"0000706d",
			7171 => x"01cf706d",
			7172 => x"09010f10",
			7173 => x"0a02bf04",
			7174 => x"fe03706d",
			7175 => x"0d066d08",
			7176 => x"03071b04",
			7177 => x"0000706d",
			7178 => x"00c5706d",
			7179 => x"0000706d",
			7180 => x"05065108",
			7181 => x"06018104",
			7182 => x"0051706d",
			7183 => x"0190706d",
			7184 => x"0e07dc08",
			7185 => x"06017704",
			7186 => x"0000706d",
			7187 => x"fe65706d",
			7188 => x"0c054608",
			7189 => x"08035304",
			7190 => x"ffb1706d",
			7191 => x"0178706d",
			7192 => x"040b8304",
			7193 => x"0050706d",
			7194 => x"ff7c706d",
			7195 => x"0b051110",
			7196 => x"02093d04",
			7197 => x"fe6b71b1",
			7198 => x"0d05a804",
			7199 => x"fec571b1",
			7200 => x"0d05c204",
			7201 => x"00ce71b1",
			7202 => x"000071b1",
			7203 => x"040a5b40",
			7204 => x"02098e20",
			7205 => x"0f097d1c",
			7206 => x"0f09600c",
			7207 => x"0a027808",
			7208 => x"0d082204",
			7209 => x"002771b1",
			7210 => x"fea071b1",
			7211 => x"017271b1",
			7212 => x"02096008",
			7213 => x"03097804",
			7214 => x"022871b1",
			7215 => x"000071b1",
			7216 => x"0c061304",
			7217 => x"ff4371b1",
			7218 => x"006e71b1",
			7219 => x"fe7671b1",
			7220 => x"0e09870c",
			7221 => x"0f09a304",
			7222 => x"ff3b71b1",
			7223 => x"07065a04",
			7224 => x"019671b1",
			7225 => x"03f371b1",
			7226 => x"0209ce0c",
			7227 => x"07065c04",
			7228 => x"fe8571b1",
			7229 => x"01012a04",
			7230 => x"ff9271b1",
			7231 => x"004771b1",
			7232 => x"0a023904",
			7233 => x"021071b1",
			7234 => x"ff4c71b1",
			7235 => x"0c04e924",
			7236 => x"0003ea0c",
			7237 => x"0003e508",
			7238 => x"08031804",
			7239 => x"ff5f71b1",
			7240 => x"00da71b1",
			7241 => x"fb6d71b1",
			7242 => x"040d0010",
			7243 => x"03065908",
			7244 => x"0c04b204",
			7245 => x"003071b1",
			7246 => x"fe3d71b1",
			7247 => x"02091104",
			7248 => x"017371b1",
			7249 => x"000c71b1",
			7250 => x"07051804",
			7251 => x"01b771b1",
			7252 => x"000071b1",
			7253 => x"0308c71c",
			7254 => x"08034410",
			7255 => x"0003b808",
			7256 => x"0a025c04",
			7257 => x"ff3871b1",
			7258 => x"014b71b1",
			7259 => x"00040304",
			7260 => x"fe3271b1",
			7261 => x"ffa971b1",
			7262 => x"040b3604",
			7263 => x"01ce71b1",
			7264 => x"0c052a04",
			7265 => x"ffd571b1",
			7266 => x"fe2871b1",
			7267 => x"0705a304",
			7268 => x"020a71b1",
			7269 => x"0003ee08",
			7270 => x"00037004",
			7271 => x"ff1c71b1",
			7272 => x"009071b1",
			7273 => x"08032b04",
			7274 => x"fccd71b1",
			7275 => x"ffba71b1",
			7276 => x"0507f688",
			7277 => x"0705e64c",
			7278 => x"08034218",
			7279 => x"0c04d008",
			7280 => x"06017004",
			7281 => x"0000735d",
			7282 => x"0011735d",
			7283 => x"0d061d04",
			7284 => x"0000735d",
			7285 => x"08027904",
			7286 => x"0000735d",
			7287 => x"06019604",
			7288 => x"ff0d735d",
			7289 => x"0000735d",
			7290 => x"0306e21c",
			7291 => x"0f082210",
			7292 => x"03063a08",
			7293 => x"0f07b904",
			7294 => x"0000735d",
			7295 => x"ff55735d",
			7296 => x"01008a04",
			7297 => x"00a1735d",
			7298 => x"fffe735d",
			7299 => x"0704f104",
			7300 => x"0000735d",
			7301 => x"06018004",
			7302 => x"fed8735d",
			7303 => x"0000735d",
			7304 => x"0f087208",
			7305 => x"05064204",
			7306 => x"0126735d",
			7307 => x"0000735d",
			7308 => x"06018c08",
			7309 => x"02093504",
			7310 => x"0000735d",
			7311 => x"ff75735d",
			7312 => x"020b2404",
			7313 => x"009b735d",
			7314 => x"0000735d",
			7315 => x"0f095614",
			7316 => x"0c05d710",
			7317 => x"0209000c",
			7318 => x"0d07f108",
			7319 => x"0f07dc04",
			7320 => x"0000735d",
			7321 => x"0039735d",
			7322 => x"0000735d",
			7323 => x"0000735d",
			7324 => x"ff57735d",
			7325 => x"07065518",
			7326 => x"07062e0c",
			7327 => x"0c05f608",
			7328 => x"0c059f04",
			7329 => x"0000735d",
			7330 => x"00a9735d",
			7331 => x"0000735d",
			7332 => x"0f097104",
			7333 => x"0000735d",
			7334 => x"07064104",
			7335 => x"ff79735d",
			7336 => x"0000735d",
			7337 => x"0f097104",
			7338 => x"0000735d",
			7339 => x"0b06cb04",
			7340 => x"0000735d",
			7341 => x"0b06fc04",
			7342 => x"00dc735d",
			7343 => x"0000735d",
			7344 => x"030a9918",
			7345 => x"0101450c",
			7346 => x"0706ca08",
			7347 => x"09020804",
			7348 => x"fed4735d",
			7349 => x"0000735d",
			7350 => x"0000735d",
			7351 => x"07066d04",
			7352 => x"003a735d",
			7353 => x"07068804",
			7354 => x"ffd0735d",
			7355 => x"0000735d",
			7356 => x"05086a08",
			7357 => x"01013f04",
			7358 => x"0000735d",
			7359 => x"00bc735d",
			7360 => x"030ba618",
			7361 => x"0601900c",
			7362 => x"0c068404",
			7363 => x"0000735d",
			7364 => x"0706de04",
			7365 => x"0000735d",
			7366 => x"005f735d",
			7367 => x"0a026404",
			7368 => x"0000735d",
			7369 => x"05091b04",
			7370 => x"fed0735d",
			7371 => x"0000735d",
			7372 => x"0c06a40c",
			7373 => x"01015404",
			7374 => x"0000735d",
			7375 => x"08032604",
			7376 => x"0000735d",
			7377 => x"00b8735d",
			7378 => x"07077d04",
			7379 => x"ff4a735d",
			7380 => x"0601d004",
			7381 => x"0085735d",
			7382 => x"0000735d",
			7383 => x"0e078e6c",
			7384 => x"0f082b34",
			7385 => x"03069624",
			7386 => x"0208f70c",
			7387 => x"040c2c08",
			7388 => x"0d069f04",
			7389 => x"fed37531",
			7390 => x"00007531",
			7391 => x"00007531",
			7392 => x"0601700c",
			7393 => x"01007508",
			7394 => x"0505df04",
			7395 => x"00007531",
			7396 => x"000f7531",
			7397 => x"ff047531",
			7398 => x"03063a08",
			7399 => x"0505ea04",
			7400 => x"000b7531",
			7401 => x"ffc57531",
			7402 => x"01347531",
			7403 => x"0208ad04",
			7404 => x"00007531",
			7405 => x"0c04cd04",
			7406 => x"00007531",
			7407 => x"0004bc04",
			7408 => x"01407531",
			7409 => x"00007531",
			7410 => x"040bb218",
			7411 => x"0c04cc08",
			7412 => x"06017404",
			7413 => x"00007531",
			7414 => x"009b7531",
			7415 => x"0100a608",
			7416 => x"06016b04",
			7417 => x"00007531",
			7418 => x"fec07531",
			7419 => x"06017404",
			7420 => x"fff97531",
			7421 => x"00387531",
			7422 => x"0004580c",
			7423 => x"06017404",
			7424 => x"00007531",
			7425 => x"05064404",
			7426 => x"01297531",
			7427 => x"00007531",
			7428 => x"06018108",
			7429 => x"0a02e804",
			7430 => x"fee07531",
			7431 => x"00007531",
			7432 => x"0a030808",
			7433 => x"0306ff04",
			7434 => x"00007531",
			7435 => x"00947531",
			7436 => x"00007531",
			7437 => x"0507f634",
			7438 => x"0309071c",
			7439 => x"0f09e118",
			7440 => x"0a029d0c",
			7441 => x"02093a08",
			7442 => x"0e081604",
			7443 => x"00d87531",
			7444 => x"ffc27531",
			7445 => x"fee77531",
			7446 => x"09012704",
			7447 => x"00007531",
			7448 => x"0e086804",
			7449 => x"01697531",
			7450 => x"00007531",
			7451 => x"fedb7531",
			7452 => x"0803a014",
			7453 => x"020a5010",
			7454 => x"0901df08",
			7455 => x"0f095604",
			7456 => x"00007531",
			7457 => x"00c37531",
			7458 => x"01013204",
			7459 => x"ff497531",
			7460 => x"002c7531",
			7461 => x"01387531",
			7462 => x"fff97531",
			7463 => x"05083e18",
			7464 => x"0508210c",
			7465 => x"00039604",
			7466 => x"ff017531",
			7467 => x"040c1804",
			7468 => x"01137531",
			7469 => x"00007531",
			7470 => x"09021908",
			7471 => x"030a9904",
			7472 => x"fe387531",
			7473 => x"00007531",
			7474 => x"00007531",
			7475 => x"0e0a4814",
			7476 => x"0d089a04",
			7477 => x"00007531",
			7478 => x"0c065008",
			7479 => x"00033504",
			7480 => x"00007531",
			7481 => x"013b7531",
			7482 => x"0100ff04",
			7483 => x"00437531",
			7484 => x"ffe17531",
			7485 => x"0508a310",
			7486 => x"0e0abb08",
			7487 => x"030a8104",
			7488 => x"00007531",
			7489 => x"fedf7531",
			7490 => x"05088604",
			7491 => x"006f7531",
			7492 => x"ff5d7531",
			7493 => x"030c6c08",
			7494 => x"01015c04",
			7495 => x"008d7531",
			7496 => x"00007531",
			7497 => x"0e0cf604",
			7498 => x"ff517531",
			7499 => x"00007531",
			7500 => x"0b051108",
			7501 => x"06017804",
			7502 => x"fe6c7655",
			7503 => x"fffb7655",
			7504 => x"040a5b30",
			7505 => x"03073b10",
			7506 => x"09010f08",
			7507 => x"07057704",
			7508 => x"feb67655",
			7509 => x"00007655",
			7510 => x"0d069104",
			7511 => x"00377655",
			7512 => x"00007655",
			7513 => x"0a02571c",
			7514 => x"0b06bc10",
			7515 => x"0d071608",
			7516 => x"07058b04",
			7517 => x"00007655",
			7518 => x"01e57655",
			7519 => x"03092e04",
			7520 => x"feb87655",
			7521 => x"00007655",
			7522 => x"0100fa04",
			7523 => x"fecd7655",
			7524 => x"06017504",
			7525 => x"01397655",
			7526 => x"ffa17655",
			7527 => x"01ac7655",
			7528 => x"0601793c",
			7529 => x"01008a1c",
			7530 => x"03067810",
			7531 => x"040c9308",
			7532 => x"0e061e04",
			7533 => x"fe3e7655",
			7534 => x"00007655",
			7535 => x"0c04d004",
			7536 => x"01247655",
			7537 => x"fefb7655",
			7538 => x"02093508",
			7539 => x"00042404",
			7540 => x"ff1f7655",
			7541 => x"02067655",
			7542 => x"feaf7655",
			7543 => x"040b5b10",
			7544 => x"00040208",
			7545 => x"0d064504",
			7546 => x"fdd27655",
			7547 => x"00007655",
			7548 => x"07050404",
			7549 => x"00007655",
			7550 => x"01a37655",
			7551 => x"0b054508",
			7552 => x"0900e704",
			7553 => x"fe6c7655",
			7554 => x"00007655",
			7555 => x"0003d804",
			7556 => x"00007655",
			7557 => x"fd8f7655",
			7558 => x"0c04e90c",
			7559 => x"0c04b508",
			7560 => x"01009004",
			7561 => x"01ad7655",
			7562 => x"fe6d7655",
			7563 => x"019e7655",
			7564 => x"00050810",
			7565 => x"01016008",
			7566 => x"0901d404",
			7567 => x"ffec7655",
			7568 => x"008f7655",
			7569 => x"00044304",
			7570 => x"fea77655",
			7571 => x"00827655",
			7572 => x"fe277655",
			7573 => x"0e078e60",
			7574 => x"0b056344",
			7575 => x"0d062a2c",
			7576 => x"0505f61c",
			7577 => x"0d05ed0c",
			7578 => x"040d6e04",
			7579 => x"fef37829",
			7580 => x"0b050404",
			7581 => x"00007829",
			7582 => x"00847829",
			7583 => x"0f082b08",
			7584 => x"0704ed04",
			7585 => x"00007829",
			7586 => x"00f47829",
			7587 => x"0704ef04",
			7588 => x"00007829",
			7589 => x"ff3c7829",
			7590 => x"02093d08",
			7591 => x"0c04cc04",
			7592 => x"00007829",
			7593 => x"fea97829",
			7594 => x"02096c04",
			7595 => x"00007829",
			7596 => x"fff87829",
			7597 => x"00043208",
			7598 => x"0f082204",
			7599 => x"00007829",
			7600 => x"016f7829",
			7601 => x"0e06ac08",
			7602 => x"07051c04",
			7603 => x"01397829",
			7604 => x"00007829",
			7605 => x"07051a04",
			7606 => x"feb27829",
			7607 => x"00b07829",
			7608 => x"01009708",
			7609 => x"0a02d104",
			7610 => x"fdd07829",
			7611 => x"00007829",
			7612 => x"05062608",
			7613 => x"0f085c04",
			7614 => x"ff6a7829",
			7615 => x"01547829",
			7616 => x"0900fb04",
			7617 => x"00007829",
			7618 => x"0409a004",
			7619 => x"00007829",
			7620 => x"fe8d7829",
			7621 => x"040b854c",
			7622 => x"0c056310",
			7623 => x"0b059908",
			7624 => x"0a028704",
			7625 => x"00007829",
			7626 => x"00ab7829",
			7627 => x"0100e904",
			7628 => x"fede7829",
			7629 => x"00007829",
			7630 => x"0802d420",
			7631 => x"0a021d10",
			7632 => x"02094908",
			7633 => x"0c05d704",
			7634 => x"00c47829",
			7635 => x"ff597829",
			7636 => x"01010204",
			7637 => x"00007829",
			7638 => x"01187829",
			7639 => x"040a0108",
			7640 => x"05079e04",
			7641 => x"00007829",
			7642 => x"fef87829",
			7643 => x"040a5b04",
			7644 => x"006d7829",
			7645 => x"ffab7829",
			7646 => x"0706f50c",
			7647 => x"01015c08",
			7648 => x"00037804",
			7649 => x"00007829",
			7650 => x"00ee7829",
			7651 => x"00007829",
			7652 => x"0f0b4408",
			7653 => x"09023704",
			7654 => x"ff937829",
			7655 => x"00007829",
			7656 => x"0e0b0e04",
			7657 => x"001a7829",
			7658 => x"00007829",
			7659 => x"08033128",
			7660 => x"0003ee1c",
			7661 => x"0901c30c",
			7662 => x"0a028b08",
			7663 => x"040bb004",
			7664 => x"00007829",
			7665 => x"01037829",
			7666 => x"00007829",
			7667 => x"0003dd08",
			7668 => x"0c061204",
			7669 => x"00007829",
			7670 => x"ff5b7829",
			7671 => x"0901e304",
			7672 => x"00007829",
			7673 => x"00547829",
			7674 => x"0e0aaa04",
			7675 => x"fe2b7829",
			7676 => x"0706c904",
			7677 => x"001f7829",
			7678 => x"00007829",
			7679 => x"0c050a04",
			7680 => x"ff357829",
			7681 => x"0705a104",
			7682 => x"01677829",
			7683 => x"0e0c7e08",
			7684 => x"0a02d104",
			7685 => x"00377829",
			7686 => x"ff1c7829",
			7687 => x"0004bc04",
			7688 => x"01157829",
			7689 => x"00007829",
			7690 => x"03063220",
			7691 => x"01009d1c",
			7692 => x"0208e904",
			7693 => x"fe64797d",
			7694 => x"0c04cf0c",
			7695 => x"0803be04",
			7696 => x"fe6a797d",
			7697 => x"05058404",
			7698 => x"fe9e797d",
			7699 => x"020a797d",
			7700 => x"0704ee08",
			7701 => x"0704ed04",
			7702 => x"fec8797d",
			7703 => x"0000797d",
			7704 => x"fe5a797d",
			7705 => x"01d7797d",
			7706 => x"0c066d64",
			7707 => x"0802fb30",
			7708 => x"00030210",
			7709 => x"0901a90c",
			7710 => x"0d070808",
			7711 => x"0100bf04",
			7712 => x"fe92797d",
			7713 => x"030b797d",
			7714 => x"fe68797d",
			7715 => x"011a797d",
			7716 => x"0507f510",
			7717 => x"0b06af08",
			7718 => x"0e095104",
			7719 => x"ff24797d",
			7720 => x"014f797d",
			7721 => x"07062a04",
			7722 => x"ff66797d",
			7723 => x"0197797d",
			7724 => x"0901bc08",
			7725 => x"05084d04",
			7726 => x"fe7c797d",
			7727 => x"01d5797d",
			7728 => x"00039504",
			7729 => x"fe92797d",
			7730 => x"002a797d",
			7731 => x"0901d220",
			7732 => x"0c04f110",
			7733 => x"0505cc08",
			7734 => x"040ca704",
			7735 => x"fe4e797d",
			7736 => x"0025797d",
			7737 => x"0100a804",
			7738 => x"0102797d",
			7739 => x"01dd797d",
			7740 => x"03088d08",
			7741 => x"07052f04",
			7742 => x"0041797d",
			7743 => x"fe7d797d",
			7744 => x"0c054c04",
			7745 => x"020a797d",
			7746 => x"0000797d",
			7747 => x"0b072f08",
			7748 => x"040c3204",
			7749 => x"01df797d",
			7750 => x"0000797d",
			7751 => x"0e0aaa04",
			7752 => x"fe1a797d",
			7753 => x"0c063a04",
			7754 => x"fed7797d",
			7755 => x"01e3797d",
			7756 => x"09026420",
			7757 => x"08033f1c",
			7758 => x"0d097510",
			7759 => x"01013008",
			7760 => x"01012a04",
			7761 => x"ffe6797d",
			7762 => x"065d797d",
			7763 => x"0d094e04",
			7764 => x"fe66797d",
			7765 => x"ff7f797d",
			7766 => x"0e0b0704",
			7767 => x"03e8797d",
			7768 => x"07073c04",
			7769 => x"fe8d797d",
			7770 => x"03ea797d",
			7771 => x"fe67797d",
			7772 => x"00040c04",
			7773 => x"ff32797d",
			7774 => x"0192797d",
			7775 => x"0601674c",
			7776 => x"09019624",
			7777 => x"06016318",
			7778 => x"0600e808",
			7779 => x"05064104",
			7780 => x"fe8b7b39",
			7781 => x"027d7b39",
			7782 => x"0408520c",
			7783 => x"0a01b604",
			7784 => x"fe7a7b39",
			7785 => x"05078e04",
			7786 => x"037c7b39",
			7787 => x"ff6c7b39",
			7788 => x"fe637b39",
			7789 => x"03069604",
			7790 => x"fe707b39",
			7791 => x"02091104",
			7792 => x"03487b39",
			7793 => x"feb17b39",
			7794 => x"07062b08",
			7795 => x"0e086804",
			7796 => x"01357b39",
			7797 => x"fe5e7b39",
			7798 => x"07064610",
			7799 => x"0e08cb04",
			7800 => x"fed07b39",
			7801 => x"01010204",
			7802 => x"ff2a7b39",
			7803 => x"07064004",
			7804 => x"045f7b39",
			7805 => x"02997b39",
			7806 => x"00032408",
			7807 => x"0b06cd04",
			7808 => x"01637b39",
			7809 => x"fe747b39",
			7810 => x"0c063204",
			7811 => x"03a27b39",
			7812 => x"fe9d7b39",
			7813 => x"0c066c68",
			7814 => x"0601963c",
			7815 => x"07051f1c",
			7816 => x"01009710",
			7817 => x"0f086408",
			7818 => x"0505cc04",
			7819 => x"ffec7b39",
			7820 => x"01c87b39",
			7821 => x"00043d04",
			7822 => x"fd1c7b39",
			7823 => x"fff27b39",
			7824 => x"06017404",
			7825 => x"fff27b39",
			7826 => x"0100a604",
			7827 => x"01977b39",
			7828 => x"022a7b39",
			7829 => x"03091a10",
			7830 => x"0b057408",
			7831 => x"01009904",
			7832 => x"fed87b39",
			7833 => x"023e7b39",
			7834 => x"06018d04",
			7835 => x"fe627b39",
			7836 => x"00007b39",
			7837 => x"05080408",
			7838 => x"0a024c04",
			7839 => x"00317b39",
			7840 => x"01b17b39",
			7841 => x"0901bc04",
			7842 => x"02c47b39",
			7843 => x"fed87b39",
			7844 => x"0b072f18",
			7845 => x"040c7f0c",
			7846 => x"0a027404",
			7847 => x"00007b39",
			7848 => x"09015804",
			7849 => x"01337b39",
			7850 => x"02057b39",
			7851 => x"0705a204",
			7852 => x"01e97b39",
			7853 => x"0601b304",
			7854 => x"fe3d7b39",
			7855 => x"ff7f7b39",
			7856 => x"0f0b6d08",
			7857 => x"0c066a04",
			7858 => x"fe157b39",
			7859 => x"00da7b39",
			7860 => x"0a029904",
			7861 => x"fef87b39",
			7862 => x"040ceb04",
			7863 => x"012c7b39",
			7864 => x"02377b39",
			7865 => x"09026424",
			7866 => x"0a02ac20",
			7867 => x"0901fe10",
			7868 => x"07070f08",
			7869 => x"06019904",
			7870 => x"01357b39",
			7871 => x"fe977b39",
			7872 => x"0a029304",
			7873 => x"06467b39",
			7874 => x"01377b39",
			7875 => x"0b07b508",
			7876 => x"0c066d04",
			7877 => x"002f7b39",
			7878 => x"fe737b39",
			7879 => x"040b4a04",
			7880 => x"06557b39",
			7881 => x"fe717b39",
			7882 => x"fe637b39",
			7883 => x"00040c04",
			7884 => x"feff7b39",
			7885 => x"022f7b39",
			7886 => x"0100954c",
			7887 => x"040bb214",
			7888 => x"0900f710",
			7889 => x"0f080e04",
			7890 => x"00007cfd",
			7891 => x"07051f08",
			7892 => x"0704f104",
			7893 => x"00007cfd",
			7894 => x"feb77cfd",
			7895 => x"00007cfd",
			7896 => x"00007cfd",
			7897 => x"0c04d420",
			7898 => x"0505db14",
			7899 => x"0601780c",
			7900 => x"0c049504",
			7901 => x"00007cfd",
			7902 => x"040d2e04",
			7903 => x"ff3c7cfd",
			7904 => x"00007cfd",
			7905 => x"0b051104",
			7906 => x"00007cfd",
			7907 => x"00647cfd",
			7908 => x"0d05f704",
			7909 => x"00007cfd",
			7910 => x"07050804",
			7911 => x"01107cfd",
			7912 => x"00007cfd",
			7913 => x"040e6310",
			7914 => x"0100900c",
			7915 => x"0900c204",
			7916 => x"00007cfd",
			7917 => x"0704ee04",
			7918 => x"00007cfd",
			7919 => x"fef07cfd",
			7920 => x"00007cfd",
			7921 => x"06018004",
			7922 => x"00007cfd",
			7923 => x"00477cfd",
			7924 => x"02095734",
			7925 => x"06017424",
			7926 => x"040b3c20",
			7927 => x"07063f10",
			7928 => x"0c056208",
			7929 => x"07051804",
			7930 => x"00697cfd",
			7931 => x"ff9b7cfd",
			7932 => x"01012604",
			7933 => x"00b47cfd",
			7934 => x"00007cfd",
			7935 => x"08025a08",
			7936 => x"0100f504",
			7937 => x"00007cfd",
			7938 => x"00207cfd",
			7939 => x"01011b04",
			7940 => x"ff7d7cfd",
			7941 => x"00007cfd",
			7942 => x"ff937cfd",
			7943 => x"040aa908",
			7944 => x"040a6904",
			7945 => x"00597cfd",
			7946 => x"00007cfd",
			7947 => x"0a029604",
			7948 => x"00007cfd",
			7949 => x"01587cfd",
			7950 => x"0f0ab234",
			7951 => x"020a8320",
			7952 => x"0f09b110",
			7953 => x"06018108",
			7954 => x"0c060f04",
			7955 => x"fece7cfd",
			7956 => x"00007cfd",
			7957 => x"0b057404",
			7958 => x"00d47cfd",
			7959 => x"ffcf7cfd",
			7960 => x"07064108",
			7961 => x"0d080e04",
			7962 => x"00437cfd",
			7963 => x"ff7e7cfd",
			7964 => x"0100fa04",
			7965 => x"00007cfd",
			7966 => x"00767cfd",
			7967 => x"06019f0c",
			7968 => x"06017c04",
			7969 => x"00007cfd",
			7970 => x"040aed04",
			7971 => x"00007cfd",
			7972 => x"fe997cfd",
			7973 => x"07064404",
			7974 => x"006a7cfd",
			7975 => x"00007cfd",
			7976 => x"0b073310",
			7977 => x"01011d04",
			7978 => x"00007cfd",
			7979 => x"0f0b9808",
			7980 => x"09022304",
			7981 => x"01307cfd",
			7982 => x"00007cfd",
			7983 => x"00007cfd",
			7984 => x"0601af10",
			7985 => x"0706b708",
			7986 => x"09022904",
			7987 => x"ffd37cfd",
			7988 => x"00007cfd",
			7989 => x"01015004",
			7990 => x"007d7cfd",
			7991 => x"00007cfd",
			7992 => x"030d4e08",
			7993 => x"0706f804",
			7994 => x"00007cfd",
			7995 => x"ff0d7cfd",
			7996 => x"020fae04",
			7997 => x"00017cfd",
			7998 => x"00007cfd",
			7999 => x"06016444",
			8000 => x"0901a120",
			8001 => x"0100a10c",
			8002 => x"03069604",
			8003 => x"fe637ecb",
			8004 => x"0e064304",
			8005 => x"00e57ecb",
			8006 => x"fe807ecb",
			8007 => x"0705ff10",
			8008 => x"0c056204",
			8009 => x"fe927ecb",
			8010 => x"0002f604",
			8011 => x"fece7ecb",
			8012 => x"0003d804",
			8013 => x"02b27ecb",
			8014 => x"ffa77ecb",
			8015 => x"fe5e7ecb",
			8016 => x"0a020808",
			8017 => x"0901a904",
			8018 => x"ff847ecb",
			8019 => x"03b07ecb",
			8020 => x"07062b04",
			8021 => x"fe957ecb",
			8022 => x"08029110",
			8023 => x"01010f08",
			8024 => x"01010604",
			8025 => x"000b7ecb",
			8026 => x"fee77ecb",
			8027 => x"08028704",
			8028 => x"00c67ecb",
			8029 => x"03607ecb",
			8030 => x"0a022804",
			8031 => x"fec97ecb",
			8032 => x"00337ecb",
			8033 => x"0c066d74",
			8034 => x"06017938",
			8035 => x"0208f018",
			8036 => x"0306a50c",
			8037 => x"040c0404",
			8038 => x"fe4f7ecb",
			8039 => x"0305b904",
			8040 => x"fea07ecb",
			8041 => x"022b7ecb",
			8042 => x"00042008",
			8043 => x"06017004",
			8044 => x"004b7ecb",
			8045 => x"01e97ecb",
			8046 => x"02787ecb",
			8047 => x"03091a10",
			8048 => x"0f088508",
			8049 => x"08032c04",
			8050 => x"fb937ecb",
			8051 => x"00437ecb",
			8052 => x"02091904",
			8053 => x"ffa07ecb",
			8054 => x"fe207ecb",
			8055 => x"0f097108",
			8056 => x"01012e04",
			8057 => x"032d7ecb",
			8058 => x"fec07ecb",
			8059 => x"00033e04",
			8060 => x"fe607ecb",
			8061 => x"008c7ecb",
			8062 => x"0802fb20",
			8063 => x"07066d10",
			8064 => x"040adc08",
			8065 => x"00036804",
			8066 => x"fe927ecb",
			8067 => x"01e17ecb",
			8068 => x"030a1204",
			8069 => x"fd857ecb",
			8070 => x"01c07ecb",
			8071 => x"0d08da08",
			8072 => x"0d085904",
			8073 => x"00937ecb",
			8074 => x"fe2d7ecb",
			8075 => x"0706c904",
			8076 => x"02f57ecb",
			8077 => x"ff547ecb",
			8078 => x"0e0a3910",
			8079 => x"07051f08",
			8080 => x"01009004",
			8081 => x"01157ecb",
			8082 => x"01c87ecb",
			8083 => x"08031704",
			8084 => x"01e77ecb",
			8085 => x"00097ecb",
			8086 => x"08036908",
			8087 => x"06019104",
			8088 => x"03497ecb",
			8089 => x"01ab7ecb",
			8090 => x"00637ecb",
			8091 => x"0d095014",
			8092 => x"01013010",
			8093 => x"01012a0c",
			8094 => x"0d093704",
			8095 => x"fe9c7ecb",
			8096 => x"0003dd04",
			8097 => x"01ae7ecb",
			8098 => x"ff697ecb",
			8099 => x"033d7ecb",
			8100 => x"fe6a7ecb",
			8101 => x"00039d0c",
			8102 => x"030b2a08",
			8103 => x"0c06a404",
			8104 => x"ff387ecb",
			8105 => x"01e27ecb",
			8106 => x"07fd7ecb",
			8107 => x"0004a70c",
			8108 => x"040be404",
			8109 => x"fe7d7ecb",
			8110 => x"0a029604",
			8111 => x"02967ecb",
			8112 => x"005f7ecb",
			8113 => x"fe657ecb",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(2750, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(5367, initial_addr_3'length));
	end generate gen_rom_9;

	gen_rom_10: if SELECT_ROM = 10 generate
		bank <= (
			0 => x"00000005",
			1 => x"00000009",
			2 => x"0000000d",
			3 => x"00000011",
			4 => x"00000015",
			5 => x"00000019",
			6 => x"0000001d",
			7 => x"00000021",
			8 => x"00000025",
			9 => x"00000029",
			10 => x"0000002d",
			11 => x"00000031",
			12 => x"00000035",
			13 => x"00000039",
			14 => x"0000003d",
			15 => x"00000041",
			16 => x"00000045",
			17 => x"00000049",
			18 => x"0000004d",
			19 => x"00000051",
			20 => x"0409db04",
			21 => x"00000065",
			22 => x"01014f04",
			23 => x"ffbd0065",
			24 => x"00000065",
			25 => x"06018604",
			26 => x"00000079",
			27 => x"0601bc04",
			28 => x"00110079",
			29 => x"00000079",
			30 => x"01014108",
			31 => x"0901d904",
			32 => x"0000008d",
			33 => x"0049008d",
			34 => x"0000008d",
			35 => x"01014f08",
			36 => x"0002f604",
			37 => x"000000a1",
			38 => x"ffe900a1",
			39 => x"000000a1",
			40 => x"09020808",
			41 => x"0e0abb04",
			42 => x"ffd200b5",
			43 => x"000000b5",
			44 => x"000000b5",
			45 => x"00038e0c",
			46 => x"00038504",
			47 => x"000000d1",
			48 => x"0802db04",
			49 => x"000000d1",
			50 => x"003000d1",
			51 => x"fff600d1",
			52 => x"0e0b320c",
			53 => x"01015108",
			54 => x"0e09c104",
			55 => x"000000ed",
			56 => x"ffe600ed",
			57 => x"000000ed",
			58 => x"000000ed",
			59 => x"040b0404",
			60 => x"00000109",
			61 => x"040d0008",
			62 => x"0901ce04",
			63 => x"00000109",
			64 => x"ffdb0109",
			65 => x"00000109",
			66 => x"0901f604",
			67 => x"00000125",
			68 => x"05094208",
			69 => x"09022a04",
			70 => x"00450125",
			71 => x"00000125",
			72 => x"00000125",
			73 => x"00038e0c",
			74 => x"09020804",
			75 => x"00000151",
			76 => x"0f0a5a04",
			77 => x"00530151",
			78 => x"00000151",
			79 => x"0f0b2608",
			80 => x"00039604",
			81 => x"00000151",
			82 => x"ffdb0151",
			83 => x"00000151",
			84 => x"0b06dd04",
			85 => x"00000175",
			86 => x"0601bc0c",
			87 => x"06018504",
			88 => x"00000175",
			89 => x"0b07b804",
			90 => x"00340175",
			91 => x"00000175",
			92 => x"00000175",
			93 => x"07064608",
			94 => x"0c05bb04",
			95 => x"000001a1",
			96 => x"000401a1",
			97 => x"01011d04",
			98 => x"000001a1",
			99 => x"09020808",
			100 => x"0901cc04",
			101 => x"000001a1",
			102 => x"ff9d01a1",
			103 => x"000001a1",
			104 => x"07065b10",
			105 => x"00038e0c",
			106 => x"07061404",
			107 => x"000001cd",
			108 => x"0002e604",
			109 => x"000001cd",
			110 => x"002f01cd",
			111 => x"000001cd",
			112 => x"0706a104",
			113 => x"ffc201cd",
			114 => x"000001cd",
			115 => x"0003960c",
			116 => x"09020804",
			117 => x"00000209",
			118 => x"030a3904",
			119 => x"008b0209",
			120 => x"00000209",
			121 => x"0e0ac108",
			122 => x"01015104",
			123 => x"ff740209",
			124 => x"00000209",
			125 => x"0d09db08",
			126 => x"0706a104",
			127 => x"00000209",
			128 => x"00450209",
			129 => x"00000209",
			130 => x"040abb14",
			131 => x"030a2810",
			132 => x"0c061a0c",
			133 => x"0c05bb04",
			134 => x"0000023d",
			135 => x"04090804",
			136 => x"0000023d",
			137 => x"0034023d",
			138 => x"0000023d",
			139 => x"0000023d",
			140 => x"030ae104",
			141 => x"ffeb023d",
			142 => x"0000023d",
			143 => x"0b06dd04",
			144 => x"00000269",
			145 => x"0601bc10",
			146 => x"06018504",
			147 => x"00000269",
			148 => x"05094208",
			149 => x"0507e404",
			150 => x"00000269",
			151 => x"003f0269",
			152 => x"00000269",
			153 => x"00000269",
			154 => x"0901dd10",
			155 => x"0706a10c",
			156 => x"0e0a4808",
			157 => x"06014704",
			158 => x"000002ad",
			159 => x"ffd402ad",
			160 => x"000002ad",
			161 => x"000002ad",
			162 => x"09022c10",
			163 => x"0601be0c",
			164 => x"0a023304",
			165 => x"000002ad",
			166 => x"0e08e104",
			167 => x"000002ad",
			168 => x"002f02ad",
			169 => x"000002ad",
			170 => x"000002ad",
			171 => x"07064614",
			172 => x"0c05bb04",
			173 => x"000002f1",
			174 => x"0802e30c",
			175 => x"08026904",
			176 => x"000002f1",
			177 => x"07060204",
			178 => x"000002f1",
			179 => x"001d02f1",
			180 => x"000002f1",
			181 => x"01011d04",
			182 => x"000002f1",
			183 => x"09020808",
			184 => x"0901cc04",
			185 => x"000002f1",
			186 => x"ff9302f1",
			187 => x"000002f1",
			188 => x"040abb14",
			189 => x"0e09fd10",
			190 => x"0802a504",
			191 => x"00000345",
			192 => x"0e08e104",
			193 => x"00000345",
			194 => x"00038e04",
			195 => x"00520345",
			196 => x"00000345",
			197 => x"00000345",
			198 => x"0e0ac10c",
			199 => x"0901b804",
			200 => x"00000345",
			201 => x"09021d04",
			202 => x"ffba0345",
			203 => x"00000345",
			204 => x"05096108",
			205 => x"0b073304",
			206 => x"00000345",
			207 => x"00300345",
			208 => x"00000345",
			209 => x"040aa918",
			210 => x"0e09fd14",
			211 => x"0d078804",
			212 => x"00000381",
			213 => x"0d08b30c",
			214 => x"08025f04",
			215 => x"00000381",
			216 => x"00039104",
			217 => x"00510381",
			218 => x"00000381",
			219 => x"00000381",
			220 => x"00000381",
			221 => x"0e0a8604",
			222 => x"ffd30381",
			223 => x"00000381",
			224 => x"0d09db18",
			225 => x"06016804",
			226 => x"000003b5",
			227 => x"0601be10",
			228 => x"0c05bb04",
			229 => x"000003b5",
			230 => x"00044308",
			231 => x"0a023304",
			232 => x"000003b5",
			233 => x"003103b5",
			234 => x"000003b5",
			235 => x"000003b5",
			236 => x"000003b5",
			237 => x"05083004",
			238 => x"000003e9",
			239 => x"0d09c414",
			240 => x"09021510",
			241 => x"00038c04",
			242 => x"000003e9",
			243 => x"0e0a1b04",
			244 => x"000003e9",
			245 => x"040d2e04",
			246 => x"006c03e9",
			247 => x"000003e9",
			248 => x"000003e9",
			249 => x"000003e9",
			250 => x"0d088d18",
			251 => x"0901e804",
			252 => x"00000435",
			253 => x"0e0a6d10",
			254 => x"0706720c",
			255 => x"0a027208",
			256 => x"0802aa04",
			257 => x"00000435",
			258 => x"00b60435",
			259 => x"00000435",
			260 => x"00000435",
			261 => x"00000435",
			262 => x"01011d04",
			263 => x"00000435",
			264 => x"020cab08",
			265 => x"0901cc04",
			266 => x"00000435",
			267 => x"ffc30435",
			268 => x"00000435",
			269 => x"00037814",
			270 => x"0309d810",
			271 => x"06014604",
			272 => x"00000491",
			273 => x"0d088d08",
			274 => x"0c05bb04",
			275 => x"00000491",
			276 => x"00920491",
			277 => x"00000491",
			278 => x"00000491",
			279 => x"0706860c",
			280 => x"09021208",
			281 => x"01014b04",
			282 => x"ff4b0491",
			283 => x"00000491",
			284 => x"00000491",
			285 => x"01013f0c",
			286 => x"0d09db08",
			287 => x"09017d04",
			288 => x"00000491",
			289 => x"007a0491",
			290 => x"00000491",
			291 => x"00000491",
			292 => x"0901d90c",
			293 => x"06018d08",
			294 => x"0c066604",
			295 => x"ffcb04dd",
			296 => x"000004dd",
			297 => x"000004dd",
			298 => x"0d088d18",
			299 => x"0e0a6d14",
			300 => x"0507e604",
			301 => x"000004dd",
			302 => x"00036304",
			303 => x"000004dd",
			304 => x"0c062e08",
			305 => x"0802fb04",
			306 => x"00d304dd",
			307 => x"000004dd",
			308 => x"000004dd",
			309 => x"000004dd",
			310 => x"000004dd",
			311 => x"0601850c",
			312 => x"040a0104",
			313 => x"00000529",
			314 => x"01015304",
			315 => x"ff830529",
			316 => x"00000529",
			317 => x"0c06c418",
			318 => x"00038c04",
			319 => x"00000529",
			320 => x"00040b10",
			321 => x"0b06ff04",
			322 => x"00000529",
			323 => x"0c05f604",
			324 => x"00000529",
			325 => x"0d098504",
			326 => x"00720529",
			327 => x"00000529",
			328 => x"00000529",
			329 => x"00000529",
			330 => x"0003961c",
			331 => x"0b072018",
			332 => x"0901e804",
			333 => x"0000056d",
			334 => x"07067110",
			335 => x"020a460c",
			336 => x"0507e404",
			337 => x"0000056d",
			338 => x"00036304",
			339 => x"0000056d",
			340 => x"00ad056d",
			341 => x"0000056d",
			342 => x"0000056d",
			343 => x"0000056d",
			344 => x"06019004",
			345 => x"ffc9056d",
			346 => x"0000056d",
			347 => x"0901dd14",
			348 => x"06018d08",
			349 => x"00036304",
			350 => x"000005d9",
			351 => x"ff2505d9",
			352 => x"040c3e08",
			353 => x"05086a04",
			354 => x"000005d9",
			355 => x"004c05d9",
			356 => x"000005d9",
			357 => x"0b080520",
			358 => x"01014110",
			359 => x"0a023304",
			360 => x"000005d9",
			361 => x"00033e04",
			362 => x"000005d9",
			363 => x"0e08e104",
			364 => x"000005d9",
			365 => x"00a305d9",
			366 => x"0003a308",
			367 => x"00038104",
			368 => x"000005d9",
			369 => x"ffac05d9",
			370 => x"0003f304",
			371 => x"002f05d9",
			372 => x"000005d9",
			373 => x"ffe705d9",
			374 => x"06018c04",
			375 => x"00000615",
			376 => x"0d09db18",
			377 => x"0601be14",
			378 => x"0d086604",
			379 => x"00000615",
			380 => x"0a02cb0c",
			381 => x"0b06ee04",
			382 => x"00000615",
			383 => x"0a026404",
			384 => x"00000615",
			385 => x"00460615",
			386 => x"00000615",
			387 => x"00000615",
			388 => x"00000615",
			389 => x"0b06dd08",
			390 => x"040a0104",
			391 => x"00000671",
			392 => x"ffbe0671",
			393 => x"0b07a418",
			394 => x"06017404",
			395 => x"00000671",
			396 => x"08032e10",
			397 => x"09022c0c",
			398 => x"0c05f404",
			399 => x"00000671",
			400 => x"07065804",
			401 => x"00000671",
			402 => x"00860671",
			403 => x"00000671",
			404 => x"00000671",
			405 => x"0803560c",
			406 => x"0c068b04",
			407 => x"00000671",
			408 => x"0706f804",
			409 => x"00000671",
			410 => x"ffcd0671",
			411 => x"00000671",
			412 => x"00038e14",
			413 => x"0901e804",
			414 => x"000006d5",
			415 => x"0706710c",
			416 => x"020a4608",
			417 => x"0e08e104",
			418 => x"000006d5",
			419 => x"00cf06d5",
			420 => x"000006d5",
			421 => x"000006d5",
			422 => x"07068604",
			423 => x"ff2906d5",
			424 => x"06018e08",
			425 => x"0706cc04",
			426 => x"000006d5",
			427 => x"ffca06d5",
			428 => x"0d09c410",
			429 => x"0902190c",
			430 => x"0601be08",
			431 => x"0e0a1b04",
			432 => x"000006d5",
			433 => x"009b06d5",
			434 => x"000006d5",
			435 => x"000006d5",
			436 => x"000006d5",
			437 => x"0901dd1c",
			438 => x"0e0a390c",
			439 => x"04091d04",
			440 => x"00000761",
			441 => x"0c068704",
			442 => x"ff3d0761",
			443 => x"00000761",
			444 => x"05090a0c",
			445 => x"07069b04",
			446 => x"00000761",
			447 => x"040c7f04",
			448 => x"002e0761",
			449 => x"00000761",
			450 => x"00000761",
			451 => x"0e09fd10",
			452 => x"0507e404",
			453 => x"00000761",
			454 => x"00039108",
			455 => x"00036304",
			456 => x"00000761",
			457 => x"00ab0761",
			458 => x"00000761",
			459 => x"0003a308",
			460 => x"0802e604",
			461 => x"00000761",
			462 => x"ffa40761",
			463 => x"05094f10",
			464 => x"06019404",
			465 => x"00000761",
			466 => x"05083004",
			467 => x"00000761",
			468 => x"0601be04",
			469 => x"00880761",
			470 => x"00000761",
			471 => x"00000761",
			472 => x"040af51c",
			473 => x"0d08b318",
			474 => x"06019214",
			475 => x"00038e10",
			476 => x"06014604",
			477 => x"000007d5",
			478 => x"020a4608",
			479 => x"07060204",
			480 => x"000007d5",
			481 => x"007a07d5",
			482 => x"000007d5",
			483 => x"000007d5",
			484 => x"000007d5",
			485 => x"000007d5",
			486 => x"05086a08",
			487 => x"00039604",
			488 => x"000007d5",
			489 => x"ff3607d5",
			490 => x"07070f10",
			491 => x"040c240c",
			492 => x"0a026d04",
			493 => x"000007d5",
			494 => x"09021904",
			495 => x"00b307d5",
			496 => x"000007d5",
			497 => x"000007d5",
			498 => x"0e0b0e04",
			499 => x"ffbe07d5",
			500 => x"000007d5",
			501 => x"0003d92c",
			502 => x"0c05f610",
			503 => x"0409ed0c",
			504 => x"0a023304",
			505 => x"00000859",
			506 => x"0e08e104",
			507 => x"00000859",
			508 => x"001c0859",
			509 => x"ffc40859",
			510 => x"0706ce14",
			511 => x"09022a10",
			512 => x"0d084a04",
			513 => x"00000859",
			514 => x"08030f08",
			515 => x"0a024f04",
			516 => x"00000859",
			517 => x"00aa0859",
			518 => x"00000859",
			519 => x"00000859",
			520 => x"0802fc04",
			521 => x"fff90859",
			522 => x"00000859",
			523 => x"0e0b3204",
			524 => x"ff2c0859",
			525 => x"09020e10",
			526 => x"0d09c40c",
			527 => x"030b2304",
			528 => x"00000859",
			529 => x"0004dd04",
			530 => x"00940859",
			531 => x"00000859",
			532 => x"00000859",
			533 => x"00000859",
			534 => x"040af51c",
			535 => x"0d08b318",
			536 => x"06019214",
			537 => x"06014604",
			538 => x"000008d5",
			539 => x"020a460c",
			540 => x"0a026c08",
			541 => x"07060204",
			542 => x"000008d5",
			543 => x"006e08d5",
			544 => x"000008d5",
			545 => x"000008d5",
			546 => x"000008d5",
			547 => x"000008d5",
			548 => x"0e0aee0c",
			549 => x"01011504",
			550 => x"000008d5",
			551 => x"0901bf04",
			552 => x"000008d5",
			553 => x"ff6608d5",
			554 => x"0d09db14",
			555 => x"0706a104",
			556 => x"000008d5",
			557 => x"01010604",
			558 => x"000008d5",
			559 => x"01015008",
			560 => x"0e0afd04",
			561 => x"000008d5",
			562 => x"00b008d5",
			563 => x"000008d5",
			564 => x"000008d5",
			565 => x"07067224",
			566 => x"0c05f60c",
			567 => x"0409ed04",
			568 => x"00000961",
			569 => x"01014b04",
			570 => x"ffc50961",
			571 => x"00000961",
			572 => x"0c061a14",
			573 => x"0d088d10",
			574 => x"0a02720c",
			575 => x"07063f04",
			576 => x"00000961",
			577 => x"06014604",
			578 => x"00000961",
			579 => x"00b40961",
			580 => x"00000961",
			581 => x"00000961",
			582 => x"00000961",
			583 => x"07068604",
			584 => x"ff4c0961",
			585 => x"05094f18",
			586 => x"01014510",
			587 => x"0100ff04",
			588 => x"00000961",
			589 => x"0c063204",
			590 => x"00000961",
			591 => x"05084d04",
			592 => x"00000961",
			593 => x"00930961",
			594 => x"07068804",
			595 => x"00000961",
			596 => x"ffc10961",
			597 => x"0c06a504",
			598 => x"00000961",
			599 => x"ffa40961",
			600 => x"0901f428",
			601 => x"07068508",
			602 => x"0409c704",
			603 => x"00000a0d",
			604 => x"feca0a0d",
			605 => x"0706f814",
			606 => x"040ba410",
			607 => x"0f09b104",
			608 => x"00000a0d",
			609 => x"00034b04",
			610 => x"00000a0d",
			611 => x"0508b204",
			612 => x"009e0a0d",
			613 => x"00000a0d",
			614 => x"00000a0d",
			615 => x"0f0b8808",
			616 => x"0c068a04",
			617 => x"00000a0d",
			618 => x"ff990a0d",
			619 => x"00000a0d",
			620 => x"0c06301c",
			621 => x"0003af18",
			622 => x"0507e408",
			623 => x"0c05db04",
			624 => x"002d0a0d",
			625 => x"00000a0d",
			626 => x"0c05f604",
			627 => x"00000a0d",
			628 => x"01013c04",
			629 => x"00000a0d",
			630 => x"0901fe04",
			631 => x"00000a0d",
			632 => x"012c0a0d",
			633 => x"00000a0d",
			634 => x"0101450c",
			635 => x"06019404",
			636 => x"00000a0d",
			637 => x"05086a04",
			638 => x"00000a0d",
			639 => x"008a0a0d",
			640 => x"040a9504",
			641 => x"00000a0d",
			642 => x"ff520a0d",
			643 => x"040ae224",
			644 => x"09020818",
			645 => x"06017914",
			646 => x"06014604",
			647 => x"00000ab1",
			648 => x"0101390c",
			649 => x"05084d08",
			650 => x"07061404",
			651 => x"00000ab1",
			652 => x"00ba0ab1",
			653 => x"00000ab1",
			654 => x"00000ab1",
			655 => x"ff830ab1",
			656 => x"07068508",
			657 => x"020a4604",
			658 => x"013a0ab1",
			659 => x"00000ab1",
			660 => x"00000ab1",
			661 => x"0e0b321c",
			662 => x"040be418",
			663 => x"05086a08",
			664 => x"01014b04",
			665 => x"ff780ab1",
			666 => x"00000ab1",
			667 => x"040b5604",
			668 => x"00000ab1",
			669 => x"0d094108",
			670 => x"01015104",
			671 => x"00b60ab1",
			672 => x"00000ab1",
			673 => x"00000ab1",
			674 => x"fefb0ab1",
			675 => x"0b080510",
			676 => x"0b077304",
			677 => x"00000ab1",
			678 => x"09021908",
			679 => x"01010b04",
			680 => x"00000ab1",
			681 => x"013d0ab1",
			682 => x"00000ab1",
			683 => x"ffba0ab1",
			684 => x"0100ff18",
			685 => x"00036310",
			686 => x"0a022b0c",
			687 => x"09010f08",
			688 => x"05068904",
			689 => x"fe830b55",
			690 => x"06520b55",
			691 => x"fe690b55",
			692 => x"06c30b55",
			693 => x"0100e804",
			694 => x"fe640b55",
			695 => x"fda30b55",
			696 => x"09021f34",
			697 => x"05082e1c",
			698 => x"0901fe0c",
			699 => x"0409db08",
			700 => x"06016f04",
			701 => x"fe8a0b55",
			702 => x"066c0b55",
			703 => x"fe470b55",
			704 => x"0209dd04",
			705 => x"04150b55",
			706 => x"01015108",
			707 => x"01014d04",
			708 => x"fe4c0b55",
			709 => x"00380b55",
			710 => x"06010b55",
			711 => x"0802e008",
			712 => x"0901a104",
			713 => x"00f00b55",
			714 => x"fe6e0b55",
			715 => x"020a8c04",
			716 => x"06460b55",
			717 => x"05094208",
			718 => x"06018c04",
			719 => x"fdc30b55",
			720 => x"01b40b55",
			721 => x"feaa0b55",
			722 => x"07065604",
			723 => x"00760b55",
			724 => x"fe670b55",
			725 => x"00040744",
			726 => x"0e0aee34",
			727 => x"0003b328",
			728 => x"0b073318",
			729 => x"05082e0c",
			730 => x"0309d808",
			731 => x"0901e804",
			732 => x"00000be9",
			733 => x"00750be9",
			734 => x"ff630be9",
			735 => x"07066d04",
			736 => x"00000be9",
			737 => x"040a6904",
			738 => x"00000be9",
			739 => x"012e0be9",
			740 => x"0003a308",
			741 => x"030a6904",
			742 => x"00000be9",
			743 => x"ff250be9",
			744 => x"0d090104",
			745 => x"00600be9",
			746 => x"00000be9",
			747 => x"0e0ac108",
			748 => x"09020e04",
			749 => x"ff000be9",
			750 => x"00000be9",
			751 => x"00000be9",
			752 => x"05086a04",
			753 => x"00000be9",
			754 => x"0a028504",
			755 => x"00000be9",
			756 => x"01015404",
			757 => x"011f0be9",
			758 => x"00000be9",
			759 => x"0e0b7704",
			760 => x"fee80be9",
			761 => x"00000be9",
			762 => x"0c05bb04",
			763 => x"fe770c6d",
			764 => x"0209ef20",
			765 => x"0601680c",
			766 => x"0100be08",
			767 => x"07062a04",
			768 => x"00000c6d",
			769 => x"011c0c6d",
			770 => x"fef20c6d",
			771 => x"0802d710",
			772 => x"0e09c10c",
			773 => x"0e08e104",
			774 => x"00000c6d",
			775 => x"0a023304",
			776 => x"00000c6d",
			777 => x"01470c6d",
			778 => x"00000c6d",
			779 => x"ffa50c6d",
			780 => x"0b06fe04",
			781 => x"fe810c6d",
			782 => x"0c06160c",
			783 => x"0c061204",
			784 => x"00000c6d",
			785 => x"01014704",
			786 => x"00000c6d",
			787 => x"018c0c6d",
			788 => x"0902120c",
			789 => x"07068504",
			790 => x"fe810c6d",
			791 => x"0d09db04",
			792 => x"005e0c6d",
			793 => x"fee10c6d",
			794 => x"fe6c0c6d",
			795 => x"05075604",
			796 => x"fe6a0cc9",
			797 => x"0d09db28",
			798 => x"09021f20",
			799 => x"06014604",
			800 => x"feaf0cc9",
			801 => x"0e0b3210",
			802 => x"0003d908",
			803 => x"06018e04",
			804 => x"00610cc9",
			805 => x"018c0cc9",
			806 => x"0e0b0404",
			807 => x"fe2c0cc9",
			808 => x"00000cc9",
			809 => x"00044e08",
			810 => x"05089404",
			811 => x"ffe90cc9",
			812 => x"01bb0cc9",
			813 => x"ffaf0cc9",
			814 => x"05080f04",
			815 => x"00940cc9",
			816 => x"fe940cc9",
			817 => x"fe3f0cc9",
			818 => x"05094f3c",
			819 => x"030b6330",
			820 => x"08030f28",
			821 => x"0601941c",
			822 => x"0e09c10c",
			823 => x"0309b004",
			824 => x"00000d45",
			825 => x"06017c04",
			826 => x"00a30d45",
			827 => x"00000d45",
			828 => x"06018608",
			829 => x"01010204",
			830 => x"00000d45",
			831 => x"ff320d45",
			832 => x"0f0ae304",
			833 => x"00000d45",
			834 => x"fff90d45",
			835 => x"07067104",
			836 => x"00000d45",
			837 => x"09021d04",
			838 => x"00ab0d45",
			839 => x"00000d45",
			840 => x"0e0aee04",
			841 => x"ff670d45",
			842 => x"00000d45",
			843 => x"09021908",
			844 => x"040e2304",
			845 => x"00d10d45",
			846 => x"00000d45",
			847 => x"00000d45",
			848 => x"ff8b0d45",
			849 => x"0706400c",
			850 => x"09020a04",
			851 => x"fe650dc9",
			852 => x"01014904",
			853 => x"02390dc9",
			854 => x"00000dc9",
			855 => x"0d09db34",
			856 => x"09021f2c",
			857 => x"0d087210",
			858 => x"0d07b004",
			859 => x"02be0dc9",
			860 => x"0901fe04",
			861 => x"fe710dc9",
			862 => x"06018804",
			863 => x"01d80dc9",
			864 => x"feb00dc9",
			865 => x"020abd10",
			866 => x"0b074408",
			867 => x"00034b04",
			868 => x"fee90dc9",
			869 => x"035a0dc9",
			870 => x"01010b04",
			871 => x"01060dc9",
			872 => x"fe9f0dc9",
			873 => x"0b073304",
			874 => x"fdf70dc9",
			875 => x"06019404",
			876 => x"fef80dc9",
			877 => x"01560dc9",
			878 => x"0b06ef04",
			879 => x"01480dc9",
			880 => x"fe740dc9",
			881 => x"fe380dc9",
			882 => x"0901fe40",
			883 => x"07068518",
			884 => x"00034b14",
			885 => x"0b06a510",
			886 => x"07061404",
			887 => x"00000ea5",
			888 => x"0c05bb04",
			889 => x"00000ea5",
			890 => x"07064204",
			891 => x"012a0ea5",
			892 => x"00000ea5",
			893 => x"ff7a0ea5",
			894 => x"fe750ea5",
			895 => x"0508fb18",
			896 => x"030ac510",
			897 => x"0f0aed0c",
			898 => x"06017404",
			899 => x"ffda0ea5",
			900 => x"0706cb04",
			901 => x"00cb0ea5",
			902 => x"00000ea5",
			903 => x"ff170ea5",
			904 => x"00044e04",
			905 => x"01200ea5",
			906 => x"00000ea5",
			907 => x"0a029604",
			908 => x"febe0ea5",
			909 => x"0d099c08",
			910 => x"0f0c9c04",
			911 => x"00520ea5",
			912 => x"00000ea5",
			913 => x"00000ea5",
			914 => x"030a2810",
			915 => x"0003910c",
			916 => x"0b06dd08",
			917 => x"0b06be04",
			918 => x"00bc0ea5",
			919 => x"00000ea5",
			920 => x"01c50ea5",
			921 => x"00000ea5",
			922 => x"00038d04",
			923 => x"ff1c0ea5",
			924 => x"0003d914",
			925 => x"0902180c",
			926 => x"0d087f04",
			927 => x"00000ea5",
			928 => x"0706de04",
			929 => x"01710ea5",
			930 => x"00000ea5",
			931 => x"0c061504",
			932 => x"000a0ea5",
			933 => x"ff1e0ea5",
			934 => x"0e0b6304",
			935 => x"ff180ea5",
			936 => x"00000ea5",
			937 => x"00038e2c",
			938 => x"0a025f20",
			939 => x"0e09c118",
			940 => x"06016f08",
			941 => x"0901ec04",
			942 => x"ffc70f71",
			943 => x"00000f71",
			944 => x"0802d50c",
			945 => x"0802b304",
			946 => x"00000f71",
			947 => x"03094004",
			948 => x"00000f71",
			949 => x"01100f71",
			950 => x"00000f71",
			951 => x"00038d04",
			952 => x"ff450f71",
			953 => x"00000f71",
			954 => x"06019208",
			955 => x"030a3904",
			956 => x"016a0f71",
			957 => x"00000f71",
			958 => x"00000f71",
			959 => x"0e0a3904",
			960 => x"fea50f71",
			961 => x"0b07b124",
			962 => x"0d08b314",
			963 => x"0601990c",
			964 => x"0c061204",
			965 => x"00000f71",
			966 => x"0b070e04",
			967 => x"00000f71",
			968 => x"00640f71",
			969 => x"07066e04",
			970 => x"00000f71",
			971 => x"ff1a0f71",
			972 => x"0902190c",
			973 => x"06019004",
			974 => x"00000f71",
			975 => x"08034504",
			976 => x"01190f71",
			977 => x"00000f71",
			978 => x"00000f71",
			979 => x"0601af08",
			980 => x"0d096904",
			981 => x"00000f71",
			982 => x"ff320f71",
			983 => x"09020208",
			984 => x"0901c804",
			985 => x"00000f71",
			986 => x"001c0f71",
			987 => x"00000f71",
			988 => x"0003fb48",
			989 => x"030af134",
			990 => x"0003c02c",
			991 => x"0b073318",
			992 => x"05082e0c",
			993 => x"0309d808",
			994 => x"0901e804",
			995 => x"fff3100d",
			996 => x"007b100d",
			997 => x"ff2b100d",
			998 => x"07066d04",
			999 => x"0000100d",
			1000 => x"040a6904",
			1001 => x"0000100d",
			1002 => x"013c100d",
			1003 => x"0003a30c",
			1004 => x"030a6904",
			1005 => x"0000100d",
			1006 => x"040b3604",
			1007 => x"ff05100d",
			1008 => x"0000100d",
			1009 => x"05089704",
			1010 => x"008c100d",
			1011 => x"0000100d",
			1012 => x"030ad104",
			1013 => x"fef6100d",
			1014 => x"0000100d",
			1015 => x"0a028504",
			1016 => x"0000100d",
			1017 => x"0101510c",
			1018 => x"040c5808",
			1019 => x"0003f704",
			1020 => x"011f100d",
			1021 => x"0000100d",
			1022 => x"0000100d",
			1023 => x"0000100d",
			1024 => x"0e0b6304",
			1025 => x"fecd100d",
			1026 => x"0000100d",
			1027 => x"040abb2c",
			1028 => x"06016f08",
			1029 => x"01013404",
			1030 => x"ff7810d9",
			1031 => x"000010d9",
			1032 => x"0e09fd1c",
			1033 => x"0507e410",
			1034 => x"02095708",
			1035 => x"03090f04",
			1036 => x"000010d9",
			1037 => x"000310d9",
			1038 => x"0c05d404",
			1039 => x"000010d9",
			1040 => x"ffe510d9",
			1041 => x"0a023904",
			1042 => x"000010d9",
			1043 => x"00034b04",
			1044 => x"000010d9",
			1045 => x"018410d9",
			1046 => x"0c061504",
			1047 => x"ffd510d9",
			1048 => x"000010d9",
			1049 => x"0e0a3908",
			1050 => x"09021d04",
			1051 => x"fe9c10d9",
			1052 => x"000010d9",
			1053 => x"00039d08",
			1054 => x"0e0a4804",
			1055 => x"000010d9",
			1056 => x"ff2c10d9",
			1057 => x"0b07b114",
			1058 => x"0b072f08",
			1059 => x"0a027404",
			1060 => x"002610d9",
			1061 => x"ff4610d9",
			1062 => x"040c2408",
			1063 => x"06018e04",
			1064 => x"000010d9",
			1065 => x"013210d9",
			1066 => x"000010d9",
			1067 => x"0601af0c",
			1068 => x"0d096904",
			1069 => x"000010d9",
			1070 => x"040be404",
			1071 => x"000010d9",
			1072 => x"ff3010d9",
			1073 => x"01014708",
			1074 => x"01011b04",
			1075 => x"000010d9",
			1076 => x"002c10d9",
			1077 => x"000010d9",
			1078 => x"0100fc18",
			1079 => x"0003a210",
			1080 => x"0309ef0c",
			1081 => x"0c061004",
			1082 => x"fe68119d",
			1083 => x"09016104",
			1084 => x"0684119d",
			1085 => x"fe75119d",
			1086 => x"0564119d",
			1087 => x"09017604",
			1088 => x"fe63119d",
			1089 => x"fcfe119d",
			1090 => x"09021f44",
			1091 => x"05082e20",
			1092 => x"040a9518",
			1093 => x"0901fe0c",
			1094 => x"0901e804",
			1095 => x"fe71119d",
			1096 => x"01012e04",
			1097 => x"07b6119d",
			1098 => x"ff8a119d",
			1099 => x"0e09a204",
			1100 => x"0640119d",
			1101 => x"030a0104",
			1102 => x"0177119d",
			1103 => x"fdeb119d",
			1104 => x"01015104",
			1105 => x"fe4c119d",
			1106 => x"0067119d",
			1107 => x"0802e510",
			1108 => x"0901a108",
			1109 => x"0b072f04",
			1110 => x"ffd0119d",
			1111 => x"0113119d",
			1112 => x"07072404",
			1113 => x"fe71119d",
			1114 => x"fccc119d",
			1115 => x"05094210",
			1116 => x"040b4a08",
			1117 => x"0c063404",
			1118 => x"06e6119d",
			1119 => x"0172119d",
			1120 => x"0e0abb04",
			1121 => x"0028119d",
			1122 => x"01ec119d",
			1123 => x"fe28119d",
			1124 => x"040aa904",
			1125 => x"013d119d",
			1126 => x"fe66119d",
			1127 => x"0b067a04",
			1128 => x"fe691201",
			1129 => x"0509612c",
			1130 => x"09021f24",
			1131 => x"06014604",
			1132 => x"fea11201",
			1133 => x"0003d910",
			1134 => x"06018e08",
			1135 => x"0f0aad04",
			1136 => x"00d51201",
			1137 => x"fe751201",
			1138 => x"07066e04",
			1139 => x"ff521201",
			1140 => x"02011201",
			1141 => x"0e0b0e08",
			1142 => x"0e0b0404",
			1143 => x"fdfe1201",
			1144 => x"00001201",
			1145 => x"05089404",
			1146 => x"feea1201",
			1147 => x"018e1201",
			1148 => x"0b06ee04",
			1149 => x"00951201",
			1150 => x"fe871201",
			1151 => x"fe251201",
			1152 => x"0901d930",
			1153 => x"0c061708",
			1154 => x"0f0ad704",
			1155 => x"fe9312e5",
			1156 => x"000012e5",
			1157 => x"0d097520",
			1158 => x"0100ff10",
			1159 => x"0c064d08",
			1160 => x"0100e004",
			1161 => x"005e12e5",
			1162 => x"000012e5",
			1163 => x"0e0a8c04",
			1164 => x"ff6012e5",
			1165 => x"000012e5",
			1166 => x"00038c04",
			1167 => x"000012e5",
			1168 => x"040c7f08",
			1169 => x"0a02a604",
			1170 => x"010412e5",
			1171 => x"000012e5",
			1172 => x"000012e5",
			1173 => x"0e0b2904",
			1174 => x"ff1d12e5",
			1175 => x"000012e5",
			1176 => x"0309ef1c",
			1177 => x"0507e414",
			1178 => x"040a010c",
			1179 => x"0901e804",
			1180 => x"000012e5",
			1181 => x"0e08fd04",
			1182 => x"000012e5",
			1183 => x"00f812e5",
			1184 => x"0c05db04",
			1185 => x"000012e5",
			1186 => x"ff9112e5",
			1187 => x"00036304",
			1188 => x"000012e5",
			1189 => x"01aa12e5",
			1190 => x"0802e504",
			1191 => x"ff0812e5",
			1192 => x"0802f910",
			1193 => x"09021f0c",
			1194 => x"05080404",
			1195 => x"000012e5",
			1196 => x"05086a04",
			1197 => x"014d12e5",
			1198 => x"000012e5",
			1199 => x"000012e5",
			1200 => x"0d08b304",
			1201 => x"fee412e5",
			1202 => x"040c2408",
			1203 => x"0c066604",
			1204 => x"014512e5",
			1205 => x"000012e5",
			1206 => x"0e0b6304",
			1207 => x"ffbd12e5",
			1208 => x"000012e5",
			1209 => x"01013440",
			1210 => x"0c05f708",
			1211 => x"030a8a04",
			1212 => x"fe7313d9",
			1213 => x"000013d9",
			1214 => x"040b2214",
			1215 => x"0601740c",
			1216 => x"02087e08",
			1217 => x"0408c304",
			1218 => x"000013d9",
			1219 => x"002a13d9",
			1220 => x"fef713d9",
			1221 => x"0b06f004",
			1222 => x"000013d9",
			1223 => x"015813d9",
			1224 => x"0e0b0410",
			1225 => x"0901b80c",
			1226 => x"09019604",
			1227 => x"ff1013d9",
			1228 => x"0003b704",
			1229 => x"001913d9",
			1230 => x"000013d9",
			1231 => x"fe7613d9",
			1232 => x"0b07f60c",
			1233 => x"030b1004",
			1234 => x"000013d9",
			1235 => x"0004bc04",
			1236 => x"013913d9",
			1237 => x"000013d9",
			1238 => x"0d09db04",
			1239 => x"000013d9",
			1240 => x"ff6813d9",
			1241 => x"0c066630",
			1242 => x"0d086614",
			1243 => x"06018810",
			1244 => x"040a6908",
			1245 => x"0901fe04",
			1246 => x"000013d9",
			1247 => x"019313d9",
			1248 => x"0c061004",
			1249 => x"ff9113d9",
			1250 => x"000013d9",
			1251 => x"feb113d9",
			1252 => x"00038908",
			1253 => x"0b06ff04",
			1254 => x"00ba13d9",
			1255 => x"ff1913d9",
			1256 => x"0e0a6d08",
			1257 => x"0003ab04",
			1258 => x"024e13d9",
			1259 => x"000013d9",
			1260 => x"040b2e04",
			1261 => x"fe9813d9",
			1262 => x"0d089a04",
			1263 => x"ffcc13d9",
			1264 => x"01bd13d9",
			1265 => x"01013f04",
			1266 => x"00c613d9",
			1267 => x"0e0bab04",
			1268 => x"feb713d9",
			1269 => x"000013d9",
			1270 => x"01013444",
			1271 => x"0c05f708",
			1272 => x"030a8a04",
			1273 => x"fe7714d5",
			1274 => x"000014d5",
			1275 => x"040b2218",
			1276 => x"0309c008",
			1277 => x"0f087a04",
			1278 => x"000214d5",
			1279 => x"ff1114d5",
			1280 => x"05086a0c",
			1281 => x"00034b04",
			1282 => x"000014d5",
			1283 => x"01012e04",
			1284 => x"017f14d5",
			1285 => x"000014d5",
			1286 => x"000014d5",
			1287 => x"0e0b0410",
			1288 => x"0901b80c",
			1289 => x"09019604",
			1290 => x"ff2914d5",
			1291 => x"0508b304",
			1292 => x"009b14d5",
			1293 => x"000014d5",
			1294 => x"fe9f14d5",
			1295 => x"0b07f60c",
			1296 => x"030b1004",
			1297 => x"000014d5",
			1298 => x"0004bc04",
			1299 => x"012814d5",
			1300 => x"000014d5",
			1301 => x"0d09db04",
			1302 => x"000014d5",
			1303 => x"ff8414d5",
			1304 => x"0c066630",
			1305 => x"0d085814",
			1306 => x"0a024508",
			1307 => x"0901f804",
			1308 => x"000014d5",
			1309 => x"014a14d5",
			1310 => x"09021208",
			1311 => x"01013904",
			1312 => x"000014d5",
			1313 => x"fec014d5",
			1314 => x"000014d5",
			1315 => x"0f0a5a08",
			1316 => x"09020804",
			1317 => x"000014d5",
			1318 => x"024014d5",
			1319 => x"0003a608",
			1320 => x"01015704",
			1321 => x"fea314d5",
			1322 => x"000014d5",
			1323 => x"05083004",
			1324 => x"ffa814d5",
			1325 => x"08032804",
			1326 => x"01bf14d5",
			1327 => x"000014d5",
			1328 => x"01013f04",
			1329 => x"009f14d5",
			1330 => x"0e0bab04",
			1331 => x"fed014d5",
			1332 => x"000014d5",
			1333 => x"0c05d908",
			1334 => x"01014d04",
			1335 => x"fe9315a1",
			1336 => x"000015a1",
			1337 => x"040b9d40",
			1338 => x"0a026924",
			1339 => x"0507900c",
			1340 => x"0409c708",
			1341 => x"0002e604",
			1342 => x"000015a1",
			1343 => x"012115a1",
			1344 => x"000015a1",
			1345 => x"00035308",
			1346 => x"0b06ae04",
			1347 => x"000015a1",
			1348 => x"fef315a1",
			1349 => x"020a1808",
			1350 => x"0d084a04",
			1351 => x"ffd315a1",
			1352 => x"012015a1",
			1353 => x"00038c04",
			1354 => x"ff2b15a1",
			1355 => x"000015a1",
			1356 => x"0d090d14",
			1357 => x"07066d08",
			1358 => x"07064004",
			1359 => x"000015a1",
			1360 => x"ffec15a1",
			1361 => x"0a029008",
			1362 => x"0d087204",
			1363 => x"000015a1",
			1364 => x"017d15a1",
			1365 => x"000015a1",
			1366 => x"08030604",
			1367 => x"ffc515a1",
			1368 => x"000015a1",
			1369 => x"0e0aee08",
			1370 => x"040ba404",
			1371 => x"000015a1",
			1372 => x"feca15a1",
			1373 => x"05091b10",
			1374 => x"09020e0c",
			1375 => x"05088604",
			1376 => x"000015a1",
			1377 => x"020cab04",
			1378 => x"012f15a1",
			1379 => x"000015a1",
			1380 => x"000015a1",
			1381 => x"0601b304",
			1382 => x"fef015a1",
			1383 => x"000015a1",
			1384 => x"0100fc1c",
			1385 => x"0003a218",
			1386 => x"0002e604",
			1387 => x"fe651665",
			1388 => x"0002ee04",
			1389 => x"00351665",
			1390 => x"00039e0c",
			1391 => x"00034b04",
			1392 => x"fe781665",
			1393 => x"00035304",
			1394 => x"03e51665",
			1395 => x"fe811665",
			1396 => x"00001665",
			1397 => x"fe611665",
			1398 => x"01015040",
			1399 => x"05083020",
			1400 => x"040aa91c",
			1401 => x"01013d10",
			1402 => x"0802cf08",
			1403 => x"02092804",
			1404 => x"ff601665",
			1405 => x"fe6a1665",
			1406 => x"0507ea04",
			1407 => x"fee81665",
			1408 => x"0abd1665",
			1409 => x"0802cc04",
			1410 => x"08fb1665",
			1411 => x"01014504",
			1412 => x"fef71665",
			1413 => x"02e41665",
			1414 => x"fe511665",
			1415 => x"06018c0c",
			1416 => x"0b072004",
			1417 => x"047a1665",
			1418 => x"0003a304",
			1419 => x"fe671665",
			1420 => x"fcb21665",
			1421 => x"020ac308",
			1422 => x"040b0204",
			1423 => x"00bc1665",
			1424 => x"06f91665",
			1425 => x"0b07e608",
			1426 => x"0e0a8404",
			1427 => x"feee1665",
			1428 => x"02391665",
			1429 => x"ff7b1665",
			1430 => x"030a3904",
			1431 => x"03a51665",
			1432 => x"fe621665",
			1433 => x"0c05bb04",
			1434 => x"fe751711",
			1435 => x"09020e40",
			1436 => x"0b069c10",
			1437 => x"00034b0c",
			1438 => x"06014604",
			1439 => x"00001711",
			1440 => x"07060204",
			1441 => x"00001711",
			1442 => x"01a01711",
			1443 => x"ffef1711",
			1444 => x"0b06ed18",
			1445 => x"0b06ae0c",
			1446 => x"02095708",
			1447 => x"02092404",
			1448 => x"00001711",
			1449 => x"00451711",
			1450 => x"00001711",
			1451 => x"0507ea04",
			1452 => x"feba1711",
			1453 => x"0507f404",
			1454 => x"00001711",
			1455 => x"ff631711",
			1456 => x"030a120c",
			1457 => x"06017404",
			1458 => x"ff6b1711",
			1459 => x"00038504",
			1460 => x"018d1711",
			1461 => x"00001711",
			1462 => x"07068504",
			1463 => x"fe6b1711",
			1464 => x"0d098504",
			1465 => x"00a21711",
			1466 => x"ff751711",
			1467 => x"0c061610",
			1468 => x"0c061208",
			1469 => x"0b06d204",
			1470 => x"00001711",
			1471 => x"ff551711",
			1472 => x"0003cf04",
			1473 => x"014d1711",
			1474 => x"00001711",
			1475 => x"fe6d1711",
			1476 => x"0c05bb04",
			1477 => x"fe8317dd",
			1478 => x"0901f62c",
			1479 => x"0706860c",
			1480 => x"02088b08",
			1481 => x"06014104",
			1482 => x"000017dd",
			1483 => x"00da17dd",
			1484 => x"fe8d17dd",
			1485 => x"0d098518",
			1486 => x"0e0aa210",
			1487 => x"0706e408",
			1488 => x"0003c004",
			1489 => x"00f017dd",
			1490 => x"ff7217dd",
			1491 => x"0601a204",
			1492 => x"fee417dd",
			1493 => x"000017dd",
			1494 => x"00042e04",
			1495 => x"013217dd",
			1496 => x"000017dd",
			1497 => x"01012304",
			1498 => x"feb617dd",
			1499 => x"000017dd",
			1500 => x"0c061714",
			1501 => x"09020808",
			1502 => x"06017b04",
			1503 => x"00c617dd",
			1504 => x"fef617dd",
			1505 => x"0003b308",
			1506 => x"0b06dd04",
			1507 => x"000017dd",
			1508 => x"01c417dd",
			1509 => x"ffe017dd",
			1510 => x"0802fc0c",
			1511 => x"09020e08",
			1512 => x"09020a04",
			1513 => x"ff1317dd",
			1514 => x"00a717dd",
			1515 => x"fe9417dd",
			1516 => x"0d09010c",
			1517 => x"08030f08",
			1518 => x"01014504",
			1519 => x"009b17dd",
			1520 => x"000017dd",
			1521 => x"ff3e17dd",
			1522 => x"0e0ad004",
			1523 => x"000017dd",
			1524 => x"01015104",
			1525 => x"01a117dd",
			1526 => x"000017dd",
			1527 => x"07060204",
			1528 => x"fe701891",
			1529 => x"0b068f10",
			1530 => x"0a023e0c",
			1531 => x"0409db08",
			1532 => x"0f087204",
			1533 => x"00001891",
			1534 => x"02311891",
			1535 => x"00001891",
			1536 => x"00001891",
			1537 => x"01014b30",
			1538 => x"0e0a841c",
			1539 => x"0209ef10",
			1540 => x"040a3a08",
			1541 => x"0b06ae04",
			1542 => x"00001891",
			1543 => x"fea31891",
			1544 => x"0507e404",
			1545 => x"ff481891",
			1546 => x"02001891",
			1547 => x"0c062e04",
			1548 => x"fe231891",
			1549 => x"07068804",
			1550 => x"005d1891",
			1551 => x"fee31891",
			1552 => x"0b08050c",
			1553 => x"06018e04",
			1554 => x"fee21891",
			1555 => x"0b072f04",
			1556 => x"ff011891",
			1557 => x"01291891",
			1558 => x"05096104",
			1559 => x"00001891",
			1560 => x"fe941891",
			1561 => x"0706b414",
			1562 => x"0b06ff08",
			1563 => x"06019604",
			1564 => x"00e11891",
			1565 => x"ff501891",
			1566 => x"08032808",
			1567 => x"09021f04",
			1568 => x"022b1891",
			1569 => x"00001891",
			1570 => x"00001891",
			1571 => x"fea11891",
			1572 => x"0c05d908",
			1573 => x"09021504",
			1574 => x"fe6b193d",
			1575 => x"0000193d",
			1576 => x"0d09db4c",
			1577 => x"0e0b293c",
			1578 => x"020ad120",
			1579 => x"0003a310",
			1580 => x"0e0a2a08",
			1581 => x"040a6904",
			1582 => x"001d193d",
			1583 => x"01b5193d",
			1584 => x"01013c04",
			1585 => x"0056193d",
			1586 => x"fdc5193d",
			1587 => x"09020208",
			1588 => x"0706a104",
			1589 => x"fe9a193d",
			1590 => x"00ea193d",
			1591 => x"0c065204",
			1592 => x"0272193d",
			1593 => x"fff9193d",
			1594 => x"0e0abb10",
			1595 => x"020aec08",
			1596 => x"01012104",
			1597 => x"0088193d",
			1598 => x"ff47193d",
			1599 => x"0a027a04",
			1600 => x"0000193d",
			1601 => x"fe0a193d",
			1602 => x"08030204",
			1603 => x"fea1193d",
			1604 => x"08032504",
			1605 => x"011c193d",
			1606 => x"fec0193d",
			1607 => x"0101490c",
			1608 => x"0004a708",
			1609 => x"0706a104",
			1610 => x"0000193d",
			1611 => x"01b8193d",
			1612 => x"0000193d",
			1613 => x"ff44193d",
			1614 => x"fe4b193d",
			1615 => x"0100da04",
			1616 => x"fe6819d3",
			1617 => x"09021f40",
			1618 => x"06016b04",
			1619 => x"fe8819d3",
			1620 => x"040abb1c",
			1621 => x"0507e710",
			1622 => x"0409db08",
			1623 => x"0901df04",
			1624 => x"000019d3",
			1625 => x"028819d3",
			1626 => x"09020804",
			1627 => x"fe9b19d3",
			1628 => x"003319d3",
			1629 => x"030a2808",
			1630 => x"00034b04",
			1631 => x"ff8f19d3",
			1632 => x"036219d3",
			1633 => x"ff0f19d3",
			1634 => x"0003a310",
			1635 => x"030a3908",
			1636 => x"06018804",
			1637 => x"fee919d3",
			1638 => x"017c19d3",
			1639 => x"00039d04",
			1640 => x"fde019d3",
			1641 => x"ffdb19d3",
			1642 => x"0003b308",
			1643 => x"0a026c04",
			1644 => x"fef919d3",
			1645 => x"02bb19d3",
			1646 => x"05086a04",
			1647 => x"fe4919d3",
			1648 => x"00d419d3",
			1649 => x"0d085b04",
			1650 => x"009519d3",
			1651 => x"fe8119d3",
			1652 => x"000019d5",
			1653 => x"000019d9",
			1654 => x"000019dd",
			1655 => x"000019e1",
			1656 => x"000019e5",
			1657 => x"000019e9",
			1658 => x"000019ed",
			1659 => x"000019f1",
			1660 => x"000019f5",
			1661 => x"000019f9",
			1662 => x"000019fd",
			1663 => x"00001a01",
			1664 => x"00001a05",
			1665 => x"00001a09",
			1666 => x"00001a0d",
			1667 => x"00001a11",
			1668 => x"00001a15",
			1669 => x"00001a19",
			1670 => x"00001a1d",
			1671 => x"00001a21",
			1672 => x"06018604",
			1673 => x"00001a35",
			1674 => x"0601bc04",
			1675 => x"00131a35",
			1676 => x"00001a35",
			1677 => x"0e0b3208",
			1678 => x"030a0104",
			1679 => x"00001a49",
			1680 => x"fff11a49",
			1681 => x"00001a49",
			1682 => x"06018c04",
			1683 => x"00001a5d",
			1684 => x"0601be04",
			1685 => x"00171a5d",
			1686 => x"00001a5d",
			1687 => x"08033608",
			1688 => x"0802aa04",
			1689 => x"00001a71",
			1690 => x"00051a71",
			1691 => x"00001a71",
			1692 => x"07068608",
			1693 => x"07065b04",
			1694 => x"00001a8d",
			1695 => x"ffe41a8d",
			1696 => x"07070c04",
			1697 => x"003b1a8d",
			1698 => x"00001a8d",
			1699 => x"00038e0c",
			1700 => x"00038504",
			1701 => x"00001aa9",
			1702 => x"0802db04",
			1703 => x"00001aa9",
			1704 => x"002f1aa9",
			1705 => x"fff61aa9",
			1706 => x"0d09db0c",
			1707 => x"0b072f04",
			1708 => x"00001ac5",
			1709 => x"0d089a04",
			1710 => x"00001ac5",
			1711 => x"00191ac5",
			1712 => x"00001ac5",
			1713 => x"01014f0c",
			1714 => x"07067104",
			1715 => x"00001ae1",
			1716 => x"00041404",
			1717 => x"ffe11ae1",
			1718 => x"00001ae1",
			1719 => x"00001ae1",
			1720 => x"0901f604",
			1721 => x"00001afd",
			1722 => x"05094208",
			1723 => x"09022a04",
			1724 => x"003d1afd",
			1725 => x"00001afd",
			1726 => x"00001afd",
			1727 => x"0003d910",
			1728 => x"0901fe04",
			1729 => x"00001b21",
			1730 => x"0c063a08",
			1731 => x"0a027004",
			1732 => x"003b1b21",
			1733 => x"00001b21",
			1734 => x"00001b21",
			1735 => x"ffeb1b21",
			1736 => x"030b6310",
			1737 => x"040aa904",
			1738 => x"00001b45",
			1739 => x"01015108",
			1740 => x"01011f04",
			1741 => x"00001b45",
			1742 => x"ffad1b45",
			1743 => x"00001b45",
			1744 => x"00001b45",
			1745 => x"040b0410",
			1746 => x"0901e804",
			1747 => x"00001b71",
			1748 => x"030a8108",
			1749 => x"0a023304",
			1750 => x"00001b71",
			1751 => x"00241b71",
			1752 => x"00001b71",
			1753 => x"0901ca04",
			1754 => x"00001b71",
			1755 => x"ffdd1b71",
			1756 => x"00038e10",
			1757 => x"0f0a5a0c",
			1758 => x"0802aa04",
			1759 => x"00001b9d",
			1760 => x"0f091504",
			1761 => x"00001b9d",
			1762 => x"002c1b9d",
			1763 => x"00001b9d",
			1764 => x"020cab04",
			1765 => x"ffdb1b9d",
			1766 => x"00001b9d",
			1767 => x"0003960c",
			1768 => x"09020804",
			1769 => x"00001bd9",
			1770 => x"020a3a04",
			1771 => x"008e1bd9",
			1772 => x"00001bd9",
			1773 => x"0e0ac108",
			1774 => x"01015104",
			1775 => x"ff7e1bd9",
			1776 => x"00001bd9",
			1777 => x"0d09db08",
			1778 => x"0706a104",
			1779 => x"00001bd9",
			1780 => x"00451bd9",
			1781 => x"00001bd9",
			1782 => x"07065b14",
			1783 => x"00038e10",
			1784 => x"030a120c",
			1785 => x"07061404",
			1786 => x"00001c0d",
			1787 => x"0002e604",
			1788 => x"00001c0d",
			1789 => x"00431c0d",
			1790 => x"00001c0d",
			1791 => x"00001c0d",
			1792 => x"0706a104",
			1793 => x"ffc71c0d",
			1794 => x"00001c0d",
			1795 => x"0901fc04",
			1796 => x"00001c39",
			1797 => x"0c066610",
			1798 => x"0601b20c",
			1799 => x"09022d08",
			1800 => x"0901fe04",
			1801 => x"00001c39",
			1802 => x"00421c39",
			1803 => x"00001c39",
			1804 => x"00001c39",
			1805 => x"00001c39",
			1806 => x"0802ed14",
			1807 => x"0507ea04",
			1808 => x"00001c7d",
			1809 => x"00035b04",
			1810 => x"00001c7d",
			1811 => x"0b072008",
			1812 => x"020a4604",
			1813 => x"008b1c7d",
			1814 => x"00001c7d",
			1815 => x"00001c7d",
			1816 => x"0e0ac10c",
			1817 => x"01015108",
			1818 => x"040af504",
			1819 => x"00001c7d",
			1820 => x"ff8d1c7d",
			1821 => x"00001c7d",
			1822 => x"00001c7d",
			1823 => x"0802ed18",
			1824 => x"0507ea08",
			1825 => x"0002f604",
			1826 => x"00001cd1",
			1827 => x"fffa1cd1",
			1828 => x"00035b04",
			1829 => x"00001cd1",
			1830 => x"030a8108",
			1831 => x"0706b404",
			1832 => x"00721cd1",
			1833 => x"00001cd1",
			1834 => x"00001cd1",
			1835 => x"05086a08",
			1836 => x"040a9504",
			1837 => x"00001cd1",
			1838 => x"ff9b1cd1",
			1839 => x"040c2408",
			1840 => x"040b5604",
			1841 => x"00001cd1",
			1842 => x"004f1cd1",
			1843 => x"00001cd1",
			1844 => x"040aa918",
			1845 => x"0e09fd14",
			1846 => x"07061404",
			1847 => x"00001d0d",
			1848 => x"08025f04",
			1849 => x"00001d0d",
			1850 => x"0d08b308",
			1851 => x"0a026c04",
			1852 => x"00611d0d",
			1853 => x"00001d0d",
			1854 => x"00001d0d",
			1855 => x"00001d0d",
			1856 => x"0e0a8604",
			1857 => x"ffc91d0d",
			1858 => x"00001d0d",
			1859 => x"08030f18",
			1860 => x"06016804",
			1861 => x"00001d49",
			1862 => x"0d090110",
			1863 => x"020b080c",
			1864 => x"0507ea04",
			1865 => x"00001d49",
			1866 => x"0802b704",
			1867 => x"00001d49",
			1868 => x"004a1d49",
			1869 => x"00001d49",
			1870 => x"00001d49",
			1871 => x"020cab04",
			1872 => x"fff81d49",
			1873 => x"00001d49",
			1874 => x"0d09db18",
			1875 => x"0100fc04",
			1876 => x"00001d7d",
			1877 => x"07068304",
			1878 => x"00001d7d",
			1879 => x"0101450c",
			1880 => x"0d089a04",
			1881 => x"00001d7d",
			1882 => x"06018d04",
			1883 => x"00001d7d",
			1884 => x"00901d7d",
			1885 => x"00001d7d",
			1886 => x"00001d7d",
			1887 => x"05083004",
			1888 => x"00001db1",
			1889 => x"0d09c414",
			1890 => x"09021510",
			1891 => x"0d088d04",
			1892 => x"00001db1",
			1893 => x"06017404",
			1894 => x"00001db1",
			1895 => x"0a02cb04",
			1896 => x"005b1db1",
			1897 => x"00001db1",
			1898 => x"00001db1",
			1899 => x"00001db1",
			1900 => x"00039618",
			1901 => x"0b072014",
			1902 => x"0c063210",
			1903 => x"06014604",
			1904 => x"00001dfd",
			1905 => x"0c05d904",
			1906 => x"00001dfd",
			1907 => x"020a4604",
			1908 => x"00671dfd",
			1909 => x"00001dfd",
			1910 => x"00001dfd",
			1911 => x"00001dfd",
			1912 => x"06019004",
			1913 => x"ffd01dfd",
			1914 => x"0a02a108",
			1915 => x"0a027504",
			1916 => x"00001dfd",
			1917 => x"002d1dfd",
			1918 => x"00001dfd",
			1919 => x"07067220",
			1920 => x"0c05f60c",
			1921 => x"0409ed04",
			1922 => x"00001e59",
			1923 => x"01014b04",
			1924 => x"ffbb1e59",
			1925 => x"00001e59",
			1926 => x"0c061a10",
			1927 => x"0003af0c",
			1928 => x"07063f04",
			1929 => x"00001e59",
			1930 => x"06014604",
			1931 => x"00001e59",
			1932 => x"00a81e59",
			1933 => x"00001e59",
			1934 => x"00001e59",
			1935 => x"020cab0c",
			1936 => x"01011d04",
			1937 => x"00001e59",
			1938 => x"0601af04",
			1939 => x"ff651e59",
			1940 => x"00001e59",
			1941 => x"00001e59",
			1942 => x"040c2420",
			1943 => x"0b06dd08",
			1944 => x"040a0104",
			1945 => x"00001ea5",
			1946 => x"ffca1ea5",
			1947 => x"07070f14",
			1948 => x"06017404",
			1949 => x"00001ea5",
			1950 => x"09022c0c",
			1951 => x"0c05f404",
			1952 => x"00001ea5",
			1953 => x"08032e04",
			1954 => x"008f1ea5",
			1955 => x"00001ea5",
			1956 => x"00001ea5",
			1957 => x"00001ea5",
			1958 => x"0a02b604",
			1959 => x"ffcc1ea5",
			1960 => x"00001ea5",
			1961 => x"0c061108",
			1962 => x"0e0a5104",
			1963 => x"ff4d1ee9",
			1964 => x"00001ee9",
			1965 => x"0d09db18",
			1966 => x"0b06ff04",
			1967 => x"00001ee9",
			1968 => x"040aa904",
			1969 => x"00001ee9",
			1970 => x"0b07a40c",
			1971 => x"040c1808",
			1972 => x"0d088204",
			1973 => x"00001ee9",
			1974 => x"007d1ee9",
			1975 => x"00001ee9",
			1976 => x"00001ee9",
			1977 => x"ffe01ee9",
			1978 => x"00038e14",
			1979 => x"0901e804",
			1980 => x"00001f4d",
			1981 => x"0706710c",
			1982 => x"020a4608",
			1983 => x"0e08e104",
			1984 => x"00001f4d",
			1985 => x"00df1f4d",
			1986 => x"00001f4d",
			1987 => x"00001f4d",
			1988 => x"07068604",
			1989 => x"ff1e1f4d",
			1990 => x"0706ce0c",
			1991 => x"08033008",
			1992 => x"09021904",
			1993 => x"009a1f4d",
			1994 => x"00001f4d",
			1995 => x"00001f4d",
			1996 => x"0601a108",
			1997 => x"040b4204",
			1998 => x"00001f4d",
			1999 => x"ffac1f4d",
			2000 => x"0601be04",
			2001 => x"00121f4d",
			2002 => x"00001f4d",
			2003 => x"0802c314",
			2004 => x"0a023304",
			2005 => x"00001fc1",
			2006 => x"0a02450c",
			2007 => x"06017c08",
			2008 => x"06016804",
			2009 => x"00001fc1",
			2010 => x"001d1fc1",
			2011 => x"00001fc1",
			2012 => x"00001fc1",
			2013 => x"06018e0c",
			2014 => x"09021208",
			2015 => x"01010204",
			2016 => x"00001fc1",
			2017 => x"ff231fc1",
			2018 => x"00001fc1",
			2019 => x"040c1210",
			2020 => x"07066d04",
			2021 => x"00001fc1",
			2022 => x"08032508",
			2023 => x"0a026a04",
			2024 => x"00001fc1",
			2025 => x"00661fc1",
			2026 => x"00001fc1",
			2027 => x"0a02ab08",
			2028 => x"040c2404",
			2029 => x"00001fc1",
			2030 => x"ffb61fc1",
			2031 => x"00001fc1",
			2032 => x"07067220",
			2033 => x"0802f618",
			2034 => x"0c061a14",
			2035 => x"0c05f604",
			2036 => x"00002035",
			2037 => x"0601920c",
			2038 => x"07063f04",
			2039 => x"00002035",
			2040 => x"06014604",
			2041 => x"00002035",
			2042 => x"00a22035",
			2043 => x"00002035",
			2044 => x"00002035",
			2045 => x"0b072004",
			2046 => x"fff52035",
			2047 => x"00002035",
			2048 => x"0e0a760c",
			2049 => x"01014b08",
			2050 => x"0706a104",
			2051 => x"ff262035",
			2052 => x"00002035",
			2053 => x"00002035",
			2054 => x"0b08050c",
			2055 => x"07068604",
			2056 => x"00002035",
			2057 => x"05083004",
			2058 => x"00002035",
			2059 => x"00442035",
			2060 => x"ffb52035",
			2061 => x"0901dd0c",
			2062 => x"0c061708",
			2063 => x"0e0a5104",
			2064 => x"ff2520a1",
			2065 => x"000020a1",
			2066 => x"000020a1",
			2067 => x"0c05f810",
			2068 => x"0802eb0c",
			2069 => x"0901e804",
			2070 => x"000020a1",
			2071 => x"0e08e104",
			2072 => x"000020a1",
			2073 => x"00d020a1",
			2074 => x"000020a1",
			2075 => x"06018e08",
			2076 => x"0309ef04",
			2077 => x"000020a1",
			2078 => x"ff7b20a1",
			2079 => x"0b080510",
			2080 => x"05083e04",
			2081 => x"000020a1",
			2082 => x"0e0a6304",
			2083 => x"000020a1",
			2084 => x"0a02c704",
			2085 => x"00d920a1",
			2086 => x"000020a1",
			2087 => x"ffeb20a1",
			2088 => x"0802f61c",
			2089 => x"0d08b314",
			2090 => x"0c05f604",
			2091 => x"00002115",
			2092 => x"0d084a04",
			2093 => x"00002115",
			2094 => x"00037004",
			2095 => x"00002115",
			2096 => x"06019104",
			2097 => x"00ed2115",
			2098 => x"00002115",
			2099 => x"06018c04",
			2100 => x"ffab2115",
			2101 => x"00002115",
			2102 => x"07068504",
			2103 => x"ff292115",
			2104 => x"01014714",
			2105 => x"01011b08",
			2106 => x"0508f804",
			2107 => x"00002115",
			2108 => x"ffe42115",
			2109 => x"0e0a5a04",
			2110 => x"00002115",
			2111 => x"05084d04",
			2112 => x"00002115",
			2113 => x"00c12115",
			2114 => x"0f0aed04",
			2115 => x"00002115",
			2116 => x"ffcf2115",
			2117 => x"0802c314",
			2118 => x"0a023304",
			2119 => x"00002191",
			2120 => x"0a02450c",
			2121 => x"06017c08",
			2122 => x"06016804",
			2123 => x"00002191",
			2124 => x"001f2191",
			2125 => x"00002191",
			2126 => x"00002191",
			2127 => x"06018e0c",
			2128 => x"09021208",
			2129 => x"0901a104",
			2130 => x"00002191",
			2131 => x"ff172191",
			2132 => x"00002191",
			2133 => x"0003d914",
			2134 => x"07066d04",
			2135 => x"00002191",
			2136 => x"0003a304",
			2137 => x"00002191",
			2138 => x"05083004",
			2139 => x"00002191",
			2140 => x"0802f104",
			2141 => x"00002191",
			2142 => x"00852191",
			2143 => x"00041808",
			2144 => x"0a02b904",
			2145 => x"ffb02191",
			2146 => x"00002191",
			2147 => x"00002191",
			2148 => x"0802f628",
			2149 => x"07065a14",
			2150 => x"0901e804",
			2151 => x"0000221d",
			2152 => x"0003910c",
			2153 => x"030a1208",
			2154 => x"0e08e104",
			2155 => x"0000221d",
			2156 => x"00d4221d",
			2157 => x"0000221d",
			2158 => x"0000221d",
			2159 => x"0003a30c",
			2160 => x"0706a108",
			2161 => x"0b06be04",
			2162 => x"0000221d",
			2163 => x"ff57221d",
			2164 => x"0000221d",
			2165 => x"0e0a9404",
			2166 => x"009c221d",
			2167 => x"0000221d",
			2168 => x"07068504",
			2169 => x"ff1b221d",
			2170 => x"01014714",
			2171 => x"01011b08",
			2172 => x"0508f804",
			2173 => x"0000221d",
			2174 => x"ffd7221d",
			2175 => x"0e0a5a04",
			2176 => x"0000221d",
			2177 => x"05084d04",
			2178 => x"0000221d",
			2179 => x"00cc221d",
			2180 => x"0f0aed04",
			2181 => x"0000221d",
			2182 => x"ffc6221d",
			2183 => x"01012a10",
			2184 => x"0e0a390c",
			2185 => x"04091d04",
			2186 => x"000022a1",
			2187 => x"0c068704",
			2188 => x"ff2422a1",
			2189 => x"000022a1",
			2190 => x"000022a1",
			2191 => x"0e09fd10",
			2192 => x"07064404",
			2193 => x"000022a1",
			2194 => x"00036304",
			2195 => x"000022a1",
			2196 => x"00038e04",
			2197 => x"00c222a1",
			2198 => x"000022a1",
			2199 => x"0003a308",
			2200 => x"0802e604",
			2201 => x"000022a1",
			2202 => x"ff9322a1",
			2203 => x"0706ce10",
			2204 => x"040c240c",
			2205 => x"0d087f04",
			2206 => x"000022a1",
			2207 => x"07066d04",
			2208 => x"000022a1",
			2209 => x"00a522a1",
			2210 => x"000022a1",
			2211 => x"040c2c08",
			2212 => x"0706e004",
			2213 => x"000022a1",
			2214 => x"ff7422a1",
			2215 => x"000022a1",
			2216 => x"040aa910",
			2217 => x"0e09fd0c",
			2218 => x"0b06ef08",
			2219 => x"0901f604",
			2220 => x"0000230d",
			2221 => x"00fa230d",
			2222 => x"0000230d",
			2223 => x"0000230d",
			2224 => x"05083004",
			2225 => x"fef2230d",
			2226 => x"0b080520",
			2227 => x"0003a30c",
			2228 => x"0e0a4804",
			2229 => x"0000230d",
			2230 => x"00039d04",
			2231 => x"ffb3230d",
			2232 => x"0000230d",
			2233 => x"0e0a5104",
			2234 => x"0000230d",
			2235 => x"0003f308",
			2236 => x"09021b04",
			2237 => x"00f0230d",
			2238 => x"0000230d",
			2239 => x"0e0b6304",
			2240 => x"ffb6230d",
			2241 => x"006c230d",
			2242 => x"ff72230d",
			2243 => x"07065814",
			2244 => x"0409ed0c",
			2245 => x"0a01fa04",
			2246 => x"000023b9",
			2247 => x"0c05bb04",
			2248 => x"000023b9",
			2249 => x"003f23b9",
			2250 => x"09021b04",
			2251 => x"feb523b9",
			2252 => x"000023b9",
			2253 => x"0c063418",
			2254 => x"0b06f008",
			2255 => x"0309c004",
			2256 => x"000023b9",
			2257 => x"ffb323b9",
			2258 => x"08030808",
			2259 => x"040a6904",
			2260 => x"000023b9",
			2261 => x"014423b9",
			2262 => x"0c063204",
			2263 => x"ffef23b9",
			2264 => x"000023b9",
			2265 => x"0e0afd18",
			2266 => x"0901ca0c",
			2267 => x"040bca08",
			2268 => x"040af704",
			2269 => x"000023b9",
			2270 => x"003123b9",
			2271 => x"ffb223b9",
			2272 => x"05083e04",
			2273 => x"000023b9",
			2274 => x"0e0ac904",
			2275 => x"ff1123b9",
			2276 => x"000023b9",
			2277 => x"0b07f610",
			2278 => x"08034c0c",
			2279 => x"09021908",
			2280 => x"040baa04",
			2281 => x"000023b9",
			2282 => x"013b23b9",
			2283 => x"000023b9",
			2284 => x"000023b9",
			2285 => x"ffe823b9",
			2286 => x"0901f418",
			2287 => x"0e0abb08",
			2288 => x"0003ab04",
			2289 => x"0000243d",
			2290 => x"ff00243d",
			2291 => x"040caf0c",
			2292 => x"0003c404",
			2293 => x"0000243d",
			2294 => x"05088604",
			2295 => x"0000243d",
			2296 => x"005f243d",
			2297 => x"0000243d",
			2298 => x"0c06e328",
			2299 => x"0b06dd08",
			2300 => x"040a5b04",
			2301 => x"0000243d",
			2302 => x"ffb9243d",
			2303 => x"00037004",
			2304 => x"0000243d",
			2305 => x"0e0a6d0c",
			2306 => x"07068808",
			2307 => x"0c05f404",
			2308 => x"0000243d",
			2309 => x"0116243d",
			2310 => x"0000243d",
			2311 => x"0e0b5108",
			2312 => x"09020a04",
			2313 => x"0000243d",
			2314 => x"ff85243d",
			2315 => x"09021904",
			2316 => x"00ec243d",
			2317 => x"0000243d",
			2318 => x"ffb9243d",
			2319 => x"0901f42c",
			2320 => x"07068508",
			2321 => x"0409c704",
			2322 => x"000024f1",
			2323 => x"febc24f1",
			2324 => x"0b07a414",
			2325 => x"040ba410",
			2326 => x"0f09b104",
			2327 => x"000024f1",
			2328 => x"0802b704",
			2329 => x"000024f1",
			2330 => x"0508b304",
			2331 => x"00b524f1",
			2332 => x"000024f1",
			2333 => x"000024f1",
			2334 => x"0c068b04",
			2335 => x"000024f1",
			2336 => x"08033f08",
			2337 => x"0706f804",
			2338 => x"000024f1",
			2339 => x"ff9724f1",
			2340 => x"000024f1",
			2341 => x"0c06301c",
			2342 => x"0003af18",
			2343 => x"0507e408",
			2344 => x"0c05db04",
			2345 => x"004024f1",
			2346 => x"000024f1",
			2347 => x"0c05f604",
			2348 => x"000024f1",
			2349 => x"01013c04",
			2350 => x"000024f1",
			2351 => x"0901fe04",
			2352 => x"000024f1",
			2353 => x"014a24f1",
			2354 => x"000024f1",
			2355 => x"0101450c",
			2356 => x"06019404",
			2357 => x"000024f1",
			2358 => x"05086a04",
			2359 => x"000024f1",
			2360 => x"009b24f1",
			2361 => x"0b072004",
			2362 => x"000024f1",
			2363 => x"ff2324f1",
			2364 => x"0e08fd10",
			2365 => x"07064304",
			2366 => x"fe6e2575",
			2367 => x"07064408",
			2368 => x"0d07fd04",
			2369 => x"00e22575",
			2370 => x"00002575",
			2371 => x"ff212575",
			2372 => x"0d09db30",
			2373 => x"0e0b511c",
			2374 => x"08032614",
			2375 => x"0a023304",
			2376 => x"fede2575",
			2377 => x"0209e808",
			2378 => x"06017904",
			2379 => x"01ca2575",
			2380 => x"00002575",
			2381 => x"0003a304",
			2382 => x"ff462575",
			2383 => x"00a92575",
			2384 => x"0e0b3204",
			2385 => x"feab2575",
			2386 => x"00002575",
			2387 => x"08036510",
			2388 => x"040c0c04",
			2389 => x"00002575",
			2390 => x"01015308",
			2391 => x"0d092904",
			2392 => x"03df2575",
			2393 => x"01a12575",
			2394 => x"00002575",
			2395 => x"00002575",
			2396 => x"fe9b2575",
			2397 => x"00038e18",
			2398 => x"01012c04",
			2399 => x"00002609",
			2400 => x"07067110",
			2401 => x"020a460c",
			2402 => x"0a023304",
			2403 => x"00002609",
			2404 => x"0e08e104",
			2405 => x"00002609",
			2406 => x"00e72609",
			2407 => x"00002609",
			2408 => x"00002609",
			2409 => x"07068604",
			2410 => x"ff122609",
			2411 => x"0706ce10",
			2412 => x"0803300c",
			2413 => x"0802ed04",
			2414 => x"00002609",
			2415 => x"01015104",
			2416 => x"00b12609",
			2417 => x"00002609",
			2418 => x"00002609",
			2419 => x"0e0afd10",
			2420 => x"040b4204",
			2421 => x"00002609",
			2422 => x"0601a608",
			2423 => x"0c06c604",
			2424 => x"ff9d2609",
			2425 => x"00002609",
			2426 => x"00002609",
			2427 => x"0d09c40c",
			2428 => x"0601be08",
			2429 => x"06019a04",
			2430 => x"00002609",
			2431 => x"00842609",
			2432 => x"00002609",
			2433 => x"00002609",
			2434 => x"040aa91c",
			2435 => x"0e09fd18",
			2436 => x"06014604",
			2437 => x"0000268d",
			2438 => x"0b06ef10",
			2439 => x"0901fe0c",
			2440 => x"02094d08",
			2441 => x"00034b04",
			2442 => x"0056268d",
			2443 => x"0000268d",
			2444 => x"0000268d",
			2445 => x"0104268d",
			2446 => x"0000268d",
			2447 => x"0000268d",
			2448 => x"06018504",
			2449 => x"fef7268d",
			2450 => x"0b080520",
			2451 => x"05086a10",
			2452 => x"040b4a0c",
			2453 => x"09021508",
			2454 => x"0d088d04",
			2455 => x"0000268d",
			2456 => x"007d268d",
			2457 => x"0000268d",
			2458 => x"ffb0268d",
			2459 => x"0601be0c",
			2460 => x"09021908",
			2461 => x"0100fc04",
			2462 => x"0000268d",
			2463 => x"00b9268d",
			2464 => x"0000268d",
			2465 => x"0000268d",
			2466 => x"ff87268d",
			2467 => x"0c061420",
			2468 => x"01012c08",
			2469 => x"0e0a6d04",
			2470 => x"ff142721",
			2471 => x"00002721",
			2472 => x"0b06f008",
			2473 => x"0b06ae04",
			2474 => x"00002721",
			2475 => x"ffd32721",
			2476 => x"0b07100c",
			2477 => x"01014d08",
			2478 => x"0507f504",
			2479 => x"00002721",
			2480 => x"00532721",
			2481 => x"00002721",
			2482 => x"00002721",
			2483 => x"05094f28",
			2484 => x"01015624",
			2485 => x"00035b04",
			2486 => x"00002721",
			2487 => x"0706ce10",
			2488 => x"06019908",
			2489 => x"040ba404",
			2490 => x"00d92721",
			2491 => x"00002721",
			2492 => x"0b074404",
			2493 => x"00002721",
			2494 => x"00032721",
			2495 => x"0e0afd08",
			2496 => x"06019004",
			2497 => x"ffa62721",
			2498 => x"00002721",
			2499 => x"0601be04",
			2500 => x"009d2721",
			2501 => x"00002721",
			2502 => x"00002721",
			2503 => x"ff752721",
			2504 => x"0901f42c",
			2505 => x"0c061008",
			2506 => x"0409c704",
			2507 => x"000027cd",
			2508 => x"ff3427cd",
			2509 => x"020a830c",
			2510 => x"08025f04",
			2511 => x"000027cd",
			2512 => x"040b0404",
			2513 => x"001d27cd",
			2514 => x"000027cd",
			2515 => x"0e0abb08",
			2516 => x"0f0aed04",
			2517 => x"000027cd",
			2518 => x"ff7c27cd",
			2519 => x"030c6c0c",
			2520 => x"0e0ae104",
			2521 => x"000027cd",
			2522 => x"0f0c9c04",
			2523 => x"004427cd",
			2524 => x"000027cd",
			2525 => x"000027cd",
			2526 => x"0c06e328",
			2527 => x"0b06dd08",
			2528 => x"040a5b04",
			2529 => x"000027cd",
			2530 => x"ffc627cd",
			2531 => x"040a9504",
			2532 => x"000027cd",
			2533 => x"0e0a6d0c",
			2534 => x"07068808",
			2535 => x"0c05f604",
			2536 => x"000027cd",
			2537 => x"011a27cd",
			2538 => x"000027cd",
			2539 => x"0e0b5108",
			2540 => x"01014904",
			2541 => x"000027cd",
			2542 => x"ff6527cd",
			2543 => x"01015104",
			2544 => x"00d527cd",
			2545 => x"000027cd",
			2546 => x"ffc527cd",
			2547 => x"0c05bb04",
			2548 => x"febd2851",
			2549 => x"0c06c434",
			2550 => x"030b5b28",
			2551 => x"07065a10",
			2552 => x"00038e0c",
			2553 => x"0901e804",
			2554 => x"00002851",
			2555 => x"030a1204",
			2556 => x"01272851",
			2557 => x"00002851",
			2558 => x"ff9f2851",
			2559 => x"040be410",
			2560 => x"07069b08",
			2561 => x"09020a04",
			2562 => x"fecb2851",
			2563 => x"00232851",
			2564 => x"09020a04",
			2565 => x"00c32851",
			2566 => x"ffd52851",
			2567 => x"0e0afd04",
			2568 => x"fefb2851",
			2569 => x"00002851",
			2570 => x"09021908",
			2571 => x"0004a004",
			2572 => x"01352851",
			2573 => x"00002851",
			2574 => x"00002851",
			2575 => x"07070f04",
			2576 => x"00002851",
			2577 => x"0a02ac04",
			2578 => x"fef82851",
			2579 => x"00002851",
			2580 => x"0901fe3c",
			2581 => x"07068518",
			2582 => x"0409db14",
			2583 => x"0b06a510",
			2584 => x"05076404",
			2585 => x"0000292d",
			2586 => x"0002ee04",
			2587 => x"0000292d",
			2588 => x"07061404",
			2589 => x"0000292d",
			2590 => x"011e292d",
			2591 => x"ffef292d",
			2592 => x"fe78292d",
			2593 => x"0d09851c",
			2594 => x"0601900c",
			2595 => x"0706ca08",
			2596 => x"06017404",
			2597 => x"0000292d",
			2598 => x"00a6292d",
			2599 => x"ff25292d",
			2600 => x"040cd808",
			2601 => x"05086a04",
			2602 => x"0000292d",
			2603 => x"0132292d",
			2604 => x"0b07c404",
			2605 => x"ffde292d",
			2606 => x"0000292d",
			2607 => x"0601b304",
			2608 => x"fee8292d",
			2609 => x"0000292d",
			2610 => x"030a2810",
			2611 => x"0003910c",
			2612 => x"0b06dd08",
			2613 => x"0b06be04",
			2614 => x"00aa292d",
			2615 => x"0000292d",
			2616 => x"01b5292d",
			2617 => x"0000292d",
			2618 => x"00038d04",
			2619 => x"ff2b292d",
			2620 => x"0003cf14",
			2621 => x"0902180c",
			2622 => x"0d087f04",
			2623 => x"0000292d",
			2624 => x"0706cb04",
			2625 => x"016b292d",
			2626 => x"0000292d",
			2627 => x"0c061a04",
			2628 => x"000e292d",
			2629 => x"ff43292d",
			2630 => x"030b6308",
			2631 => x"0003d904",
			2632 => x"0000292d",
			2633 => x"ff26292d",
			2634 => x"0000292d",
			2635 => x"0901fe3c",
			2636 => x"07068518",
			2637 => x"0409db14",
			2638 => x"0b06a510",
			2639 => x"05076404",
			2640 => x"00002a09",
			2641 => x"0002ee04",
			2642 => x"00002a09",
			2643 => x"07061404",
			2644 => x"00002a09",
			2645 => x"01452a09",
			2646 => x"ffcc2a09",
			2647 => x"fe712a09",
			2648 => x"0d09851c",
			2649 => x"0601900c",
			2650 => x"0706ca08",
			2651 => x"06017404",
			2652 => x"00002a09",
			2653 => x"00b22a09",
			2654 => x"ff0c2a09",
			2655 => x"040cd808",
			2656 => x"05086a04",
			2657 => x"00002a09",
			2658 => x"013f2a09",
			2659 => x"0b07c404",
			2660 => x"ffc32a09",
			2661 => x"00002a09",
			2662 => x"0601b304",
			2663 => x"fecc2a09",
			2664 => x"00002a09",
			2665 => x"040aa910",
			2666 => x"020a2d0c",
			2667 => x"0507e608",
			2668 => x"0507cc04",
			2669 => x"00b12a09",
			2670 => x"00002a09",
			2671 => x"01d32a09",
			2672 => x"00002a09",
			2673 => x"0b06ff04",
			2674 => x"ff142a09",
			2675 => x"0003d918",
			2676 => x"00038c08",
			2677 => x"040ab204",
			2678 => x"00002a09",
			2679 => x"ff3e2a09",
			2680 => x"0d090d08",
			2681 => x"0003cf04",
			2682 => x"01372a09",
			2683 => x"00002a09",
			2684 => x"0c065004",
			2685 => x"00002a09",
			2686 => x"ffba2a09",
			2687 => x"020ba004",
			2688 => x"ff332a09",
			2689 => x"00002a09",
			2690 => x"0100ff14",
			2691 => x"0003a210",
			2692 => x"0309ef0c",
			2693 => x"0c061004",
			2694 => x"fe6b2ab5",
			2695 => x"0e086804",
			2696 => x"03cd2ab5",
			2697 => x"fe7b2ab5",
			2698 => x"04982ab5",
			2699 => x"fe612ab5",
			2700 => x"09021f3c",
			2701 => x"05082e20",
			2702 => x"040abb1c",
			2703 => x"0901f60c",
			2704 => x"02092808",
			2705 => x"02092004",
			2706 => x"feb52ab5",
			2707 => x"022c2ab5",
			2708 => x"fe762ab5",
			2709 => x"0209dd08",
			2710 => x"06017904",
			2711 => x"042c2ab5",
			2712 => x"02012ab5",
			2713 => x"0b06ff04",
			2714 => x"fe2d2ab5",
			2715 => x"03f32ab5",
			2716 => x"fe462ab5",
			2717 => x"0802e008",
			2718 => x"0901a104",
			2719 => x"00cd2ab5",
			2720 => x"fe722ab5",
			2721 => x"020a9908",
			2722 => x"030a6904",
			2723 => x"06052ab5",
			2724 => x"01262ab5",
			2725 => x"0e0a5104",
			2726 => x"fe3d2ab5",
			2727 => x"0b07d604",
			2728 => x"01ab2ab5",
			2729 => x"ff702ab5",
			2730 => x"01015004",
			2731 => x"00702ab5",
			2732 => x"fe692ab5",
			2733 => x"0b068d04",
			2734 => x"fe6f2b21",
			2735 => x"0d09db30",
			2736 => x"0e0b5120",
			2737 => x"0003f21c",
			2738 => x"0a02390c",
			2739 => x"0b06ae08",
			2740 => x"07064004",
			2741 => x"00002b21",
			2742 => x"00f42b21",
			2743 => x"feac2b21",
			2744 => x"06017908",
			2745 => x"0209e804",
			2746 => x"01cd2b21",
			2747 => x"ff692b21",
			2748 => x"0c05fc04",
			2749 => x"fedf2b21",
			2750 => x"00572b21",
			2751 => x"feaf2b21",
			2752 => x"0803650c",
			2753 => x"040c0c04",
			2754 => x"00002b21",
			2755 => x"01015304",
			2756 => x"020b2b21",
			2757 => x"00002b21",
			2758 => x"00002b21",
			2759 => x"feaa2b21",
			2760 => x"0003782c",
			2761 => x"0e09c128",
			2762 => x"0a023918",
			2763 => x"0b069c10",
			2764 => x"0b067a04",
			2765 => x"00002bf5",
			2766 => x"0409a008",
			2767 => x"04090804",
			2768 => x"00002bf5",
			2769 => x"00972bf5",
			2770 => x"00002bf5",
			2771 => x"0b06ae04",
			2772 => x"00002bf5",
			2773 => x"ffb22bf5",
			2774 => x"0e08fd04",
			2775 => x"00002bf5",
			2776 => x"0d07ee04",
			2777 => x"00002bf5",
			2778 => x"040a8804",
			2779 => x"013c2bf5",
			2780 => x"00002bf5",
			2781 => x"ff752bf5",
			2782 => x"0e0a4810",
			2783 => x"09021d08",
			2784 => x"01015304",
			2785 => x"fea92bf5",
			2786 => x"00002bf5",
			2787 => x"01015804",
			2788 => x"002b2bf5",
			2789 => x"00002bf5",
			2790 => x"00039d08",
			2791 => x"020ad104",
			2792 => x"fee52bf5",
			2793 => x"00002bf5",
			2794 => x"020ac30c",
			2795 => x"0d087f04",
			2796 => x"00002bf5",
			2797 => x"0d08f404",
			2798 => x"01112bf5",
			2799 => x"00002bf5",
			2800 => x"0b07a410",
			2801 => x"0c066c08",
			2802 => x"0d090f04",
			2803 => x"ffca2bf5",
			2804 => x"00002bf5",
			2805 => x"06019004",
			2806 => x"00002bf5",
			2807 => x"00642bf5",
			2808 => x"0c068b04",
			2809 => x"00002bf5",
			2810 => x"0f0c0904",
			2811 => x"ff2a2bf5",
			2812 => x"00002bf5",
			2813 => x"0100ff14",
			2814 => x"00036310",
			2815 => x"0309ef0c",
			2816 => x"0100b008",
			2817 => x"0705a104",
			2818 => x"fe882c99",
			2819 => x"03d82c99",
			2820 => x"fe6c2c99",
			2821 => x"04452c99",
			2822 => x"fe632c99",
			2823 => x"0101583c",
			2824 => x"05082e1c",
			2825 => x"040abb18",
			2826 => x"0101360c",
			2827 => x"02092808",
			2828 => x"02092004",
			2829 => x"fec22c99",
			2830 => x"02022c99",
			2831 => x"fe7b2c99",
			2832 => x"030a1208",
			2833 => x"00039204",
			2834 => x"02a32c99",
			2835 => x"fef32c99",
			2836 => x"fe122c99",
			2837 => x"fe4a2c99",
			2838 => x"0802e008",
			2839 => x"01010604",
			2840 => x"006f2c99",
			2841 => x"fe712c99",
			2842 => x"0d09850c",
			2843 => x"020a7204",
			2844 => x"05022c99",
			2845 => x"0a026c04",
			2846 => x"fef22c99",
			2847 => x"018e2c99",
			2848 => x"0601af04",
			2849 => x"fbac2c99",
			2850 => x"08033f04",
			2851 => x"00cb2c99",
			2852 => x"02de2c99",
			2853 => x"fe6b2c99",
			2854 => x"0901961c",
			2855 => x"0003a218",
			2856 => x"0002e604",
			2857 => x"fe642d55",
			2858 => x"0002ee04",
			2859 => x"00482d55",
			2860 => x"00039e0c",
			2861 => x"00034b04",
			2862 => x"fe762d55",
			2863 => x"00035304",
			2864 => x"058a2d55",
			2865 => x"fe7e2d55",
			2866 => x"00002d55",
			2867 => x"fe602d55",
			2868 => x"0902193c",
			2869 => x"0d088d1c",
			2870 => x"09020a14",
			2871 => x"02093008",
			2872 => x"0a023304",
			2873 => x"fe7c2d55",
			2874 => x"175b2d55",
			2875 => x"040a8808",
			2876 => x"00037004",
			2877 => x"fe6a2d55",
			2878 => x"05c62d55",
			2879 => x"fe532d55",
			2880 => x"0a026704",
			2881 => x"04822d55",
			2882 => x"fe672d55",
			2883 => x"06018c0c",
			2884 => x"05083e04",
			2885 => x"03942d55",
			2886 => x"0003a604",
			2887 => x"fe642d55",
			2888 => x"fcb22d55",
			2889 => x"020ac304",
			2890 => x"0b1b2d55",
			2891 => x"0901f608",
			2892 => x"0d098504",
			2893 => x"02272d55",
			2894 => x"00392d55",
			2895 => x"040c2404",
			2896 => x"06472d55",
			2897 => x"01382d55",
			2898 => x"030a3904",
			2899 => x"04392d55",
			2900 => x"fe612d55",
			2901 => x"0c05d908",
			2902 => x"01014d04",
			2903 => x"fe982e11",
			2904 => x"00002e11",
			2905 => x"040ba43c",
			2906 => x"0802de20",
			2907 => x"0507900c",
			2908 => x"0409c708",
			2909 => x"02087c04",
			2910 => x"00002e11",
			2911 => x"010d2e11",
			2912 => x"00002e11",
			2913 => x"0d089a0c",
			2914 => x"09020808",
			2915 => x"0b06ae04",
			2916 => x"00002e11",
			2917 => x"fef02e11",
			2918 => x"00002e11",
			2919 => x"0b072f04",
			2920 => x"00482e11",
			2921 => x"00002e11",
			2922 => x"0d08da10",
			2923 => x"0b06dd04",
			2924 => x"fff82e11",
			2925 => x"08030808",
			2926 => x"0c05f404",
			2927 => x"00002e11",
			2928 => x"01552e11",
			2929 => x"00002e11",
			2930 => x"06019004",
			2931 => x"ff132e11",
			2932 => x"01014e04",
			2933 => x"00d22e11",
			2934 => x"00002e11",
			2935 => x"0e0ae104",
			2936 => x"fec62e11",
			2937 => x"05091b10",
			2938 => x"0d08f404",
			2939 => x"fff12e11",
			2940 => x"01014d08",
			2941 => x"01010b04",
			2942 => x"00002e11",
			2943 => x"012d2e11",
			2944 => x"00002e11",
			2945 => x"0601b304",
			2946 => x"feff2e11",
			2947 => x"00002e11",
			2948 => x"0c05bb04",
			2949 => x"feb72ea5",
			2950 => x"0c06c43c",
			2951 => x"07065a14",
			2952 => x"00038e10",
			2953 => x"0901e804",
			2954 => x"00002ea5",
			2955 => x"0c061608",
			2956 => x"040abb04",
			2957 => x"013a2ea5",
			2958 => x"00002ea5",
			2959 => x"00002ea5",
			2960 => x"ff942ea5",
			2961 => x"0e0aee18",
			2962 => x"040ba410",
			2963 => x"0003a308",
			2964 => x"0100e704",
			2965 => x"00002ea5",
			2966 => x"ff752ea5",
			2967 => x"0b072f04",
			2968 => x"fffa2ea5",
			2969 => x"00c82ea5",
			2970 => x"0e0ae104",
			2971 => x"fef02ea5",
			2972 => x"00002ea5",
			2973 => x"0b077304",
			2974 => x"00002ea5",
			2975 => x"09021908",
			2976 => x"0004c904",
			2977 => x"014d2ea5",
			2978 => x"00002ea5",
			2979 => x"00002ea5",
			2980 => x"07070f04",
			2981 => x"00002ea5",
			2982 => x"0601af04",
			2983 => x"fece2ea5",
			2984 => x"00002ea5",
			2985 => x"0100da04",
			2986 => x"fe672f21",
			2987 => x"09021f34",
			2988 => x"00033e04",
			2989 => x"fe812f21",
			2990 => x"040aa918",
			2991 => x"0507e70c",
			2992 => x"0409db04",
			2993 => x"02bb2f21",
			2994 => x"01014104",
			2995 => x"fe9a2f21",
			2996 => x"00162f21",
			2997 => x"0e09fd08",
			2998 => x"00034b04",
			2999 => x"00002f21",
			3000 => x"047c2f21",
			3001 => x"ff432f21",
			3002 => x"0e0b320c",
			3003 => x"040c1208",
			3004 => x"0b06ff04",
			3005 => x"fe7c2f21",
			3006 => x"00dd2f21",
			3007 => x"fdc82f21",
			3008 => x"08031804",
			3009 => x"ff442f21",
			3010 => x"0901fc04",
			3011 => x"01532f21",
			3012 => x"03122f21",
			3013 => x"040aa904",
			3014 => x"00b02f21",
			3015 => x"fe7a2f21",
			3016 => x"0c05bb04",
			3017 => x"fe862fed",
			3018 => x"0901f62c",
			3019 => x"0e0b0418",
			3020 => x"0901a910",
			3021 => x"040b5d0c",
			3022 => x"06014604",
			3023 => x"00002fed",
			3024 => x"0c05f404",
			3025 => x"00002fed",
			3026 => x"00bd2fed",
			3027 => x"ffb92fed",
			3028 => x"0e0abb04",
			3029 => x"feda2fed",
			3030 => x"00002fed",
			3031 => x"030c250c",
			3032 => x"030b1004",
			3033 => x"00002fed",
			3034 => x"0004a704",
			3035 => x"01092fed",
			3036 => x"00002fed",
			3037 => x"05092904",
			3038 => x"00002fed",
			3039 => x"ffc82fed",
			3040 => x"0c061714",
			3041 => x"09020808",
			3042 => x"06017b04",
			3043 => x"00b72fed",
			3044 => x"ff042fed",
			3045 => x"0003b308",
			3046 => x"0b06dd04",
			3047 => x"00002fed",
			3048 => x"01b02fed",
			3049 => x"ffe42fed",
			3050 => x"0802fc0c",
			3051 => x"09020e08",
			3052 => x"09020a04",
			3053 => x"ff1b2fed",
			3054 => x"009c2fed",
			3055 => x"fea12fed",
			3056 => x"0508a30c",
			3057 => x"08031208",
			3058 => x"09020e04",
			3059 => x"00a62fed",
			3060 => x"00002fed",
			3061 => x"ff412fed",
			3062 => x"0e0ad004",
			3063 => x"00002fed",
			3064 => x"09021f04",
			3065 => x"017b2fed",
			3066 => x"00002fed",
			3067 => x"05076404",
			3068 => x"fe713081",
			3069 => x"030a1220",
			3070 => x"0a023308",
			3071 => x"0100cd04",
			3072 => x"013a3081",
			3073 => x"fec23081",
			3074 => x"00038d14",
			3075 => x"0507ea0c",
			3076 => x"0409db04",
			3077 => x"01d83081",
			3078 => x"09020a04",
			3079 => x"feb73081",
			3080 => x"00f83081",
			3081 => x"040a3a04",
			3082 => x"00003081",
			3083 => x"01e23081",
			3084 => x"ff313081",
			3085 => x"00038c04",
			3086 => x"fe4a3081",
			3087 => x"0b070104",
			3088 => x"fe9c3081",
			3089 => x"0c066610",
			3090 => x"01014b08",
			3091 => x"05083004",
			3092 => x"feb03081",
			3093 => x"00b93081",
			3094 => x"08032804",
			3095 => x"01f33081",
			3096 => x"00003081",
			3097 => x"0a027b08",
			3098 => x"0706b704",
			3099 => x"00003081",
			3100 => x"fea43081",
			3101 => x"0d09db04",
			3102 => x"00703081",
			3103 => x"fe9f3081",
			3104 => x"01013448",
			3105 => x"0c05f708",
			3106 => x"030a8a04",
			3107 => x"fe75318d",
			3108 => x"0000318d",
			3109 => x"0003a21c",
			3110 => x"0601740c",
			3111 => x"02087e08",
			3112 => x"0d07fd04",
			3113 => x"0010318d",
			3114 => x"0000318d",
			3115 => x"ff04318d",
			3116 => x"0b06f004",
			3117 => x"0000318d",
			3118 => x"05086a08",
			3119 => x"01012e04",
			3120 => x"018e318d",
			3121 => x"0000318d",
			3122 => x"0000318d",
			3123 => x"0e0b0410",
			3124 => x"0901b80c",
			3125 => x"09019604",
			3126 => x"fefe318d",
			3127 => x"0901a904",
			3128 => x"0057318d",
			3129 => x"0000318d",
			3130 => x"fe8a318d",
			3131 => x"0b07f60c",
			3132 => x"030b1004",
			3133 => x"0000318d",
			3134 => x"0004bc04",
			3135 => x"0130318d",
			3136 => x"0000318d",
			3137 => x"0d09db04",
			3138 => x"0000318d",
			3139 => x"ff76318d",
			3140 => x"0c066634",
			3141 => x"0d086610",
			3142 => x"0309d80c",
			3143 => x"0901fe04",
			3144 => x"ffd2318d",
			3145 => x"00037d04",
			3146 => x"0158318d",
			3147 => x"0000318d",
			3148 => x"febe318d",
			3149 => x"05080f08",
			3150 => x"09020804",
			3151 => x"0000318d",
			3152 => x"02ca318d",
			3153 => x"0003a60c",
			3154 => x"030a3908",
			3155 => x"0a025304",
			3156 => x"0000318d",
			3157 => x"0144318d",
			3158 => x"fe8e318d",
			3159 => x"08032808",
			3160 => x"05083004",
			3161 => x"0000318d",
			3162 => x"01d2318d",
			3163 => x"020ba004",
			3164 => x"fff1318d",
			3165 => x"0000318d",
			3166 => x"01013f04",
			3167 => x"00b1318d",
			3168 => x"0e0bab04",
			3169 => x"fec3318d",
			3170 => x"0000318d",
			3171 => x"0c05bb04",
			3172 => x"fe743249",
			3173 => x"09020e48",
			3174 => x"0b069c14",
			3175 => x"00034b10",
			3176 => x"06014604",
			3177 => x"00003249",
			3178 => x"0409db08",
			3179 => x"07060204",
			3180 => x"00003249",
			3181 => x"01c23249",
			3182 => x"00003249",
			3183 => x"ffda3249",
			3184 => x"0b06ed18",
			3185 => x"0b06ae0c",
			3186 => x"0409db08",
			3187 => x"0901db04",
			3188 => x"00003249",
			3189 => x"006c3249",
			3190 => x"00003249",
			3191 => x"0507ea04",
			3192 => x"feaf3249",
			3193 => x"0507f404",
			3194 => x"00003249",
			3195 => x"ff563249",
			3196 => x"0003b70c",
			3197 => x"06017404",
			3198 => x"ff413249",
			3199 => x"01012e04",
			3200 => x"018b3249",
			3201 => x"00493249",
			3202 => x"0e0abb08",
			3203 => x"0003c004",
			3204 => x"00003249",
			3205 => x"fe593249",
			3206 => x"0d09db04",
			3207 => x"00f33249",
			3208 => x"feca3249",
			3209 => x"0c061610",
			3210 => x"0c061208",
			3211 => x"0b06d204",
			3212 => x"00003249",
			3213 => x"ff493249",
			3214 => x"0003cf04",
			3215 => x"015e3249",
			3216 => x"00003249",
			3217 => x"fe613249",
			3218 => x"0c05d708",
			3219 => x"01014904",
			3220 => x"fe6c32f5",
			3221 => x"000032f5",
			3222 => x"0d09db4c",
			3223 => x"0e0b293c",
			3224 => x"020ad120",
			3225 => x"0003a310",
			3226 => x"0e0a2a08",
			3227 => x"040a6904",
			3228 => x"000232f5",
			3229 => x"016c32f5",
			3230 => x"01013c04",
			3231 => x"003d32f5",
			3232 => x"fde632f5",
			3233 => x"09020208",
			3234 => x"0706a104",
			3235 => x"fea132f5",
			3236 => x"00c832f5",
			3237 => x"0c065204",
			3238 => x"021332f5",
			3239 => x"ffe332f5",
			3240 => x"0e0abb10",
			3241 => x"020aec08",
			3242 => x"01012104",
			3243 => x"005e32f5",
			3244 => x"ff4532f5",
			3245 => x"0a027a04",
			3246 => x"000032f5",
			3247 => x"fe3132f5",
			3248 => x"08030204",
			3249 => x"feb832f5",
			3250 => x"08032604",
			3251 => x"010632f5",
			3252 => x"fedf32f5",
			3253 => x"0101490c",
			3254 => x"0004a708",
			3255 => x"05089404",
			3256 => x"000032f5",
			3257 => x"01af32f5",
			3258 => x"000032f5",
			3259 => x"ff6d32f5",
			3260 => x"fe6332f5",
			3261 => x"0e08fd04",
			3262 => x"fe683393",
			3263 => x"0d09db48",
			3264 => x"0e0b3234",
			3265 => x"0706cc1c",
			3266 => x"08030f0c",
			3267 => x"06016b04",
			3268 => x"fea43393",
			3269 => x"06017b04",
			3270 => x"02d53393",
			3271 => x"01363393",
			3272 => x"0d08f408",
			3273 => x"0b074404",
			3274 => x"fe293393",
			3275 => x"ff7a3393",
			3276 => x"040be404",
			3277 => x"02023393",
			3278 => x"00003393",
			3279 => x"0e0b040c",
			3280 => x"040bca08",
			3281 => x"0802fc04",
			3282 => x"fe8b3393",
			3283 => x"00cb3393",
			3284 => x"fded3393",
			3285 => x"0003c804",
			3286 => x"ff173393",
			3287 => x"0003f704",
			3288 => x"01713393",
			3289 => x"00003393",
			3290 => x"08036510",
			3291 => x"05089404",
			3292 => x"ffba3393",
			3293 => x"0706ca04",
			3294 => x"058c3393",
			3295 => x"08030f04",
			3296 => x"fff23393",
			3297 => x"01c43393",
			3298 => x"ff463393",
			3299 => x"fe493393",
			3300 => x"00003395",
			3301 => x"00003399",
			3302 => x"0000339d",
			3303 => x"000033a1",
			3304 => x"000033a5",
			3305 => x"000033a9",
			3306 => x"000033ad",
			3307 => x"000033b1",
			3308 => x"000033b5",
			3309 => x"000033b9",
			3310 => x"000033bd",
			3311 => x"000033c1",
			3312 => x"000033c5",
			3313 => x"000033c9",
			3314 => x"000033cd",
			3315 => x"000033d1",
			3316 => x"000033d5",
			3317 => x"000033d9",
			3318 => x"000033dd",
			3319 => x"09020804",
			3320 => x"fffc33e9",
			3321 => x"000033e9",
			3322 => x"06018604",
			3323 => x"000033fd",
			3324 => x"0601bc04",
			3325 => x"001333fd",
			3326 => x"000033fd",
			3327 => x"01014108",
			3328 => x"01012504",
			3329 => x"00003411",
			3330 => x"00513411",
			3331 => x"00003411",
			3332 => x"01014f08",
			3333 => x"0002f604",
			3334 => x"00003425",
			3335 => x"ffe63425",
			3336 => x"00003425",
			3337 => x"09020808",
			3338 => x"0601af04",
			3339 => x"ffcc3439",
			3340 => x"00003439",
			3341 => x"00003439",
			3342 => x"07068608",
			3343 => x"07065b04",
			3344 => x"00003455",
			3345 => x"ffea3455",
			3346 => x"07070c04",
			3347 => x"00363455",
			3348 => x"00003455",
			3349 => x"00038e0c",
			3350 => x"0802aa04",
			3351 => x"00003471",
			3352 => x"0802eb04",
			3353 => x"001e3471",
			3354 => x"00003471",
			3355 => x"fff63471",
			3356 => x"040b0404",
			3357 => x"0000348d",
			3358 => x"020cab08",
			3359 => x"01011d04",
			3360 => x"0000348d",
			3361 => x"ffcc348d",
			3362 => x"0000348d",
			3363 => x"0901f604",
			3364 => x"000034a9",
			3365 => x"05094208",
			3366 => x"09022a04",
			3367 => x"004d34a9",
			3368 => x"000034a9",
			3369 => x"000034a9",
			3370 => x"00038e0c",
			3371 => x"09020804",
			3372 => x"000034d5",
			3373 => x"0f0a5a04",
			3374 => x"006134d5",
			3375 => x"000034d5",
			3376 => x"030af108",
			3377 => x"00039604",
			3378 => x"000034d5",
			3379 => x"ffbe34d5",
			3380 => x"000034d5",
			3381 => x"0b06dd04",
			3382 => x"000034f9",
			3383 => x"0601bc0c",
			3384 => x"06018504",
			3385 => x"000034f9",
			3386 => x"0b07b804",
			3387 => x"003534f9",
			3388 => x"000034f9",
			3389 => x"000034f9",
			3390 => x"0901fc04",
			3391 => x"0000351d",
			3392 => x"0b07a10c",
			3393 => x"09022c08",
			3394 => x"0901fe04",
			3395 => x"0000351d",
			3396 => x"002c351d",
			3397 => x"0000351d",
			3398 => x"0000351d",
			3399 => x"0003b710",
			3400 => x"0a023904",
			3401 => x"00003549",
			3402 => x"05089708",
			3403 => x"0507ea04",
			3404 => x"00003549",
			3405 => x"00443549",
			3406 => x"00003549",
			3407 => x"020cab04",
			3408 => x"fff53549",
			3409 => x"00003549",
			3410 => x"0901dd04",
			3411 => x"00003575",
			3412 => x"01014108",
			3413 => x"0802aa04",
			3414 => x"00003575",
			3415 => x"00363575",
			3416 => x"030a0104",
			3417 => x"00003575",
			3418 => x"030b6304",
			3419 => x"ffdb3575",
			3420 => x"00003575",
			3421 => x"09020a14",
			3422 => x"0706a108",
			3423 => x"0409db04",
			3424 => x"000035b1",
			3425 => x"ff6c35b1",
			3426 => x"07070f08",
			3427 => x"0b073304",
			3428 => x"000035b1",
			3429 => x"002035b1",
			3430 => x"000035b1",
			3431 => x"07068808",
			3432 => x"09022d04",
			3433 => x"003335b1",
			3434 => x"000035b1",
			3435 => x"000035b1",
			3436 => x"0003d914",
			3437 => x"0a023304",
			3438 => x"000035dd",
			3439 => x"09020e0c",
			3440 => x"09015504",
			3441 => x"000035dd",
			3442 => x"00033e04",
			3443 => x"000035dd",
			3444 => x"001135dd",
			3445 => x"000035dd",
			3446 => x"fff235dd",
			3447 => x"0802ed0c",
			3448 => x"09020804",
			3449 => x"00003621",
			3450 => x"020a3a04",
			3451 => x"00783621",
			3452 => x"00003621",
			3453 => x"0e0ac10c",
			3454 => x"01015108",
			3455 => x"040a9504",
			3456 => x"00003621",
			3457 => x"ff9f3621",
			3458 => x"00003621",
			3459 => x"0d09db08",
			3460 => x"0706a104",
			3461 => x"00003621",
			3462 => x"00473621",
			3463 => x"00003621",
			3464 => x"0802ed10",
			3465 => x"0507ea04",
			3466 => x"00003665",
			3467 => x"00035b04",
			3468 => x"00003665",
			3469 => x"05083e04",
			3470 => x"005c3665",
			3471 => x"00003665",
			3472 => x"0e0ac110",
			3473 => x"0101510c",
			3474 => x"040af504",
			3475 => x"00003665",
			3476 => x"0901b804",
			3477 => x"00003665",
			3478 => x"ff853665",
			3479 => x"00003665",
			3480 => x"00003665",
			3481 => x"0901dd10",
			3482 => x"0706a10c",
			3483 => x"0e0a4808",
			3484 => x"06014704",
			3485 => x"000036b9",
			3486 => x"ffd136b9",
			3487 => x"000036b9",
			3488 => x"000036b9",
			3489 => x"0101410c",
			3490 => x"0a023304",
			3491 => x"000036b9",
			3492 => x"0e08e104",
			3493 => x"000036b9",
			3494 => x"004b36b9",
			3495 => x"030a0104",
			3496 => x"000036b9",
			3497 => x"030b6308",
			3498 => x"0c061404",
			3499 => x"000036b9",
			3500 => x"ffbb36b9",
			3501 => x"000036b9",
			3502 => x"040aa918",
			3503 => x"0e09fd14",
			3504 => x"0d078804",
			3505 => x"000036f5",
			3506 => x"08025f04",
			3507 => x"000036f5",
			3508 => x"0d08b308",
			3509 => x"00039104",
			3510 => x"005836f5",
			3511 => x"000036f5",
			3512 => x"000036f5",
			3513 => x"000036f5",
			3514 => x"0e0a8604",
			3515 => x"ffce36f5",
			3516 => x"000036f5",
			3517 => x"0b072018",
			3518 => x"0802f314",
			3519 => x"0b06dd04",
			3520 => x"00003741",
			3521 => x"0f09e104",
			3522 => x"00003741",
			3523 => x"0c05f404",
			3524 => x"00003741",
			3525 => x"040a4904",
			3526 => x"00003741",
			3527 => x"008c3741",
			3528 => x"00003741",
			3529 => x"0802fc08",
			3530 => x"0e095104",
			3531 => x"00003741",
			3532 => x"ffca3741",
			3533 => x"08033704",
			3534 => x"00153741",
			3535 => x"00003741",
			3536 => x"05083004",
			3537 => x"00003775",
			3538 => x"0d09c414",
			3539 => x"09021510",
			3540 => x"00038c04",
			3541 => x"00003775",
			3542 => x"0e0a1b04",
			3543 => x"00003775",
			3544 => x"08036504",
			3545 => x"00723775",
			3546 => x"00003775",
			3547 => x"00003775",
			3548 => x"00003775",
			3549 => x"0901fc04",
			3550 => x"000037a9",
			3551 => x"0706ce14",
			3552 => x"040c1810",
			3553 => x"0901fe04",
			3554 => x"000037a9",
			3555 => x"09022d08",
			3556 => x"0508b504",
			3557 => x"004437a9",
			3558 => x"000037a9",
			3559 => x"000037a9",
			3560 => x"000037a9",
			3561 => x"000037a9",
			3562 => x"040abb18",
			3563 => x"030a2814",
			3564 => x"0802a504",
			3565 => x"000037f5",
			3566 => x"0802eb0c",
			3567 => x"0b06dc04",
			3568 => x"000037f5",
			3569 => x"0309a304",
			3570 => x"000037f5",
			3571 => x"005737f5",
			3572 => x"000037f5",
			3573 => x"000037f5",
			3574 => x"030ae104",
			3575 => x"ffeb37f5",
			3576 => x"0b083508",
			3577 => x"0b073304",
			3578 => x"000037f5",
			3579 => x"001037f5",
			3580 => x"000037f5",
			3581 => x"0802c314",
			3582 => x"0a023304",
			3583 => x"00003859",
			3584 => x"0a02450c",
			3585 => x"06017c08",
			3586 => x"06016804",
			3587 => x"00003859",
			3588 => x"00223859",
			3589 => x"00003859",
			3590 => x"00003859",
			3591 => x"06018e08",
			3592 => x"01014b04",
			3593 => x"ff333859",
			3594 => x"00003859",
			3595 => x"0003d90c",
			3596 => x"020a9304",
			3597 => x"00003859",
			3598 => x"0802f104",
			3599 => x"00003859",
			3600 => x"00653859",
			3601 => x"00041808",
			3602 => x"0a02b904",
			3603 => x"ffa13859",
			3604 => x"00003859",
			3605 => x"00003859",
			3606 => x"0601850c",
			3607 => x"040a0104",
			3608 => x"000038a5",
			3609 => x"09021b04",
			3610 => x"ff7938a5",
			3611 => x"000038a5",
			3612 => x"0c06c418",
			3613 => x"00038c04",
			3614 => x"000038a5",
			3615 => x"00040b10",
			3616 => x"0b06ff04",
			3617 => x"000038a5",
			3618 => x"09021f08",
			3619 => x"0d086604",
			3620 => x"000038a5",
			3621 => x"008438a5",
			3622 => x"000038a5",
			3623 => x"000038a5",
			3624 => x"000038a5",
			3625 => x"0c061108",
			3626 => x"0f0a9e04",
			3627 => x"ff5c38e9",
			3628 => x"000038e9",
			3629 => x"0d09db18",
			3630 => x"0b06ff04",
			3631 => x"000038e9",
			3632 => x"040aa904",
			3633 => x"000038e9",
			3634 => x"07070c0c",
			3635 => x"040c1808",
			3636 => x"0d088204",
			3637 => x"000038e9",
			3638 => x"006c38e9",
			3639 => x"000038e9",
			3640 => x"000038e9",
			3641 => x"ffe738e9",
			3642 => x"09020814",
			3643 => x"0c061708",
			3644 => x"00037804",
			3645 => x"00003945",
			3646 => x"ffb73945",
			3647 => x"0c06fe08",
			3648 => x"040d1b04",
			3649 => x"00153945",
			3650 => x"00003945",
			3651 => x"00003945",
			3652 => x"0c066618",
			3653 => x"09022d14",
			3654 => x"00038504",
			3655 => x"00003945",
			3656 => x"0c05f604",
			3657 => x"00003945",
			3658 => x"08032808",
			3659 => x"0802de04",
			3660 => x"00003945",
			3661 => x"009a3945",
			3662 => x"00003945",
			3663 => x"00003945",
			3664 => x"00003945",
			3665 => x"0e09c118",
			3666 => x"00037d14",
			3667 => x"06014604",
			3668 => x"000039b1",
			3669 => x"05084d0c",
			3670 => x"0c05bb04",
			3671 => x"000039b1",
			3672 => x"08025f04",
			3673 => x"000039b1",
			3674 => x"009e39b1",
			3675 => x"000039b1",
			3676 => x"000039b1",
			3677 => x"0c06500c",
			3678 => x"020aa608",
			3679 => x"01014b04",
			3680 => x"ff4539b1",
			3681 => x"000039b1",
			3682 => x"000039b1",
			3683 => x"0d09db10",
			3684 => x"0e0b3204",
			3685 => x"000039b1",
			3686 => x"09021908",
			3687 => x"0004c904",
			3688 => x"006f39b1",
			3689 => x"000039b1",
			3690 => x"000039b1",
			3691 => x"000039b1",
			3692 => x"0c061108",
			3693 => x"0e0a5104",
			3694 => x"ff3f3a0d",
			3695 => x"00003a0d",
			3696 => x"07070c18",
			3697 => x"0b06ff04",
			3698 => x"00003a0d",
			3699 => x"040c2410",
			3700 => x"040aa904",
			3701 => x"00003a0d",
			3702 => x"0d088204",
			3703 => x"00003a0d",
			3704 => x"0d093704",
			3705 => x"00923a0d",
			3706 => x"00003a0d",
			3707 => x"00003a0d",
			3708 => x"040cf50c",
			3709 => x"0c068b04",
			3710 => x"00003a0d",
			3711 => x"0b07a404",
			3712 => x"00003a0d",
			3713 => x"ffad3a0d",
			3714 => x"00003a0d",
			3715 => x"0901dd14",
			3716 => x"0e0a390c",
			3717 => x"04091d04",
			3718 => x"00003a89",
			3719 => x"0c068704",
			3720 => x"ff323a89",
			3721 => x"00003a89",
			3722 => x"05090a04",
			3723 => x"00143a89",
			3724 => x"00003a89",
			3725 => x"0e09fd10",
			3726 => x"0507e404",
			3727 => x"00003a89",
			3728 => x"00036304",
			3729 => x"00003a89",
			3730 => x"00039104",
			3731 => x"00b93a89",
			3732 => x"00003a89",
			3733 => x"0003a308",
			3734 => x"0802e604",
			3735 => x"00003a89",
			3736 => x"ff9c3a89",
			3737 => x"05094f10",
			3738 => x"06019404",
			3739 => x"00003a89",
			3740 => x"05083004",
			3741 => x"00003a89",
			3742 => x"0601be04",
			3743 => x"00953a89",
			3744 => x"00003a89",
			3745 => x"00003a89",
			3746 => x"0c061414",
			3747 => x"0901e808",
			3748 => x"0e0a8404",
			3749 => x"ff1b3afd",
			3750 => x"00003afd",
			3751 => x"0507f508",
			3752 => x"05079e04",
			3753 => x"00003afd",
			3754 => x"fff63afd",
			3755 => x"000a3afd",
			3756 => x"05094f24",
			3757 => x"030b6318",
			3758 => x"0f0aed10",
			3759 => x"06019d0c",
			3760 => x"00035b04",
			3761 => x"00003afd",
			3762 => x"09021f04",
			3763 => x"00be3afd",
			3764 => x"00003afd",
			3765 => x"00003afd",
			3766 => x"030ac504",
			3767 => x"ff9e3afd",
			3768 => x"00003afd",
			3769 => x"09021908",
			3770 => x"00048204",
			3771 => x"00d93afd",
			3772 => x"00003afd",
			3773 => x"00003afd",
			3774 => x"ff813afd",
			3775 => x"0e09c118",
			3776 => x"00037d14",
			3777 => x"06014604",
			3778 => x"00003b79",
			3779 => x"0b07330c",
			3780 => x"0c05bb04",
			3781 => x"00003b79",
			3782 => x"08025f04",
			3783 => x"00003b79",
			3784 => x"00a93b79",
			3785 => x"00003b79",
			3786 => x"00003b79",
			3787 => x"0c065010",
			3788 => x"040b560c",
			3789 => x"07064004",
			3790 => x"00003b79",
			3791 => x"06019d04",
			3792 => x"ff583b79",
			3793 => x"00003b79",
			3794 => x"00003b79",
			3795 => x"0d09db14",
			3796 => x"0e0b3208",
			3797 => x"040bca04",
			3798 => x"00003b79",
			3799 => x"ffff3b79",
			3800 => x"09021908",
			3801 => x"0004c904",
			3802 => x"00793b79",
			3803 => x"00003b79",
			3804 => x"00003b79",
			3805 => x"00003b79",
			3806 => x"0901dd18",
			3807 => x"0c061708",
			3808 => x"0e0a5104",
			3809 => x"ff173c05",
			3810 => x"00003c05",
			3811 => x"0508fb08",
			3812 => x"0d089a04",
			3813 => x"00003c05",
			3814 => x"00053c05",
			3815 => x"0d096904",
			3816 => x"00003c05",
			3817 => x"ffea3c05",
			3818 => x"0c05f810",
			3819 => x"0802eb0c",
			3820 => x"0901e804",
			3821 => x"00003c05",
			3822 => x"0e08e104",
			3823 => x"00003c05",
			3824 => x"00e73c05",
			3825 => x"00003c05",
			3826 => x"06018e08",
			3827 => x"0209c904",
			3828 => x"00003c05",
			3829 => x"ff6c3c05",
			3830 => x"0b080514",
			3831 => x"0b071e08",
			3832 => x"0f0a5a04",
			3833 => x"00003c05",
			3834 => x"fff53c05",
			3835 => x"0003a304",
			3836 => x"00003c05",
			3837 => x"08036504",
			3838 => x"00e83c05",
			3839 => x"00003c05",
			3840 => x"ffde3c05",
			3841 => x"040af51c",
			3842 => x"0d08b318",
			3843 => x"06019214",
			3844 => x"00038e10",
			3845 => x"06014604",
			3846 => x"00003c79",
			3847 => x"020a4608",
			3848 => x"07060204",
			3849 => x"00003c79",
			3850 => x"00813c79",
			3851 => x"00003c79",
			3852 => x"00003c79",
			3853 => x"00003c79",
			3854 => x"00003c79",
			3855 => x"0e0aee08",
			3856 => x"01011504",
			3857 => x"00003c79",
			3858 => x"ff4f3c79",
			3859 => x"0d09db14",
			3860 => x"0706a104",
			3861 => x"00003c79",
			3862 => x"01010604",
			3863 => x"00003c79",
			3864 => x"01015008",
			3865 => x"0e0afd04",
			3866 => x"00003c79",
			3867 => x"00c23c79",
			3868 => x"00003c79",
			3869 => x"00003c79",
			3870 => x"0e08fd10",
			3871 => x"07064304",
			3872 => x"fe6d3ced",
			3873 => x"07064408",
			3874 => x"0d07fd04",
			3875 => x"00f73ced",
			3876 => x"00003ced",
			3877 => x"ff0f3ced",
			3878 => x"0d09db28",
			3879 => x"0e0b5118",
			3880 => x"0003f214",
			3881 => x"0a023304",
			3882 => x"fed13ced",
			3883 => x"0209e808",
			3884 => x"01013704",
			3885 => x"02443ced",
			3886 => x"00743ced",
			3887 => x"0003a304",
			3888 => x"ff2f3ced",
			3889 => x"00b83ced",
			3890 => x"fe9e3ced",
			3891 => x"0803650c",
			3892 => x"0706cb04",
			3893 => x"04203ced",
			3894 => x"01015104",
			3895 => x"01ab3ced",
			3896 => x"00003ced",
			3897 => x"00003ced",
			3898 => x"fe933ced",
			3899 => x"0003d92c",
			3900 => x"06016804",
			3901 => x"00003d51",
			3902 => x"030a2814",
			3903 => x"0507ea04",
			3904 => x"00003d51",
			3905 => x"06017404",
			3906 => x"00003d51",
			3907 => x"00039108",
			3908 => x"00034b04",
			3909 => x"00003d51",
			3910 => x"00c93d51",
			3911 => x"00003d51",
			3912 => x"0f0a9204",
			3913 => x"ffce3d51",
			3914 => x"06018e04",
			3915 => x"00003d51",
			3916 => x"030a8a04",
			3917 => x"00003d51",
			3918 => x"0a026c04",
			3919 => x"00003d51",
			3920 => x"00633d51",
			3921 => x"020cab04",
			3922 => x"ffe33d51",
			3923 => x"00003d51",
			3924 => x"0901f428",
			3925 => x"0c061008",
			3926 => x"0409c704",
			3927 => x"00003de5",
			3928 => x"ff293de5",
			3929 => x"020a8310",
			3930 => x"06014604",
			3931 => x"00003de5",
			3932 => x"040b0408",
			3933 => x"08025f04",
			3934 => x"00003de5",
			3935 => x"00223de5",
			3936 => x"00003de5",
			3937 => x"0e0abb04",
			3938 => x"ff7d3de5",
			3939 => x"030c2508",
			3940 => x"0e0ae104",
			3941 => x"00003de5",
			3942 => x"00403de5",
			3943 => x"00003de5",
			3944 => x"0c06e320",
			3945 => x"0b06dd08",
			3946 => x"040a5b04",
			3947 => x"00003de5",
			3948 => x"ffbf3de5",
			3949 => x"00037004",
			3950 => x"00003de5",
			3951 => x"01015810",
			3952 => x"0e0a6d08",
			3953 => x"0d08da04",
			3954 => x"011d3de5",
			3955 => x"00003de5",
			3956 => x"0e0b5104",
			3957 => x"ffdb3de5",
			3958 => x"00d33de5",
			3959 => x"00003de5",
			3960 => x"ffbe3de5",
			3961 => x"0901f42c",
			3962 => x"07068508",
			3963 => x"0409c704",
			3964 => x"00003e99",
			3965 => x"fec33e99",
			3966 => x"0b07a414",
			3967 => x"040ba410",
			3968 => x"0f09b104",
			3969 => x"00003e99",
			3970 => x"0a023904",
			3971 => x"00003e99",
			3972 => x"0508b304",
			3973 => x"00a83e99",
			3974 => x"00003e99",
			3975 => x"00003e99",
			3976 => x"030b930c",
			3977 => x"0c068b04",
			3978 => x"00003e99",
			3979 => x"0c06c504",
			3980 => x"ff8d3e99",
			3981 => x"00003e99",
			3982 => x"00003e99",
			3983 => x"0c06301c",
			3984 => x"0003af18",
			3985 => x"0507e408",
			3986 => x"0c05db04",
			3987 => x"00343e99",
			3988 => x"00003e99",
			3989 => x"0c05f604",
			3990 => x"00003e99",
			3991 => x"01013c04",
			3992 => x"00003e99",
			3993 => x"0901fe04",
			3994 => x"00003e99",
			3995 => x"013a3e99",
			3996 => x"00003e99",
			3997 => x"0101450c",
			3998 => x"0e0a5a04",
			3999 => x"00003e99",
			4000 => x"05086a04",
			4001 => x"00003e99",
			4002 => x"00843e99",
			4003 => x"0b072004",
			4004 => x"00003e99",
			4005 => x"ff323e99",
			4006 => x"0706400c",
			4007 => x"01013d04",
			4008 => x"fe653f15",
			4009 => x"0d080b04",
			4010 => x"026b3f15",
			4011 => x"feda3f15",
			4012 => x"0d09db30",
			4013 => x"01015428",
			4014 => x"05082110",
			4015 => x"0d07b004",
			4016 => x"034a3f15",
			4017 => x"01013804",
			4018 => x"fe673f15",
			4019 => x"0e09fd04",
			4020 => x"01373f15",
			4021 => x"fe903f15",
			4022 => x"040cd80c",
			4023 => x"0100e704",
			4024 => x"068c3f15",
			4025 => x"06018604",
			4026 => x"fe8a3f15",
			4027 => x"017c3f15",
			4028 => x"0e0c0604",
			4029 => x"fdb33f15",
			4030 => x"07074e04",
			4031 => x"00ed3f15",
			4032 => x"04c13f15",
			4033 => x"0c061504",
			4034 => x"02003f15",
			4035 => x"fe713f15",
			4036 => x"fe323f15",
			4037 => x"0706400c",
			4038 => x"01013d04",
			4039 => x"fe663f99",
			4040 => x"0d080b04",
			4041 => x"01ef3f99",
			4042 => x"ff003f99",
			4043 => x"0d09db34",
			4044 => x"0e0b5120",
			4045 => x"0003ed18",
			4046 => x"01015410",
			4047 => x"06018e08",
			4048 => x"0100dc04",
			4049 => x"027a3f99",
			4050 => x"ffd73f99",
			4051 => x"0d087204",
			4052 => x"feaf3f99",
			4053 => x"01cb3f99",
			4054 => x"0d088d04",
			4055 => x"01a73f99",
			4056 => x"fe783f99",
			4057 => x"0e0b3204",
			4058 => x"fdfe3f99",
			4059 => x"00003f99",
			4060 => x"0706b704",
			4061 => x"079d3f99",
			4062 => x"0803650c",
			4063 => x"01015108",
			4064 => x"040cce04",
			4065 => x"01a93f99",
			4066 => x"02dd3f99",
			4067 => x"ffb63f99",
			4068 => x"ff1e3f99",
			4069 => x"fe3f3f99",
			4070 => x"00038e24",
			4071 => x"09020818",
			4072 => x"06017914",
			4073 => x"0d084b10",
			4074 => x"06014604",
			4075 => x"0000403d",
			4076 => x"07065a08",
			4077 => x"07061404",
			4078 => x"0000403d",
			4079 => x"0098403d",
			4080 => x"0000403d",
			4081 => x"0000403d",
			4082 => x"ff9d403d",
			4083 => x"07068508",
			4084 => x"030a3904",
			4085 => x"013d403d",
			4086 => x"0000403d",
			4087 => x"0000403d",
			4088 => x"0e0a3904",
			4089 => x"fef1403d",
			4090 => x"0e0b3218",
			4091 => x"040be414",
			4092 => x"09020a0c",
			4093 => x"07070d08",
			4094 => x"05084d04",
			4095 => x"0000403d",
			4096 => x"00e8403d",
			4097 => x"0000403d",
			4098 => x"0e0a5a04",
			4099 => x"0000403d",
			4100 => x"ff8d403d",
			4101 => x"ff4e403d",
			4102 => x"0b080510",
			4103 => x"0b077104",
			4104 => x"0000403d",
			4105 => x"09021908",
			4106 => x"0004bc04",
			4107 => x"012a403d",
			4108 => x"0000403d",
			4109 => x"0000403d",
			4110 => x"ffcf403d",
			4111 => x"0c05d908",
			4112 => x"09021504",
			4113 => x"fe6b40b9",
			4114 => x"000040b9",
			4115 => x"0d09db34",
			4116 => x"0e0b2924",
			4117 => x"040be41c",
			4118 => x"0e0a6d10",
			4119 => x"09020808",
			4120 => x"06017b04",
			4121 => x"00d540b9",
			4122 => x"ff1d40b9",
			4123 => x"0c061704",
			4124 => x"022040b9",
			4125 => x"fffe40b9",
			4126 => x"09021508",
			4127 => x"07069b04",
			4128 => x"ff5540b9",
			4129 => x"011040b9",
			4130 => x"fdfa40b9",
			4131 => x"0e0aee04",
			4132 => x"fe3140b9",
			4133 => x"000040b9",
			4134 => x"0101490c",
			4135 => x"0004a708",
			4136 => x"030b1b04",
			4137 => x"000040b9",
			4138 => x"01b440b9",
			4139 => x"000040b9",
			4140 => x"ff5940b9",
			4141 => x"fe5840b9",
			4142 => x"040a8828",
			4143 => x"0e09c124",
			4144 => x"06016810",
			4145 => x"04091d0c",
			4146 => x"04090804",
			4147 => x"0000417d",
			4148 => x"09016f04",
			4149 => x"001b417d",
			4150 => x"0000417d",
			4151 => x"ffd4417d",
			4152 => x"0a025710",
			4153 => x"0a023304",
			4154 => x"0000417d",
			4155 => x"0e08e104",
			4156 => x"0000417d",
			4157 => x"05078e04",
			4158 => x"0000417d",
			4159 => x"0137417d",
			4160 => x"0000417d",
			4161 => x"ff9e417d",
			4162 => x"0e0a4810",
			4163 => x"09021d08",
			4164 => x"01015304",
			4165 => x"fea2417d",
			4166 => x"0000417d",
			4167 => x"01015804",
			4168 => x"0033417d",
			4169 => x"0000417d",
			4170 => x"0e0a6310",
			4171 => x"0601960c",
			4172 => x"020a8604",
			4173 => x"0000417d",
			4174 => x"06018904",
			4175 => x"0000417d",
			4176 => x"00d1417d",
			4177 => x"0000417d",
			4178 => x"01014918",
			4179 => x"0c06a90c",
			4180 => x"06018e04",
			4181 => x"0000417d",
			4182 => x"0c063204",
			4183 => x"0000417d",
			4184 => x"00aa417d",
			4185 => x"0601af08",
			4186 => x"0901bf04",
			4187 => x"0000417d",
			4188 => x"ff18417d",
			4189 => x"0000417d",
			4190 => x"feb4417d",
			4191 => x"0b080540",
			4192 => x"0e0b3230",
			4193 => x"0003dd28",
			4194 => x"0f0a6e10",
			4195 => x"0d08b30c",
			4196 => x"0901f604",
			4197 => x"00004201",
			4198 => x"09020e04",
			4199 => x"00d44201",
			4200 => x"00004201",
			4201 => x"00004201",
			4202 => x"0b072f08",
			4203 => x"07068304",
			4204 => x"ff164201",
			4205 => x"00004201",
			4206 => x"0003a308",
			4207 => x"030a8104",
			4208 => x"00004201",
			4209 => x"ffdd4201",
			4210 => x"0e0a6304",
			4211 => x"00004201",
			4212 => x"00bf4201",
			4213 => x"0003ea04",
			4214 => x"00004201",
			4215 => x"ff224201",
			4216 => x"0c064d04",
			4217 => x"00004201",
			4218 => x"09021908",
			4219 => x"0004c904",
			4220 => x"010b4201",
			4221 => x"00004201",
			4222 => x"00004201",
			4223 => x"ff5c4201",
			4224 => x"040a8828",
			4225 => x"0e09c124",
			4226 => x"0802d520",
			4227 => x"0a023914",
			4228 => x"0b069c0c",
			4229 => x"0b067a04",
			4230 => x"000042cd",
			4231 => x"0409a004",
			4232 => x"008c42cd",
			4233 => x"000042cd",
			4234 => x"0b06ae04",
			4235 => x"000042cd",
			4236 => x"ffc042cd",
			4237 => x"0d07ee04",
			4238 => x"000042cd",
			4239 => x"0e08fd04",
			4240 => x"000042cd",
			4241 => x"012a42cd",
			4242 => x"000042cd",
			4243 => x"ffc642cd",
			4244 => x"0e0a4814",
			4245 => x"09021d0c",
			4246 => x"040aa904",
			4247 => x"000042cd",
			4248 => x"01015304",
			4249 => x"fe9a42cd",
			4250 => x"000042cd",
			4251 => x"01015804",
			4252 => x"003642cd",
			4253 => x"000042cd",
			4254 => x"01014920",
			4255 => x"0b07a410",
			4256 => x"0d089a04",
			4257 => x"000042cd",
			4258 => x"040c2408",
			4259 => x"040b0204",
			4260 => x"000042cd",
			4261 => x"011342cd",
			4262 => x"000042cd",
			4263 => x"0e0b0e04",
			4264 => x"ff2942cd",
			4265 => x"0d09b608",
			4266 => x"0b07f604",
			4267 => x"009042cd",
			4268 => x"000042cd",
			4269 => x"ff5842cd",
			4270 => x"0e0a5a08",
			4271 => x"0c063404",
			4272 => x"005842cd",
			4273 => x"000042cd",
			4274 => x"fed042cd",
			4275 => x"020b1644",
			4276 => x"020ac32c",
			4277 => x"0e08e10c",
			4278 => x"0c061004",
			4279 => x"bf8f43a9",
			4280 => x"0c061104",
			4281 => x"c18c43a9",
			4282 => x"bfa543a9",
			4283 => x"0d08f41c",
			4284 => x"01014910",
			4285 => x"0706a108",
			4286 => x"0901fe04",
			4287 => x"bfbb43a9",
			4288 => x"c2f543a9",
			4289 => x"00037804",
			4290 => x"c4f443a9",
			4291 => x"e6ad43a9",
			4292 => x"020a2004",
			4293 => x"f80043a9",
			4294 => x"01014e04",
			4295 => x"cafe43a9",
			4296 => x"c15d43a9",
			4297 => x"bf9243a9",
			4298 => x"0901d408",
			4299 => x"0003f204",
			4300 => x"0aa943a9",
			4301 => x"c02343a9",
			4302 => x"0902120c",
			4303 => x"05084d04",
			4304 => x"bf9d43a9",
			4305 => x"0706b704",
			4306 => x"ed4043a9",
			4307 => x"c55a43a9",
			4308 => x"bf9443a9",
			4309 => x"08035a24",
			4310 => x"0901ee08",
			4311 => x"030ae504",
			4312 => x"bfe443a9",
			4313 => x"0ffb43a9",
			4314 => x"0e0bab14",
			4315 => x"09020a08",
			4316 => x"05086a04",
			4317 => x"bfab43a9",
			4318 => x"ec3443a9",
			4319 => x"09021908",
			4320 => x"020b4904",
			4321 => x"c00343a9",
			4322 => x"c5cf43a9",
			4323 => x"bf9643a9",
			4324 => x"01015b04",
			4325 => x"f62e43a9",
			4326 => x"c00343a9",
			4327 => x"08036504",
			4328 => x"c55a43a9",
			4329 => x"bf9143a9",
			4330 => x"0901d92c",
			4331 => x"0c061708",
			4332 => x"0f0ad704",
			4333 => x"fe98448d",
			4334 => x"0000448d",
			4335 => x"0d09751c",
			4336 => x"0100fc0c",
			4337 => x"0100e008",
			4338 => x"0f0abc04",
			4339 => x"002c448d",
			4340 => x"0000448d",
			4341 => x"ff80448d",
			4342 => x"00038c04",
			4343 => x"0000448d",
			4344 => x"040c7f08",
			4345 => x"0a02a604",
			4346 => x"0107448d",
			4347 => x"0000448d",
			4348 => x"0000448d",
			4349 => x"0e0b2904",
			4350 => x"ff2d448d",
			4351 => x"0000448d",
			4352 => x"040aa91c",
			4353 => x"0b06fc14",
			4354 => x"0901e804",
			4355 => x"0000448d",
			4356 => x"00038e0c",
			4357 => x"0d07ee04",
			4358 => x"0000448d",
			4359 => x"0a023904",
			4360 => x"0000448d",
			4361 => x"015c448d",
			4362 => x"0000448d",
			4363 => x"030a0104",
			4364 => x"0000448d",
			4365 => x"ff91448d",
			4366 => x"0706860c",
			4367 => x"01015304",
			4368 => x"feca448d",
			4369 => x"0003c804",
			4370 => x"007f448d",
			4371 => x"0000448d",
			4372 => x"0706ce10",
			4373 => x"0803280c",
			4374 => x"0003a304",
			4375 => x"0000448d",
			4376 => x"09021d04",
			4377 => x"0169448d",
			4378 => x"0000448d",
			4379 => x"0000448d",
			4380 => x"0101450c",
			4381 => x"0a028e04",
			4382 => x"0000448d",
			4383 => x"0c06c504",
			4384 => x"0076448d",
			4385 => x"0000448d",
			4386 => x"ff56448d",
			4387 => x"0c05bb04",
			4388 => x"fec54531",
			4389 => x"0706ce38",
			4390 => x"09020a24",
			4391 => x"06017914",
			4392 => x"0901e808",
			4393 => x"0100e704",
			4394 => x"00004531",
			4395 => x"ffdd4531",
			4396 => x"0c05f808",
			4397 => x"0d07ee04",
			4398 => x"00004531",
			4399 => x"012a4531",
			4400 => x"00004531",
			4401 => x"07069b04",
			4402 => x"fea64531",
			4403 => x"040be908",
			4404 => x"0c067104",
			4405 => x"01064531",
			4406 => x"00004531",
			4407 => x"00004531",
			4408 => x"06019208",
			4409 => x"07068504",
			4410 => x"01054531",
			4411 => x"00004531",
			4412 => x"0b071e04",
			4413 => x"ff414531",
			4414 => x"09021904",
			4415 => x"00f54531",
			4416 => x"00004531",
			4417 => x"0e0ae108",
			4418 => x"0100fa04",
			4419 => x"00004531",
			4420 => x"fef24531",
			4421 => x"07074e0c",
			4422 => x"01014708",
			4423 => x"0004d204",
			4424 => x"00ea4531",
			4425 => x"00004531",
			4426 => x"00004531",
			4427 => x"ff214531",
			4428 => x"0802eb2c",
			4429 => x"0d08b328",
			4430 => x"06014604",
			4431 => x"000045ed",
			4432 => x"0b06dd18",
			4433 => x"03094f0c",
			4434 => x"0802bb08",
			4435 => x"0b06ae04",
			4436 => x"00ce45ed",
			4437 => x"000045ed",
			4438 => x"000045ed",
			4439 => x"0c05c204",
			4440 => x"000045ed",
			4441 => x"0507f604",
			4442 => x"ffe445ed",
			4443 => x"000045ed",
			4444 => x"0802b704",
			4445 => x"000045ed",
			4446 => x"07065804",
			4447 => x"000045ed",
			4448 => x"014e45ed",
			4449 => x"ffae45ed",
			4450 => x"0d08b308",
			4451 => x"0b072f04",
			4452 => x"fedd45ed",
			4453 => x"000045ed",
			4454 => x"07070c10",
			4455 => x"040c240c",
			4456 => x"06019004",
			4457 => x"000045ed",
			4458 => x"09021904",
			4459 => x"011f45ed",
			4460 => x"000045ed",
			4461 => x"000045ed",
			4462 => x"0601af10",
			4463 => x"07070f04",
			4464 => x"000045ed",
			4465 => x"0b07a404",
			4466 => x"000045ed",
			4467 => x"0c068b04",
			4468 => x"000045ed",
			4469 => x"ff2b45ed",
			4470 => x"01014708",
			4471 => x"040d2e04",
			4472 => x"00db45ed",
			4473 => x"000045ed",
			4474 => x"000045ed",
			4475 => x"0100fc18",
			4476 => x"0003a214",
			4477 => x"0e09770c",
			4478 => x"0c061004",
			4479 => x"fe6746b1",
			4480 => x"0507ba04",
			4481 => x"08b646b1",
			4482 => x"fe7346b1",
			4483 => x"0b072f04",
			4484 => x"0c2946b1",
			4485 => x"000046b1",
			4486 => x"fe5e46b1",
			4487 => x"09021f44",
			4488 => x"05082e20",
			4489 => x"040a9518",
			4490 => x"0901fe0c",
			4491 => x"0901e804",
			4492 => x"fe6e46b1",
			4493 => x"0409db04",
			4494 => x"0cdc46b1",
			4495 => x"ff7a46b1",
			4496 => x"0e09a204",
			4497 => x"07fe46b1",
			4498 => x"0a025404",
			4499 => x"fdd246b1",
			4500 => x"016c46b1",
			4501 => x"01015104",
			4502 => x"fe4a46b1",
			4503 => x"007c46b1",
			4504 => x"0802e510",
			4505 => x"0901a108",
			4506 => x"0b072f04",
			4507 => x"ffbb46b1",
			4508 => x"014246b1",
			4509 => x"07072404",
			4510 => x"fe6d46b1",
			4511 => x"fcaf46b1",
			4512 => x"05094210",
			4513 => x"0c061708",
			4514 => x"0e0a6d04",
			4515 => x"0d5e46b1",
			4516 => x"010646b1",
			4517 => x"06018c04",
			4518 => x"ff2746b1",
			4519 => x"01e546b1",
			4520 => x"fe1146b1",
			4521 => x"040aa904",
			4522 => x"016546b1",
			4523 => x"fe6546b1",
			4524 => x"0100fc14",
			4525 => x"0003a210",
			4526 => x"0309ef0c",
			4527 => x"0c061004",
			4528 => x"fe66476d",
			4529 => x"0b06bb04",
			4530 => x"0f73476d",
			4531 => x"fe71476d",
			4532 => x"07af476d",
			4533 => x"fe5e476d",
			4534 => x"09021d44",
			4535 => x"05084d28",
			4536 => x"0901fe18",
			4537 => x"02094d08",
			4538 => x"0a023904",
			4539 => x"fe77476d",
			4540 => x"0d2e476d",
			4541 => x"0d086d08",
			4542 => x"0507f504",
			4543 => x"fe68476d",
			4544 => x"ff2b476d",
			4545 => x"05081304",
			4546 => x"fd48476d",
			4547 => x"fe90476d",
			4548 => x"0209dd04",
			4549 => x"08e0476d",
			4550 => x"01014b04",
			4551 => x"fe45476d",
			4552 => x"0a027404",
			4553 => x"03ca476d",
			4554 => x"fed3476d",
			4555 => x"0a026c0c",
			4556 => x"0706b404",
			4557 => x"021b476d",
			4558 => x"07072504",
			4559 => x"fe65476d",
			4560 => x"fc75476d",
			4561 => x"0509420c",
			4562 => x"020ab504",
			4563 => x"0653476d",
			4564 => x"0a027504",
			4565 => x"fcd1476d",
			4566 => x"0203476d",
			4567 => x"fdca476d",
			4568 => x"030a5c04",
			4569 => x"0354476d",
			4570 => x"fe64476d",
			4571 => x"00038e38",
			4572 => x"0901e810",
			4573 => x"06017404",
			4574 => x"ff6f4841",
			4575 => x"0a024108",
			4576 => x"00034b04",
			4577 => x"00004841",
			4578 => x"00144841",
			4579 => x"00004841",
			4580 => x"030a2820",
			4581 => x"0b06dd18",
			4582 => x"0a02450c",
			4583 => x"07064608",
			4584 => x"0e08fd04",
			4585 => x"00004841",
			4586 => x"00c74841",
			4587 => x"00004841",
			4588 => x"0f09a304",
			4589 => x"00004841",
			4590 => x"0b06bd04",
			4591 => x"00004841",
			4592 => x"ffb94841",
			4593 => x"00037004",
			4594 => x"00004841",
			4595 => x"01934841",
			4596 => x"00038d04",
			4597 => x"ffdf4841",
			4598 => x"00004841",
			4599 => x"0e0a3904",
			4600 => x"fea14841",
			4601 => x"07073c28",
			4602 => x"0d08b314",
			4603 => x"0601990c",
			4604 => x"0c061204",
			4605 => x"00004841",
			4606 => x"0d086604",
			4607 => x"00004841",
			4608 => x"00694841",
			4609 => x"07066e04",
			4610 => x"00004841",
			4611 => x"ff0c4841",
			4612 => x"06019004",
			4613 => x"00004841",
			4614 => x"0003f308",
			4615 => x"09021904",
			4616 => x"01334841",
			4617 => x"00004841",
			4618 => x"0e0b5104",
			4619 => x"ffd84841",
			4620 => x"00004841",
			4621 => x"0d099c04",
			4622 => x"00004841",
			4623 => x"ff6f4841",
			4624 => x"0b067a04",
			4625 => x"fe6a48b5",
			4626 => x"05096134",
			4627 => x"0e0b3224",
			4628 => x"040c0c20",
			4629 => x"0706cc10",
			4630 => x"07068508",
			4631 => x"0c061a04",
			4632 => x"009348b5",
			4633 => x"fe1448b5",
			4634 => x"0a029304",
			4635 => x"01a348b5",
			4636 => x"ff4348b5",
			4637 => x"08030208",
			4638 => x"0a027b04",
			4639 => x"fe9f48b5",
			4640 => x"000048b5",
			4641 => x"01014b04",
			4642 => x"016d48b5",
			4643 => x"ffb748b5",
			4644 => x"fdf948b5",
			4645 => x"0101490c",
			4646 => x"0004a008",
			4647 => x"030b4604",
			4648 => x"000048b5",
			4649 => x"01c148b5",
			4650 => x"ff7448b5",
			4651 => x"ff2748b5",
			4652 => x"fe3248b5",
			4653 => x"0901d934",
			4654 => x"0c061708",
			4655 => x"0f0ad704",
			4656 => x"fe8e49b1",
			4657 => x"000049b1",
			4658 => x"0508fb24",
			4659 => x"0100ff14",
			4660 => x"0c06300c",
			4661 => x"05083e08",
			4662 => x"08026904",
			4663 => x"000049b1",
			4664 => x"008349b1",
			4665 => x"000049b1",
			4666 => x"05089404",
			4667 => x"ff5649b1",
			4668 => x"000049b1",
			4669 => x"00038c04",
			4670 => x"000049b1",
			4671 => x"040c7f08",
			4672 => x"08033404",
			4673 => x"010b49b1",
			4674 => x"000049b1",
			4675 => x"000049b1",
			4676 => x"01011b04",
			4677 => x"ff0e49b1",
			4678 => x"000049b1",
			4679 => x"040aa920",
			4680 => x"0b06fc18",
			4681 => x"0901e804",
			4682 => x"000049b1",
			4683 => x"00038e10",
			4684 => x"0507e408",
			4685 => x"03096804",
			4686 => x"00d949b1",
			4687 => x"000049b1",
			4688 => x"0a024104",
			4689 => x"000049b1",
			4690 => x"01bc49b1",
			4691 => x"000049b1",
			4692 => x"030a0104",
			4693 => x"000049b1",
			4694 => x"ff6d49b1",
			4695 => x"0706860c",
			4696 => x"01015304",
			4697 => x"feb949b1",
			4698 => x"0003c804",
			4699 => x"009c49b1",
			4700 => x"000049b1",
			4701 => x"0706ce10",
			4702 => x"0803280c",
			4703 => x"0003a304",
			4704 => x"000049b1",
			4705 => x"09021d04",
			4706 => x"018149b1",
			4707 => x"000049b1",
			4708 => x"000049b1",
			4709 => x"0101450c",
			4710 => x"0601a604",
			4711 => x"000049b1",
			4712 => x"0c06c504",
			4713 => x"009b49b1",
			4714 => x"000049b1",
			4715 => x"ff4549b1",
			4716 => x"0c05bd04",
			4717 => x"fe9f4a6d",
			4718 => x"040b9d3c",
			4719 => x"0a026920",
			4720 => x"030a1214",
			4721 => x"09020810",
			4722 => x"0100e708",
			4723 => x"06014204",
			4724 => x"00004a6d",
			4725 => x"00854a6d",
			4726 => x"0b06ae04",
			4727 => x"00004a6d",
			4728 => x"ff0e4a6d",
			4729 => x"00f34a6d",
			4730 => x"0c061404",
			4731 => x"00004a6d",
			4732 => x"0802eb04",
			4733 => x"ff6d4a6d",
			4734 => x"00004a6d",
			4735 => x"0d090d14",
			4736 => x"07066d08",
			4737 => x"0a026c04",
			4738 => x"00004a6d",
			4739 => x"ffd04a6d",
			4740 => x"0a029008",
			4741 => x"0d087204",
			4742 => x"00004a6d",
			4743 => x"015f4a6d",
			4744 => x"00004a6d",
			4745 => x"08030604",
			4746 => x"ffe44a6d",
			4747 => x"00004a6d",
			4748 => x"0e0aee08",
			4749 => x"040ba404",
			4750 => x"00004a6d",
			4751 => x"fee64a6d",
			4752 => x"05091b10",
			4753 => x"09020e0c",
			4754 => x"05088604",
			4755 => x"00004a6d",
			4756 => x"01010b04",
			4757 => x"00004a6d",
			4758 => x"011e4a6d",
			4759 => x"00004a6d",
			4760 => x"0601b304",
			4761 => x"ff0d4a6d",
			4762 => x"00004a6d",
			4763 => x"0100fc04",
			4764 => x"fe684b09",
			4765 => x"01014e44",
			4766 => x"05083020",
			4767 => x"0901fe0c",
			4768 => x"02094d08",
			4769 => x"0901e804",
			4770 => x"fe964b09",
			4771 => x"04ca4b09",
			4772 => x"fe634b09",
			4773 => x"040a5b04",
			4774 => x"03834b09",
			4775 => x"0d087208",
			4776 => x"01014b04",
			4777 => x"fe484b09",
			4778 => x"00004b09",
			4779 => x"0b06fc04",
			4780 => x"0c6e4b09",
			4781 => x"ff334b09",
			4782 => x"06018d0c",
			4783 => x"0d08b308",
			4784 => x"06016b04",
			4785 => x"ff884b09",
			4786 => x"03114b09",
			4787 => x"fdb24b09",
			4788 => x"040bf10c",
			4789 => x"01013d04",
			4790 => x"01d04b09",
			4791 => x"040b1c04",
			4792 => x"00fa4b09",
			4793 => x"03cb4b09",
			4794 => x"0e0b1604",
			4795 => x"fd994b09",
			4796 => x"0c06de04",
			4797 => x"01bd4b09",
			4798 => x"fff24b09",
			4799 => x"030a3904",
			4800 => x"027b4b09",
			4801 => x"fe694b09",
			4802 => x"09019604",
			4803 => x"fe694bb5",
			4804 => x"09021f4c",
			4805 => x"05083028",
			4806 => x"09020814",
			4807 => x"02094d08",
			4808 => x"0901e804",
			4809 => x"fe9d4bb5",
			4810 => x"03484bb5",
			4811 => x"0c061a04",
			4812 => x"fe694bb5",
			4813 => x"07065804",
			4814 => x"05e94bb5",
			4815 => x"fe7a4bb5",
			4816 => x"05080f0c",
			4817 => x"0d086508",
			4818 => x"040a9504",
			4819 => x"03264bb5",
			4820 => x"fee24bb5",
			4821 => x"08fd4bb5",
			4822 => x"0b071004",
			4823 => x"fe364bb5",
			4824 => x"00004bb5",
			4825 => x"06018d0c",
			4826 => x"0d08b308",
			4827 => x"030a0104",
			4828 => x"ff884bb5",
			4829 => x"02ed4bb5",
			4830 => x"fe234bb5",
			4831 => x"0003dd0c",
			4832 => x"09021908",
			4833 => x"0901fc04",
			4834 => x"01b64bb5",
			4835 => x"02bd4bb5",
			4836 => x"fed24bb5",
			4837 => x"0e0afd04",
			4838 => x"fdcb4bb5",
			4839 => x"0a029304",
			4840 => x"ffbd4bb5",
			4841 => x"01b24bb5",
			4842 => x"0c05de04",
			4843 => x"00304bb5",
			4844 => x"fe6d4bb5",
			4845 => x"0100fc04",
			4846 => x"fe6a4c59",
			4847 => x"01014e48",
			4848 => x"05083028",
			4849 => x"0901f60c",
			4850 => x"02092808",
			4851 => x"0f093d04",
			4852 => x"fee24c59",
			4853 => x"012a4c59",
			4854 => x"fe6a4c59",
			4855 => x"040a5b0c",
			4856 => x"06017c04",
			4857 => x"03e04c59",
			4858 => x"07065804",
			4859 => x"fefa4c59",
			4860 => x"02044c59",
			4861 => x"0d087208",
			4862 => x"01014b04",
			4863 => x"fe584c59",
			4864 => x"00004c59",
			4865 => x"05080f04",
			4866 => x"0acf4c59",
			4867 => x"ff0c4c59",
			4868 => x"06018504",
			4869 => x"fe5a4c59",
			4870 => x"040be410",
			4871 => x"00038c08",
			4872 => x"040ac204",
			4873 => x"03424c59",
			4874 => x"fe884c59",
			4875 => x"0706df04",
			4876 => x"02834c59",
			4877 => x"014f4c59",
			4878 => x"030b3204",
			4879 => x"fe1a4c59",
			4880 => x"0d098504",
			4881 => x"01aa4c59",
			4882 => x"fff54c59",
			4883 => x"030a3904",
			4884 => x"01e44c59",
			4885 => x"fe6c4c59",
			4886 => x"07060204",
			4887 => x"fe734d0d",
			4888 => x"0e09c11c",
			4889 => x"0a023308",
			4890 => x"0100cd04",
			4891 => x"010d4d0d",
			4892 => x"fecf4d0d",
			4893 => x"00037d10",
			4894 => x"0e08e104",
			4895 => x"00004d0d",
			4896 => x"040a8808",
			4897 => x"00033e04",
			4898 => x"00004d0d",
			4899 => x"01a04d0d",
			4900 => x"00004d0d",
			4901 => x"ff1b4d0d",
			4902 => x"00038504",
			4903 => x"fe644d0d",
			4904 => x"0c06661c",
			4905 => x"01014b0c",
			4906 => x"05083004",
			4907 => x"fe7a4d0d",
			4908 => x"0e0a8404",
			4909 => x"ffdf4d0d",
			4910 => x"011f4d0d",
			4911 => x"0b06ff08",
			4912 => x"0b06ef04",
			4913 => x"00c14d0d",
			4914 => x"ff8c4d0d",
			4915 => x"09021f04",
			4916 => x"01e04d0d",
			4917 => x"00004d0d",
			4918 => x"0e0afd0c",
			4919 => x"040bca08",
			4920 => x"0802fc04",
			4921 => x"ff084d0d",
			4922 => x"00634d0d",
			4923 => x"fe834d0d",
			4924 => x"0b080508",
			4925 => x"01014704",
			4926 => x"016e4d0d",
			4927 => x"ff474d0d",
			4928 => x"0d09db04",
			4929 => x"00004d0d",
			4930 => x"feaf4d0d",
			4931 => x"07061404",
			4932 => x"fe804e03",
			4933 => x"0101342c",
			4934 => x"0706a114",
			4935 => x"0f087a0c",
			4936 => x"0f087204",
			4937 => x"00004e03",
			4938 => x"08023004",
			4939 => x"00004e03",
			4940 => x"00ef4e03",
			4941 => x"07069b04",
			4942 => x"fe814e03",
			4943 => x"00004e03",
			4944 => x"0d096910",
			4945 => x"01012e0c",
			4946 => x"06018504",
			4947 => x"00004e03",
			4948 => x"00042904",
			4949 => x"014d4e03",
			4950 => x"00004e03",
			4951 => x"ffb84e03",
			4952 => x"01011b04",
			4953 => x"fea54e03",
			4954 => x"00004e03",
			4955 => x"01014120",
			4956 => x"0d087210",
			4957 => x"06017b0c",
			4958 => x"01013908",
			4959 => x"01013604",
			4960 => x"00004e03",
			4961 => x"011a4e03",
			4962 => x"00004e03",
			4963 => x"ff224e03",
			4964 => x"06018e04",
			4965 => x"00004e03",
			4966 => x"01013a04",
			4967 => x"00004e03",
			4968 => x"07066e04",
			4969 => x"00004e03",
			4970 => x"02074e03",
			4971 => x"01014f1c",
			4972 => x"030a120c",
			4973 => x"0b06de08",
			4974 => x"0b06be04",
			4975 => x"00004e03",
			4976 => x"ffe44e03",
			4977 => x"01274e03",
			4978 => x"0003a308",
			4979 => x"0b070e04",
			4980 => x"00004e03",
			4981 => x"fea14e03",
			4982 => x"0802f404",
			4983 => x"00fa4e03",
			4984 => x"ffaf4e03",
			4985 => x"0706b40c",
			4986 => x"0b06dd04",
			4987 => x"00004e03",
			4988 => x"08032804",
			4989 => x"018f4e03",
			4990 => x"00004e03",
			4991 => x"ff814e03",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1652, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(3300, initial_addr_3'length));
	end generate gen_rom_10;

	gen_rom_11: if SELECT_ROM = 11 generate
		bank <= (
			0 => x"00000005",
			1 => x"00000009",
			2 => x"0000000d",
			3 => x"00000011",
			4 => x"00000015",
			5 => x"00000019",
			6 => x"0000001d",
			7 => x"00000021",
			8 => x"00000025",
			9 => x"00000029",
			10 => x"0000002d",
			11 => x"00000031",
			12 => x"00000035",
			13 => x"00000039",
			14 => x"0000003d",
			15 => x"00000041",
			16 => x"00000045",
			17 => x"00000049",
			18 => x"0000004d",
			19 => x"00000051",
			20 => x"00000055",
			21 => x"00000059",
			22 => x"0000005d",
			23 => x"00000061",
			24 => x"00000065",
			25 => x"00000069",
			26 => x"0000006d",
			27 => x"00000071",
			28 => x"01013704",
			29 => x"ffff007d",
			30 => x"0000007d",
			31 => x"0802be04",
			32 => x"00000089",
			33 => x"fffb0089",
			34 => x"0209be08",
			35 => x"0e08e104",
			36 => x"0000009d",
			37 => x"ffdf009d",
			38 => x"0000009d",
			39 => x"0901d908",
			40 => x"00034b04",
			41 => x"000000b1",
			42 => x"ffa000b1",
			43 => x"000000b1",
			44 => x"01012408",
			45 => x"0901d904",
			46 => x"ffea00c5",
			47 => x"000000c5",
			48 => x"000000c5",
			49 => x"0901f008",
			50 => x"01013804",
			51 => x"fff800d9",
			52 => x"000000d9",
			53 => x"000000d9",
			54 => x"0802e60c",
			55 => x"01011104",
			56 => x"000000f5",
			57 => x"01014904",
			58 => x"003500f5",
			59 => x"000000f5",
			60 => x"000000f5",
			61 => x"01013f0c",
			62 => x"0e08e104",
			63 => x"00000111",
			64 => x"040b9d04",
			65 => x"ffc90111",
			66 => x"00000111",
			67 => x"00000111",
			68 => x"0901bc08",
			69 => x"04091d04",
			70 => x"0000013d",
			71 => x"ff98013d",
			72 => x"0e093308",
			73 => x"0409db04",
			74 => x"0000013d",
			75 => x"003c013d",
			76 => x"040a6904",
			77 => x"ff80013d",
			78 => x"0000013d",
			79 => x"0e08e10c",
			80 => x"09019c04",
			81 => x"00000169",
			82 => x"00030204",
			83 => x"00000169",
			84 => x"002e0169",
			85 => x"0901d908",
			86 => x"0d078804",
			87 => x"00000169",
			88 => x"ffa80169",
			89 => x"00000169",
			90 => x"01011704",
			91 => x"0000018d",
			92 => x"0902080c",
			93 => x"0802fb08",
			94 => x"0802aa04",
			95 => x"0000018d",
			96 => x"002a018d",
			97 => x"0000018d",
			98 => x"0000018d",
			99 => x"0e08e104",
			100 => x"000001b1",
			101 => x"0101370c",
			102 => x"0c060f08",
			103 => x"0c059f04",
			104 => x"000001b1",
			105 => x"ffbc01b1",
			106 => x"000001b1",
			107 => x"000001b1",
			108 => x"0901d908",
			109 => x"0b06ae04",
			110 => x"000001dd",
			111 => x"ffa001dd",
			112 => x"0c05da04",
			113 => x"000001dd",
			114 => x"0d082208",
			115 => x"0a026204",
			116 => x"007f01dd",
			117 => x"000001dd",
			118 => x"000001dd",
			119 => x"0901d90c",
			120 => x"02099508",
			121 => x"0802a504",
			122 => x"00000211",
			123 => x"ff9d0211",
			124 => x"00000211",
			125 => x"06017c08",
			126 => x"0c061004",
			127 => x"006b0211",
			128 => x"00000211",
			129 => x"020a1004",
			130 => x"fffb0211",
			131 => x"00000211",
			132 => x"01011708",
			133 => x"00031a04",
			134 => x"00000245",
			135 => x"fff10245",
			136 => x"0d086d10",
			137 => x"040a3a04",
			138 => x"00000245",
			139 => x"0e09c108",
			140 => x"00034b04",
			141 => x"00000245",
			142 => x"007c0245",
			143 => x"00000245",
			144 => x"00000245",
			145 => x"02097010",
			146 => x"0c06140c",
			147 => x"0e08cb04",
			148 => x"00000289",
			149 => x"06017404",
			150 => x"ffaf0289",
			151 => x"00000289",
			152 => x"00000289",
			153 => x"0f09950c",
			154 => x"040a0104",
			155 => x"00000289",
			156 => x"0a026d04",
			157 => x"00720289",
			158 => x"00000289",
			159 => x"040a8804",
			160 => x"ffc90289",
			161 => x"00000289",
			162 => x"01013f18",
			163 => x"0e08e110",
			164 => x"0e07dc04",
			165 => x"000002bd",
			166 => x"06015204",
			167 => x"000002bd",
			168 => x"0f09b104",
			169 => x"003902bd",
			170 => x"000002bd",
			171 => x"040b9d04",
			172 => x"ff9202bd",
			173 => x"000002bd",
			174 => x"000002bd",
			175 => x"0c05d818",
			176 => x"0d07e40c",
			177 => x"01010b04",
			178 => x"ff790319",
			179 => x"0802f804",
			180 => x"00500319",
			181 => x"00000319",
			182 => x"040a2808",
			183 => x"05079c04",
			184 => x"00000319",
			185 => x"feed0319",
			186 => x"00000319",
			187 => x"0d083810",
			188 => x"0901bc04",
			189 => x"00000319",
			190 => x"040a3a04",
			191 => x"00000319",
			192 => x"0e09c104",
			193 => x"00d00319",
			194 => x"00000319",
			195 => x"0e096204",
			196 => x"00000319",
			197 => x"ffe40319",
			198 => x"0101170c",
			199 => x"0901c308",
			200 => x"04091d04",
			201 => x"0000035d",
			202 => x"ffe5035d",
			203 => x"0000035d",
			204 => x"0d086d14",
			205 => x"040a3a04",
			206 => x"0000035d",
			207 => x"0e09c10c",
			208 => x"06018908",
			209 => x"00034b04",
			210 => x"0000035d",
			211 => x"0093035d",
			212 => x"0000035d",
			213 => x"0000035d",
			214 => x"0000035d",
			215 => x"0209be18",
			216 => x"0a024c14",
			217 => x"03096810",
			218 => x"0409db08",
			219 => x"0308f704",
			220 => x"000003b1",
			221 => x"ffc403b1",
			222 => x"0f08d404",
			223 => x"000003b1",
			224 => x"007a03b1",
			225 => x"000003b1",
			226 => x"fee603b1",
			227 => x"0309c00c",
			228 => x"06018808",
			229 => x"01010604",
			230 => x"000003b1",
			231 => x"00f603b1",
			232 => x"000003b1",
			233 => x"01013904",
			234 => x"ffae03b1",
			235 => x"000003b1",
			236 => x"02093004",
			237 => x"000003e5",
			238 => x"020a6b14",
			239 => x"01010604",
			240 => x"000003e5",
			241 => x"0101490c",
			242 => x"06015c04",
			243 => x"000003e5",
			244 => x"06018d04",
			245 => x"002d03e5",
			246 => x"000003e5",
			247 => x"000003e5",
			248 => x"000003e5",
			249 => x"0c05b80c",
			250 => x"01012108",
			251 => x"08029104",
			252 => x"00000441",
			253 => x"ff950441",
			254 => x"00000441",
			255 => x"0e08fd0c",
			256 => x"0a020004",
			257 => x"00000441",
			258 => x"09019c04",
			259 => x"00000441",
			260 => x"00a40441",
			261 => x"040a5b0c",
			262 => x"0901f208",
			263 => x"01012804",
			264 => x"00000441",
			265 => x"ff850441",
			266 => x"00000441",
			267 => x"0309d808",
			268 => x"01011f04",
			269 => x"00000441",
			270 => x"00730441",
			271 => x"00000441",
			272 => x"0c05d710",
			273 => x"0802be04",
			274 => x"000004a5",
			275 => x"0901ea08",
			276 => x"07062c04",
			277 => x"fe4904a5",
			278 => x"000004a5",
			279 => x"000004a5",
			280 => x"0c05fa10",
			281 => x"00035304",
			282 => x"000004a5",
			283 => x"0802e808",
			284 => x"0e09c104",
			285 => x"00dd04a5",
			286 => x"000004a5",
			287 => x"000004a5",
			288 => x"0e091508",
			289 => x"01011704",
			290 => x"000004a5",
			291 => x"001304a5",
			292 => x"040abb08",
			293 => x"0802ae04",
			294 => x"000004a5",
			295 => x"fef804a5",
			296 => x"000004a5",
			297 => x"0c05b810",
			298 => x"0101210c",
			299 => x"00033e04",
			300 => x"00000509",
			301 => x"07061504",
			302 => x"ff740509",
			303 => x"00000509",
			304 => x"00000509",
			305 => x"07062a0c",
			306 => x"0901f608",
			307 => x"01010604",
			308 => x"00000509",
			309 => x"00c00509",
			310 => x"00000509",
			311 => x"0e09240c",
			312 => x"02093004",
			313 => x"00000509",
			314 => x"01011304",
			315 => x"00000509",
			316 => x"00570509",
			317 => x"01013408",
			318 => x"0c061404",
			319 => x"ff500509",
			320 => x"00000509",
			321 => x"00000509",
			322 => x"0209700c",
			323 => x"0802a504",
			324 => x"00000565",
			325 => x"06017404",
			326 => x"ff480565",
			327 => x"00000565",
			328 => x"0e092408",
			329 => x"09019c04",
			330 => x"00000565",
			331 => x"00ac0565",
			332 => x"0901ee10",
			333 => x"0c06140c",
			334 => x"0d07fd04",
			335 => x"00000565",
			336 => x"01013404",
			337 => x"ff520565",
			338 => x"00000565",
			339 => x"00000565",
			340 => x"0b06cb08",
			341 => x"0a026a04",
			342 => x"00490565",
			343 => x"00000565",
			344 => x"00000565",
			345 => x"01011108",
			346 => x"06017804",
			347 => x"ff3a05c1",
			348 => x"000005c1",
			349 => x"0e09330c",
			350 => x"0409db04",
			351 => x"000005c1",
			352 => x"0c061104",
			353 => x"00b905c1",
			354 => x"000005c1",
			355 => x"040a7b0c",
			356 => x"01013c08",
			357 => x"0f098b04",
			358 => x"000005c1",
			359 => x"ff2d05c1",
			360 => x"000005c1",
			361 => x"0d086d0c",
			362 => x"00039d08",
			363 => x"0f0a4204",
			364 => x"007c05c1",
			365 => x"000005c1",
			366 => x"000005c1",
			367 => x"000005c1",
			368 => x"0209be18",
			369 => x"0a024c14",
			370 => x"0e09240c",
			371 => x"0409db04",
			372 => x"0000062d",
			373 => x"0f08d404",
			374 => x"0000062d",
			375 => x"0078062d",
			376 => x"040a4904",
			377 => x"ffd3062d",
			378 => x"0000062d",
			379 => x"fed3062d",
			380 => x"0309c014",
			381 => x"06018810",
			382 => x"0d08380c",
			383 => x"0705d204",
			384 => x"0000062d",
			385 => x"06016b04",
			386 => x"0000062d",
			387 => x"010f062d",
			388 => x"0000062d",
			389 => x"0000062d",
			390 => x"0b069c04",
			391 => x"0000062d",
			392 => x"07066e04",
			393 => x"ffb2062d",
			394 => x"0000062d",
			395 => x"02095110",
			396 => x"0f09600c",
			397 => x"06017408",
			398 => x"04091d04",
			399 => x"00000689",
			400 => x"ffa60689",
			401 => x"00000689",
			402 => x"00000689",
			403 => x"040a3a08",
			404 => x"0f099504",
			405 => x"00000689",
			406 => x"fffd0689",
			407 => x"0f0a5a14",
			408 => x"06016004",
			409 => x"00000689",
			410 => x"0c05a004",
			411 => x"00000689",
			412 => x"06018608",
			413 => x"01010604",
			414 => x"00000689",
			415 => x"00ad0689",
			416 => x"00000689",
			417 => x"00000689",
			418 => x"0c05d818",
			419 => x"0d07e40c",
			420 => x"01010b04",
			421 => x"ff8106fd",
			422 => x"020a5b04",
			423 => x"005006fd",
			424 => x"000006fd",
			425 => x"040a2808",
			426 => x"0308e704",
			427 => x"000006fd",
			428 => x"fefc06fd",
			429 => x"000006fd",
			430 => x"0d08381c",
			431 => x"0901bc04",
			432 => x"000006fd",
			433 => x"0209700c",
			434 => x"0e08e104",
			435 => x"000006fd",
			436 => x"0802a504",
			437 => x"000006fd",
			438 => x"ffcb06fd",
			439 => x"0e09c108",
			440 => x"00034604",
			441 => x"000006fd",
			442 => x"00c806fd",
			443 => x"000006fd",
			444 => x"0e096204",
			445 => x"000006fd",
			446 => x"fff006fd",
			447 => x"0901bc04",
			448 => x"00000739",
			449 => x"0d086d18",
			450 => x"0c05d804",
			451 => x"00000739",
			452 => x"06018610",
			453 => x"0e09c10c",
			454 => x"0c061a08",
			455 => x"0901d204",
			456 => x"00000739",
			457 => x"007f0739",
			458 => x"00000739",
			459 => x"00000739",
			460 => x"00000739",
			461 => x"00000739",
			462 => x"01010604",
			463 => x"00000775",
			464 => x"0b06cf18",
			465 => x"0a020804",
			466 => x"00000775",
			467 => x"0c061310",
			468 => x"07065a0c",
			469 => x"09020808",
			470 => x"0e09c104",
			471 => x"00840775",
			472 => x"00000775",
			473 => x"00000775",
			474 => x"00000775",
			475 => x"00000775",
			476 => x"00000775",
			477 => x"01011108",
			478 => x"0901b804",
			479 => x"fe7b07e1",
			480 => x"000007e1",
			481 => x"0e095110",
			482 => x"0409db08",
			483 => x"0e08e104",
			484 => x"00c507e1",
			485 => x"feb407e1",
			486 => x"0c061304",
			487 => x"017107e1",
			488 => x"000007e1",
			489 => x"0901f008",
			490 => x"0d07d604",
			491 => x"000007e1",
			492 => x"fe5f07e1",
			493 => x"0d081708",
			494 => x"0003a704",
			495 => x"011a07e1",
			496 => x"000007e1",
			497 => x"0901f608",
			498 => x"0b06f004",
			499 => x"000007e1",
			500 => x"003f07e1",
			501 => x"0b06bc04",
			502 => x"000007e1",
			503 => x"fef907e1",
			504 => x"0c05d710",
			505 => x"00036804",
			506 => x"0000085d",
			507 => x"0901ea08",
			508 => x"07062c04",
			509 => x"fe6a085d",
			510 => x"0000085d",
			511 => x"0000085d",
			512 => x"07064314",
			513 => x"0d081810",
			514 => x"02093004",
			515 => x"0000085d",
			516 => x"0901c804",
			517 => x"0000085d",
			518 => x"0e09c104",
			519 => x"00f8085d",
			520 => x"0000085d",
			521 => x"0000085d",
			522 => x"07066d0c",
			523 => x"0e091504",
			524 => x"0000085d",
			525 => x"0b06f004",
			526 => x"ff14085d",
			527 => x"0000085d",
			528 => x"05080f0c",
			529 => x"0f0a1908",
			530 => x"02097004",
			531 => x"0000085d",
			532 => x"002c085d",
			533 => x"0000085d",
			534 => x"0000085d",
			535 => x"09019c04",
			536 => x"fea308c1",
			537 => x"040a8820",
			538 => x"0e095114",
			539 => x"0409db08",
			540 => x"0e08cb04",
			541 => x"004008c1",
			542 => x"ff4708c1",
			543 => x"0c060f04",
			544 => x"011508c1",
			545 => x"00035b04",
			546 => x"004408c1",
			547 => x"ff9c08c1",
			548 => x"0f09b104",
			549 => x"000008c1",
			550 => x"040a7b04",
			551 => x"fec308c1",
			552 => x"000008c1",
			553 => x"0e09c10c",
			554 => x"0d083808",
			555 => x"06018d04",
			556 => x"017c08c1",
			557 => x"000008c1",
			558 => x"000008c1",
			559 => x"ffa908c1",
			560 => x"01010604",
			561 => x"fe630905",
			562 => x"0e09c11c",
			563 => x"0802fb18",
			564 => x"0d083110",
			565 => x"0a020804",
			566 => x"fdaa0905",
			567 => x"0003a708",
			568 => x"0c061304",
			569 => x"01cd0905",
			570 => x"00a10905",
			571 => x"03d90905",
			572 => x"0209dd04",
			573 => x"fe860905",
			574 => x"026f0905",
			575 => x"fdf00905",
			576 => x"fe650905",
			577 => x"0802fb2c",
			578 => x"0309c024",
			579 => x"040a1514",
			580 => x"0e08e108",
			581 => x"01011104",
			582 => x"00000961",
			583 => x"00af0961",
			584 => x"0b06de08",
			585 => x"0b069e04",
			586 => x"00000961",
			587 => x"ff210961",
			588 => x"00000961",
			589 => x"01010604",
			590 => x"00000961",
			591 => x"06018908",
			592 => x"0802aa04",
			593 => x"00000961",
			594 => x"015b0961",
			595 => x"00000961",
			596 => x"01014504",
			597 => x"ff130961",
			598 => x"00000961",
			599 => x"feb00961",
			600 => x"0802fb2c",
			601 => x"0309c024",
			602 => x"040a1510",
			603 => x"0e08e108",
			604 => x"01011104",
			605 => x"000009bd",
			606 => x"00a609bd",
			607 => x"00034604",
			608 => x"ff3509bd",
			609 => x"000009bd",
			610 => x"01010604",
			611 => x"000009bd",
			612 => x"0601890c",
			613 => x"0802aa04",
			614 => x"000009bd",
			615 => x"0d083804",
			616 => x"015509bd",
			617 => x"000009bd",
			618 => x"000009bd",
			619 => x"01014504",
			620 => x"ff2009bd",
			621 => x"000009bd",
			622 => x"feb709bd",
			623 => x"0c05d724",
			624 => x"0209a414",
			625 => x"0a024c10",
			626 => x"0b068d04",
			627 => x"00000a49",
			628 => x"07061404",
			629 => x"00000a49",
			630 => x"0b06be04",
			631 => x"ffcb0a49",
			632 => x"00000a49",
			633 => x"fe890a49",
			634 => x"0e09770c",
			635 => x"0b062a04",
			636 => x"00000a49",
			637 => x"020a1004",
			638 => x"00230a49",
			639 => x"00000a49",
			640 => x"00000a49",
			641 => x"0901d90c",
			642 => x"0c05f904",
			643 => x"00000a49",
			644 => x"0c061404",
			645 => x"ff630a49",
			646 => x"00000a49",
			647 => x"02096004",
			648 => x"00000a49",
			649 => x"0e096204",
			650 => x"00e50a49",
			651 => x"040abb04",
			652 => x"ffd30a49",
			653 => x"07065a08",
			654 => x"040b1c04",
			655 => x"00410a49",
			656 => x"00000a49",
			657 => x"00000a49",
			658 => x"01010b04",
			659 => x"fe650a95",
			660 => x"0309d820",
			661 => x"0e08e104",
			662 => x"01ba0a95",
			663 => x"0a023008",
			664 => x"07062a04",
			665 => x"00000a95",
			666 => x"fdb00a95",
			667 => x"01012308",
			668 => x"06017804",
			669 => x"00870a95",
			670 => x"fdfd0a95",
			671 => x"09020a08",
			672 => x"00034604",
			673 => x"ffb70a95",
			674 => x"01900a95",
			675 => x"fe4e0a95",
			676 => x"fe680a95",
			677 => x"01010604",
			678 => x"fe680b19",
			679 => x"0e095120",
			680 => x"0b06af0c",
			681 => x"040a0108",
			682 => x"0e08e104",
			683 => x"01900b19",
			684 => x"fec90b19",
			685 => x"01b80b19",
			686 => x"040a3a0c",
			687 => x"0e08e104",
			688 => x"01210b19",
			689 => x"0507ba04",
			690 => x"ff910b19",
			691 => x"fe1d0b19",
			692 => x"0209ce04",
			693 => x"01950b19",
			694 => x"00000b19",
			695 => x"0706400c",
			696 => x"040a8804",
			697 => x"fe8e0b19",
			698 => x"0e09c104",
			699 => x"01a40b19",
			700 => x"ff270b19",
			701 => x"040a5b08",
			702 => x"0802cc04",
			703 => x"fe9c0b19",
			704 => x"fb710b19",
			705 => x"0f0a1908",
			706 => x"040a8804",
			707 => x"ff6f0b19",
			708 => x"01880b19",
			709 => x"fe780b19",
			710 => x"0901a90c",
			711 => x"09019c04",
			712 => x"fe5f0b8d",
			713 => x"0901a104",
			714 => x"00000b8d",
			715 => x"feb70b8d",
			716 => x"0d083024",
			717 => x"0802f820",
			718 => x"020a2d1c",
			719 => x"0d081710",
			720 => x"0c05fa08",
			721 => x"020a1004",
			722 => x"028a0b8d",
			723 => x"03c10b8d",
			724 => x"02098e04",
			725 => x"007a0b8d",
			726 => x"023c0b8d",
			727 => x"0a023604",
			728 => x"fe630b8d",
			729 => x"0e098704",
			730 => x"02ff0b8d",
			731 => x"fea10b8d",
			732 => x"05cf0b8d",
			733 => x"fe460b8d",
			734 => x"0e096208",
			735 => x"0901ce04",
			736 => x"fe5f0b8d",
			737 => x"01920b8d",
			738 => x"fe600b8d",
			739 => x"0901bc14",
			740 => x"01010604",
			741 => x"fe720c31",
			742 => x"0802ee0c",
			743 => x"0802ae08",
			744 => x"01010f04",
			745 => x"ffcb0c31",
			746 => x"00000c31",
			747 => x"00530c31",
			748 => x"fee80c31",
			749 => x"07065824",
			750 => x"0309c018",
			751 => x"0c061310",
			752 => x"01013d08",
			753 => x"0e09a204",
			754 => x"016a0c31",
			755 => x"00000c31",
			756 => x"01013f04",
			757 => x"ffbb0c31",
			758 => x"008b0c31",
			759 => x"01012c04",
			760 => x"ff640c31",
			761 => x"00000c31",
			762 => x"01014504",
			763 => x"fea90c31",
			764 => x"0507d704",
			765 => x"009c0c31",
			766 => x"00000c31",
			767 => x"0802c308",
			768 => x"03097804",
			769 => x"00980c31",
			770 => x"00000c31",
			771 => x"0c05dc04",
			772 => x"00000c31",
			773 => x"040b1c04",
			774 => x"fe430c31",
			775 => x"01013208",
			776 => x"01012c04",
			777 => x"00000c31",
			778 => x"000c0c31",
			779 => x"ff420c31",
			780 => x"01010604",
			781 => x"fe6c0c95",
			782 => x"0e08e108",
			783 => x"06015704",
			784 => x"00000c95",
			785 => x"01940c95",
			786 => x"040a1514",
			787 => x"0409c704",
			788 => x"fe1d0c95",
			789 => x"03092e04",
			790 => x"00750c95",
			791 => x"06017708",
			792 => x"06016704",
			793 => x"00000c95",
			794 => x"fe600c95",
			795 => x"00000c95",
			796 => x"0e09c110",
			797 => x"01011f04",
			798 => x"fed30c95",
			799 => x"040a8808",
			800 => x"0e096204",
			801 => x"01570c95",
			802 => x"fe8e0c95",
			803 => x"01d80c95",
			804 => x"fe980c95",
			805 => x"01010604",
			806 => x"fe9e0d19",
			807 => x"07062a14",
			808 => x"040a150c",
			809 => x"00033e04",
			810 => x"00110d19",
			811 => x"0802a504",
			812 => x"00000d19",
			813 => x"ff6c0d19",
			814 => x"0e09a204",
			815 => x"01810d19",
			816 => x"00000d19",
			817 => x"0901f014",
			818 => x"0e09150c",
			819 => x"00031a04",
			820 => x"ff540d19",
			821 => x"00035b04",
			822 => x"009d0d19",
			823 => x"00000d19",
			824 => x"0c05bf04",
			825 => x"00000d19",
			826 => x"feed0d19",
			827 => x"0c05fa10",
			828 => x"00035304",
			829 => x"00000d19",
			830 => x"0802e808",
			831 => x"0e09c104",
			832 => x"01010d19",
			833 => x"00000d19",
			834 => x"00000d19",
			835 => x"0802c304",
			836 => x"00000d19",
			837 => x"ffe80d19",
			838 => x"0901bc08",
			839 => x"04093104",
			840 => x"00000d8d",
			841 => x"fe930d8d",
			842 => x"040a7b24",
			843 => x"0d07ee04",
			844 => x"01010d8d",
			845 => x"0c05d704",
			846 => x"fed40d8d",
			847 => x"0802c310",
			848 => x"0e095108",
			849 => x"0802ae04",
			850 => x"00000d8d",
			851 => x"01120d8d",
			852 => x"040a5b04",
			853 => x"ff910d8d",
			854 => x"00000d8d",
			855 => x"00035b04",
			856 => x"00000d8d",
			857 => x"0c05f404",
			858 => x"00000d8d",
			859 => x"ff150d8d",
			860 => x"0d086d0c",
			861 => x"01011f04",
			862 => x"00000d8d",
			863 => x"0e09c104",
			864 => x"01b20d8d",
			865 => x"00000d8d",
			866 => x"ff760d8d",
			867 => x"0802e640",
			868 => x"0d082220",
			869 => x"06015204",
			870 => x"fe660e31",
			871 => x"0c061318",
			872 => x"040a5b10",
			873 => x"0e093308",
			874 => x"03091a04",
			875 => x"02190e31",
			876 => x"01b70e31",
			877 => x"02099504",
			878 => x"fffe0e31",
			879 => x"fe150e31",
			880 => x"020a1004",
			881 => x"02180e31",
			882 => x"02c50e31",
			883 => x"00960e31",
			884 => x"0507bc08",
			885 => x"0002e604",
			886 => x"feed0e31",
			887 => x"02c10e31",
			888 => x"0c05f70c",
			889 => x"00036304",
			890 => x"fe730e31",
			891 => x"06018104",
			892 => x"02ed0e31",
			893 => x"ff000e31",
			894 => x"0507e408",
			895 => x"0507d904",
			896 => x"fe720e31",
			897 => x"00e10e31",
			898 => x"fe650e31",
			899 => x"0802fb10",
			900 => x"0e09a20c",
			901 => x"0c059b04",
			902 => x"fe750e31",
			903 => x"040b7804",
			904 => x"01500e31",
			905 => x"02d40e31",
			906 => x"fe680e31",
			907 => x"fe600e31",
			908 => x"01010604",
			909 => x"fe990ebd",
			910 => x"07062a14",
			911 => x"040a150c",
			912 => x"00033e04",
			913 => x"00150ebd",
			914 => x"0802a504",
			915 => x"00000ebd",
			916 => x"ff590ebd",
			917 => x"0e09a204",
			918 => x"018b0ebd",
			919 => x"00000ebd",
			920 => x"0901f018",
			921 => x"0e091510",
			922 => x"00031a04",
			923 => x"ff4b0ebd",
			924 => x"00035b08",
			925 => x"02092804",
			926 => x"00000ebd",
			927 => x"00c00ebd",
			928 => x"00000ebd",
			929 => x"0c05bf04",
			930 => x"00000ebd",
			931 => x"fedc0ebd",
			932 => x"0c05fa10",
			933 => x"00035304",
			934 => x"00000ebd",
			935 => x"0802e808",
			936 => x"0e09c104",
			937 => x"010b0ebd",
			938 => x"00000ebd",
			939 => x"00000ebd",
			940 => x"0802c304",
			941 => x"00000ebd",
			942 => x"ffe10ebd",
			943 => x"01010604",
			944 => x"fe660f19",
			945 => x"030a0128",
			946 => x"03091a04",
			947 => x"01b00f19",
			948 => x"040a010c",
			949 => x"0f095608",
			950 => x"02093504",
			951 => x"feea0f19",
			952 => x"00000f19",
			953 => x"fdae0f19",
			954 => x"01011f08",
			955 => x"05079e04",
			956 => x"00000f19",
			957 => x"fe610f19",
			958 => x"040a5b08",
			959 => x"06017904",
			960 => x"00dd0f19",
			961 => x"fd210f19",
			962 => x"06018d04",
			963 => x"01d10f19",
			964 => x"ff380f19",
			965 => x"fe6f0f19",
			966 => x"01010604",
			967 => x"fe6b0f8d",
			968 => x"0e08e108",
			969 => x"06015704",
			970 => x"00000f8d",
			971 => x"01990f8d",
			972 => x"040a1518",
			973 => x"0409db04",
			974 => x"fe330f8d",
			975 => x"03092e08",
			976 => x"0901e604",
			977 => x"00000f8d",
			978 => x"00c50f8d",
			979 => x"06017708",
			980 => x"06016704",
			981 => x"00000f8d",
			982 => x"fe730f8d",
			983 => x"00000f8d",
			984 => x"0e09c114",
			985 => x"01011f04",
			986 => x"fec20f8d",
			987 => x"040a8808",
			988 => x"0e096204",
			989 => x"01600f8d",
			990 => x"fe820f8d",
			991 => x"06018904",
			992 => x"01f20f8d",
			993 => x"00000f8d",
			994 => x"fe920f8d",
			995 => x"01010604",
			996 => x"fe691021",
			997 => x"07062c1c",
			998 => x"040b9d14",
			999 => x"03092204",
			1000 => x"01971021",
			1001 => x"040a0104",
			1002 => x"fe461021",
			1003 => x"0e09c108",
			1004 => x"040a2804",
			1005 => x"00001021",
			1006 => x"01851021",
			1007 => x"ffbe1021",
			1008 => x"040bd804",
			1009 => x"047d1021",
			1010 => x"00001021",
			1011 => x"0e095114",
			1012 => x"0a022b08",
			1013 => x"03091a04",
			1014 => x"005e1021",
			1015 => x"fe5e1021",
			1016 => x"0901c804",
			1017 => x"ff031021",
			1018 => x"02093a04",
			1019 => x"00131021",
			1020 => x"019f1021",
			1021 => x"03098704",
			1022 => x"fd891021",
			1023 => x"0507e410",
			1024 => x"07064008",
			1025 => x"0309d804",
			1026 => x"00941021",
			1027 => x"00001021",
			1028 => x"0b06e004",
			1029 => x"ff411021",
			1030 => x"00001021",
			1031 => x"fe8c1021",
			1032 => x"01010604",
			1033 => x"fe6f10ad",
			1034 => x"0e08e108",
			1035 => x"06015704",
			1036 => x"000010ad",
			1037 => x"018a10ad",
			1038 => x"01012410",
			1039 => x"0901d90c",
			1040 => x"07064204",
			1041 => x"fe8110ad",
			1042 => x"0c05fa04",
			1043 => x"000010ad",
			1044 => x"ff6610ad",
			1045 => x"000010ad",
			1046 => x"07065814",
			1047 => x"040a7b0c",
			1048 => x"0e095108",
			1049 => x"0409db04",
			1050 => x"fee610ad",
			1051 => x"013510ad",
			1052 => x"fe8710ad",
			1053 => x"0e09c104",
			1054 => x"01be10ad",
			1055 => x"ff9210ad",
			1056 => x"0c05f40c",
			1057 => x"00035b04",
			1058 => x"000010ad",
			1059 => x"09020204",
			1060 => x"010910ad",
			1061 => x"000010ad",
			1062 => x"0802be04",
			1063 => x"000010ad",
			1064 => x"040b1c04",
			1065 => x"fe0d10ad",
			1066 => x"ff8b10ad",
			1067 => x"01010604",
			1068 => x"fe631123",
			1069 => x"0e09c134",
			1070 => x"0802fb30",
			1071 => x"040a3a1c",
			1072 => x"0e08fd0c",
			1073 => x"01011104",
			1074 => x"fd991123",
			1075 => x"01013404",
			1076 => x"01da1123",
			1077 => x"00e41123",
			1078 => x"040a0108",
			1079 => x"0a023604",
			1080 => x"fe921123",
			1081 => x"fce51123",
			1082 => x"0c05f904",
			1083 => x"01371123",
			1084 => x"fd8b1123",
			1085 => x"020a2d10",
			1086 => x"0d082208",
			1087 => x"0f09e104",
			1088 => x"01e61123",
			1089 => x"01421123",
			1090 => x"0f09e104",
			1091 => x"00171123",
			1092 => x"ff0c1123",
			1093 => x"03bf1123",
			1094 => x"fdfd1123",
			1095 => x"fe661123",
			1096 => x"00001125",
			1097 => x"00001129",
			1098 => x"0000112d",
			1099 => x"00001131",
			1100 => x"00001135",
			1101 => x"00001139",
			1102 => x"0000113d",
			1103 => x"00001141",
			1104 => x"00001145",
			1105 => x"00001149",
			1106 => x"0000114d",
			1107 => x"00001151",
			1108 => x"00001155",
			1109 => x"00001159",
			1110 => x"0000115d",
			1111 => x"00001161",
			1112 => x"00001165",
			1113 => x"00001169",
			1114 => x"0000116d",
			1115 => x"00001171",
			1116 => x"00001175",
			1117 => x"00001179",
			1118 => x"0000117d",
			1119 => x"00001181",
			1120 => x"00001185",
			1121 => x"00001189",
			1122 => x"0000118d",
			1123 => x"0802e604",
			1124 => x"00001199",
			1125 => x"ffb71199",
			1126 => x"0802be04",
			1127 => x"000011a5",
			1128 => x"ffed11a5",
			1129 => x"01013704",
			1130 => x"fff911b1",
			1131 => x"000011b1",
			1132 => x"0e08e108",
			1133 => x"0e081604",
			1134 => x"000011c5",
			1135 => x"002b11c5",
			1136 => x"fff511c5",
			1137 => x"0802e608",
			1138 => x"040a5b04",
			1139 => x"000011d9",
			1140 => x"002511d9",
			1141 => x"ffac11d9",
			1142 => x"0e093304",
			1143 => x"000011ed",
			1144 => x"0f099504",
			1145 => x"000011ed",
			1146 => x"fff811ed",
			1147 => x"01011104",
			1148 => x"ffc41209",
			1149 => x"01014908",
			1150 => x"01011304",
			1151 => x"00001209",
			1152 => x"00091209",
			1153 => x"00001209",
			1154 => x"0802e60c",
			1155 => x"01011104",
			1156 => x"00001225",
			1157 => x"09020804",
			1158 => x"00381225",
			1159 => x"00001225",
			1160 => x"00001225",
			1161 => x"01012408",
			1162 => x"0901d904",
			1163 => x"ffe11249",
			1164 => x"00001249",
			1165 => x"02097004",
			1166 => x"00001249",
			1167 => x"020a6b04",
			1168 => x"001c1249",
			1169 => x"00001249",
			1170 => x"0e08e10c",
			1171 => x"09019c04",
			1172 => x"00001275",
			1173 => x"00030204",
			1174 => x"00001275",
			1175 => x"00351275",
			1176 => x"01013f08",
			1177 => x"0c059f04",
			1178 => x"00001275",
			1179 => x"ffad1275",
			1180 => x"00001275",
			1181 => x"0901bc04",
			1182 => x"ffa91299",
			1183 => x"0601860c",
			1184 => x"06015704",
			1185 => x"00001299",
			1186 => x"09020504",
			1187 => x"00301299",
			1188 => x"00001299",
			1189 => x"00001299",
			1190 => x"01011704",
			1191 => x"000012bd",
			1192 => x"0902080c",
			1193 => x"0802fb08",
			1194 => x"0802aa04",
			1195 => x"000012bd",
			1196 => x"002612bd",
			1197 => x"000012bd",
			1198 => x"000012bd",
			1199 => x"0901f010",
			1200 => x"0e08e104",
			1201 => x"000012e1",
			1202 => x"040b6b08",
			1203 => x"03092204",
			1204 => x"000012e1",
			1205 => x"ffc812e1",
			1206 => x"000012e1",
			1207 => x"000012e1",
			1208 => x"0901d908",
			1209 => x"0b06ae04",
			1210 => x"0000130d",
			1211 => x"ffa8130d",
			1212 => x"0c05da04",
			1213 => x"0000130d",
			1214 => x"0d082208",
			1215 => x"0a026204",
			1216 => x"0078130d",
			1217 => x"0000130d",
			1218 => x"0000130d",
			1219 => x"0e08e110",
			1220 => x"0e081604",
			1221 => x"00001341",
			1222 => x"0d080108",
			1223 => x"020a0604",
			1224 => x"00401341",
			1225 => x"00001341",
			1226 => x"00001341",
			1227 => x"040a5b08",
			1228 => x"0d07d604",
			1229 => x"00001341",
			1230 => x"ffb61341",
			1231 => x"00001341",
			1232 => x"0901bc04",
			1233 => x"ffaf136d",
			1234 => x"06018610",
			1235 => x"06015704",
			1236 => x"0000136d",
			1237 => x"09020508",
			1238 => x"01011304",
			1239 => x"0000136d",
			1240 => x"002b136d",
			1241 => x"0000136d",
			1242 => x"0000136d",
			1243 => x"0901d90c",
			1244 => x"0802a504",
			1245 => x"000013a9",
			1246 => x"0c05b804",
			1247 => x"ffe213a9",
			1248 => x"000013a9",
			1249 => x"0802d710",
			1250 => x"0c05d804",
			1251 => x"000013a9",
			1252 => x"09020808",
			1253 => x"0c061004",
			1254 => x"006813a9",
			1255 => x"000013a9",
			1256 => x"000013a9",
			1257 => x"000013a9",
			1258 => x"0901bc08",
			1259 => x"04091d04",
			1260 => x"000013ed",
			1261 => x"ffa613ed",
			1262 => x"0e093310",
			1263 => x"0409db04",
			1264 => x"000013ed",
			1265 => x"0a022b04",
			1266 => x"000013ed",
			1267 => x"0a024504",
			1268 => x"00a413ed",
			1269 => x"000013ed",
			1270 => x"040a6908",
			1271 => x"0f099504",
			1272 => x"000013ed",
			1273 => x"ff8813ed",
			1274 => x"000013ed",
			1275 => x"0209a41c",
			1276 => x"0e08e10c",
			1277 => x"01011108",
			1278 => x"02093d04",
			1279 => x"ffb91449",
			1280 => x"00001449",
			1281 => x"005e1449",
			1282 => x"040a280c",
			1283 => x"0b06ce08",
			1284 => x"0c061404",
			1285 => x"ff281449",
			1286 => x"00001449",
			1287 => x"00001449",
			1288 => x"00001449",
			1289 => x"0e09870c",
			1290 => x"09019c04",
			1291 => x"00001449",
			1292 => x"040a4904",
			1293 => x"00001449",
			1294 => x"00b71449",
			1295 => x"01013904",
			1296 => x"ffc51449",
			1297 => x"00001449",
			1298 => x"0901bc08",
			1299 => x"06017804",
			1300 => x"ff431495",
			1301 => x"00001495",
			1302 => x"0e093310",
			1303 => x"0101360c",
			1304 => x"0507bc08",
			1305 => x"0e092404",
			1306 => x"00ce1495",
			1307 => x"00001495",
			1308 => x"00001495",
			1309 => x"00001495",
			1310 => x"0101370c",
			1311 => x"0a025b08",
			1312 => x"0f098b04",
			1313 => x"00001495",
			1314 => x"ff441495",
			1315 => x"00001495",
			1316 => x"00001495",
			1317 => x"0c05b804",
			1318 => x"000014c9",
			1319 => x"0d083814",
			1320 => x"0a022b04",
			1321 => x"000014c9",
			1322 => x"0601880c",
			1323 => x"040a2804",
			1324 => x"000014c9",
			1325 => x"09019c04",
			1326 => x"000014c9",
			1327 => x"00b314c9",
			1328 => x"000014c9",
			1329 => x"000014c9",
			1330 => x"0c05d710",
			1331 => x"0e08e104",
			1332 => x"00001515",
			1333 => x"0b066c04",
			1334 => x"00001515",
			1335 => x"0d081704",
			1336 => x"ffdc1515",
			1337 => x"00001515",
			1338 => x"0d083814",
			1339 => x"0c061310",
			1340 => x"0601880c",
			1341 => x"01011104",
			1342 => x"00001515",
			1343 => x"0d083104",
			1344 => x"00a01515",
			1345 => x"00001515",
			1346 => x"00001515",
			1347 => x"00001515",
			1348 => x"00001515",
			1349 => x"02097010",
			1350 => x"0e08e104",
			1351 => x"00001571",
			1352 => x"06017408",
			1353 => x"0f097d04",
			1354 => x"ffa51571",
			1355 => x"00001571",
			1356 => x"00001571",
			1357 => x"0f099510",
			1358 => x"040a0104",
			1359 => x"00001571",
			1360 => x"0a026d08",
			1361 => x"06016304",
			1362 => x"00001571",
			1363 => x"00821571",
			1364 => x"00001571",
			1365 => x"040ae20c",
			1366 => x"0e092404",
			1367 => x"00001571",
			1368 => x"0d07d604",
			1369 => x"00001571",
			1370 => x"ffbc1571",
			1371 => x"00001571",
			1372 => x"0c05d710",
			1373 => x"0a024c04",
			1374 => x"000015d5",
			1375 => x"01013808",
			1376 => x"07062c04",
			1377 => x"fee215d5",
			1378 => x"000015d5",
			1379 => x"000015d5",
			1380 => x"07062c0c",
			1381 => x"02092804",
			1382 => x"000015d5",
			1383 => x"0a027504",
			1384 => x"00d015d5",
			1385 => x"000015d5",
			1386 => x"0c05f90c",
			1387 => x"0d081708",
			1388 => x"01011304",
			1389 => x"000015d5",
			1390 => x"005d15d5",
			1391 => x"000015d5",
			1392 => x"0802c304",
			1393 => x"000015d5",
			1394 => x"040b1c04",
			1395 => x"ff3a15d5",
			1396 => x"000015d5",
			1397 => x"0c05d818",
			1398 => x"0d07ee0c",
			1399 => x"09019c04",
			1400 => x"ffab1649",
			1401 => x"0e095104",
			1402 => x"00911649",
			1403 => x"00001649",
			1404 => x"0b06ac04",
			1405 => x"00001649",
			1406 => x"07061704",
			1407 => x"00001649",
			1408 => x"ff371649",
			1409 => x"07063f0c",
			1410 => x"0901c604",
			1411 => x"00001649",
			1412 => x"0e09c104",
			1413 => x"00b41649",
			1414 => x"00001649",
			1415 => x"0802d70c",
			1416 => x"0802aa04",
			1417 => x"00001649",
			1418 => x"0c061a04",
			1419 => x"005b1649",
			1420 => x"00001649",
			1421 => x"0c05dc04",
			1422 => x"00001649",
			1423 => x"0901ea04",
			1424 => x"00001649",
			1425 => x"ff961649",
			1426 => x"0c05d710",
			1427 => x"0a024c04",
			1428 => x"000016b5",
			1429 => x"01013808",
			1430 => x"07062c04",
			1431 => x"fed416b5",
			1432 => x"000016b5",
			1433 => x"000016b5",
			1434 => x"07062c10",
			1435 => x"02092804",
			1436 => x"000016b5",
			1437 => x"0a027508",
			1438 => x"01011904",
			1439 => x"000016b5",
			1440 => x"00da16b5",
			1441 => x"000016b5",
			1442 => x"0c05f90c",
			1443 => x"0d081708",
			1444 => x"01011304",
			1445 => x"000016b5",
			1446 => x"006216b5",
			1447 => x"000016b5",
			1448 => x"0802c304",
			1449 => x"000016b5",
			1450 => x"040b1c04",
			1451 => x"ff2d16b5",
			1452 => x"000016b5",
			1453 => x"0209510c",
			1454 => x"06017408",
			1455 => x"04091d04",
			1456 => x"00001701",
			1457 => x"ffb91701",
			1458 => x"00001701",
			1459 => x"040a3a04",
			1460 => x"00001701",
			1461 => x"06018614",
			1462 => x"0c05a004",
			1463 => x"00001701",
			1464 => x"0a023604",
			1465 => x"00001701",
			1466 => x"020a6b08",
			1467 => x"01010604",
			1468 => x"00001701",
			1469 => x"00a51701",
			1470 => x"00001701",
			1471 => x"00001701",
			1472 => x"0f099520",
			1473 => x"0705e80c",
			1474 => x"01010f08",
			1475 => x"0d079604",
			1476 => x"ff88176d",
			1477 => x"0000176d",
			1478 => x"0000176d",
			1479 => x"0409db0c",
			1480 => x"0308f704",
			1481 => x"0000176d",
			1482 => x"0e08e104",
			1483 => x"0000176d",
			1484 => x"ffc9176d",
			1485 => x"01010604",
			1486 => x"0000176d",
			1487 => x"00ce176d",
			1488 => x"0c061214",
			1489 => x"01013410",
			1490 => x"0e092404",
			1491 => x"0000176d",
			1492 => x"0d07d604",
			1493 => x"0000176d",
			1494 => x"0901ee04",
			1495 => x"ff25176d",
			1496 => x"0000176d",
			1497 => x"0000176d",
			1498 => x"0000176d",
			1499 => x"0802fb28",
			1500 => x"040a5b18",
			1501 => x"0e092410",
			1502 => x"0a020804",
			1503 => x"000017c1",
			1504 => x"0d080a08",
			1505 => x"01011104",
			1506 => x"000017c1",
			1507 => x"00bb17c1",
			1508 => x"000017c1",
			1509 => x"0901f804",
			1510 => x"ff0d17c1",
			1511 => x"000017c1",
			1512 => x"0d086d0c",
			1513 => x"01010604",
			1514 => x"000017c1",
			1515 => x"0e09c104",
			1516 => x"00ea17c1",
			1517 => x"000017c1",
			1518 => x"000017c1",
			1519 => x"ff7c17c1",
			1520 => x"0c05b80c",
			1521 => x"01012108",
			1522 => x"08029104",
			1523 => x"0000182d",
			1524 => x"ff8a182d",
			1525 => x"0000182d",
			1526 => x"0e08fd0c",
			1527 => x"0a020004",
			1528 => x"0000182d",
			1529 => x"09019c04",
			1530 => x"0000182d",
			1531 => x"00ac182d",
			1532 => x"040a5b10",
			1533 => x"0901f20c",
			1534 => x"0c05d504",
			1535 => x"0000182d",
			1536 => x"01012804",
			1537 => x"0000182d",
			1538 => x"ff75182d",
			1539 => x"0000182d",
			1540 => x"0309d80c",
			1541 => x"01011f04",
			1542 => x"0000182d",
			1543 => x"0c05d604",
			1544 => x"0000182d",
			1545 => x"0087182d",
			1546 => x"0000182d",
			1547 => x"0901bc04",
			1548 => x"00001869",
			1549 => x"05080418",
			1550 => x"00031a04",
			1551 => x"00001869",
			1552 => x"06018810",
			1553 => x"0e09c10c",
			1554 => x"0705ff04",
			1555 => x"00001869",
			1556 => x"07067004",
			1557 => x"004b1869",
			1558 => x"00001869",
			1559 => x"00001869",
			1560 => x"00001869",
			1561 => x"00001869",
			1562 => x"0c05d818",
			1563 => x"00036810",
			1564 => x"0d07e404",
			1565 => x"000018dd",
			1566 => x"0507ad08",
			1567 => x"05079c04",
			1568 => x"000018dd",
			1569 => x"ffd018dd",
			1570 => x"000018dd",
			1571 => x"0209a404",
			1572 => x"ff2b18dd",
			1573 => x"000018dd",
			1574 => x"0d08381c",
			1575 => x"0901bc04",
			1576 => x"000018dd",
			1577 => x"0209700c",
			1578 => x"0e08e104",
			1579 => x"000018dd",
			1580 => x"01012804",
			1581 => x"000018dd",
			1582 => x"ffcb18dd",
			1583 => x"0e09c108",
			1584 => x"00034604",
			1585 => x"000018dd",
			1586 => x"00be18dd",
			1587 => x"000018dd",
			1588 => x"0e096204",
			1589 => x"000018dd",
			1590 => x"fffe18dd",
			1591 => x"0901bc0c",
			1592 => x"06017808",
			1593 => x"04091d04",
			1594 => x"00001949",
			1595 => x"ff481949",
			1596 => x"00001949",
			1597 => x"0e093310",
			1598 => x"0409db04",
			1599 => x"00001949",
			1600 => x"0802c308",
			1601 => x"0802aa04",
			1602 => x"00001949",
			1603 => x"00a51949",
			1604 => x"00001949",
			1605 => x"040a5b08",
			1606 => x"0f098b04",
			1607 => x"00001949",
			1608 => x"ff2c1949",
			1609 => x"0802e610",
			1610 => x"040a7b04",
			1611 => x"00001949",
			1612 => x"0d086d08",
			1613 => x"0f0a4204",
			1614 => x"008c1949",
			1615 => x"00001949",
			1616 => x"00001949",
			1617 => x"00001949",
			1618 => x"0c05d710",
			1619 => x"0a024c04",
			1620 => x"000019c5",
			1621 => x"0901ea08",
			1622 => x"07062c04",
			1623 => x"fe7a19c5",
			1624 => x"000019c5",
			1625 => x"000019c5",
			1626 => x"07064314",
			1627 => x"0d081810",
			1628 => x"02093004",
			1629 => x"000019c5",
			1630 => x"0901c804",
			1631 => x"000019c5",
			1632 => x"0e09c104",
			1633 => x"00f219c5",
			1634 => x"000019c5",
			1635 => x"000019c5",
			1636 => x"07066d0c",
			1637 => x"0e091504",
			1638 => x"000019c5",
			1639 => x"0507f604",
			1640 => x"ff2d19c5",
			1641 => x"000019c5",
			1642 => x"05080f0c",
			1643 => x"0f0a1908",
			1644 => x"02097004",
			1645 => x"000019c5",
			1646 => x"002b19c5",
			1647 => x"000019c5",
			1648 => x"000019c5",
			1649 => x"0901a904",
			1650 => x"fe671a19",
			1651 => x"0e096218",
			1652 => x"0e08e104",
			1653 => x"01a71a19",
			1654 => x"0409db04",
			1655 => x"fdd01a19",
			1656 => x"0901d204",
			1657 => x"feb71a19",
			1658 => x"06018108",
			1659 => x"0802aa04",
			1660 => x"00611a19",
			1661 => x"01b71a19",
			1662 => x"00621a19",
			1663 => x"0e09c10c",
			1664 => x"0901f204",
			1665 => x"fe6c1a19",
			1666 => x"040a8804",
			1667 => x"fe9f1a19",
			1668 => x"01ce1a19",
			1669 => x"fe731a19",
			1670 => x"0209be24",
			1671 => x"0a024c20",
			1672 => x"0802aa14",
			1673 => x"0b069e04",
			1674 => x"00001a85",
			1675 => x"0706590c",
			1676 => x"0308f704",
			1677 => x"00001a85",
			1678 => x"0e08cb04",
			1679 => x"00001a85",
			1680 => x"ff671a85",
			1681 => x"00001a85",
			1682 => x"0e096208",
			1683 => x"01010b04",
			1684 => x"00001a85",
			1685 => x"00c21a85",
			1686 => x"00001a85",
			1687 => x"ff121a85",
			1688 => x"0d086d10",
			1689 => x"0802fb0c",
			1690 => x"040abb04",
			1691 => x"00001a85",
			1692 => x"0e09c104",
			1693 => x"01071a85",
			1694 => x"00001a85",
			1695 => x"00001a85",
			1696 => x"00001a85",
			1697 => x"0802f834",
			1698 => x"0e08fd14",
			1699 => x"02091308",
			1700 => x"01011104",
			1701 => x"ff4a1af1",
			1702 => x"00001af1",
			1703 => x"03092e08",
			1704 => x"01010604",
			1705 => x"00001af1",
			1706 => x"01581af1",
			1707 => x"00001af1",
			1708 => x"01013410",
			1709 => x"0b069c04",
			1710 => x"00001af1",
			1711 => x"07065b08",
			1712 => x"06016c04",
			1713 => x"00001af1",
			1714 => x"feb51af1",
			1715 => x"00001af1",
			1716 => x"0802dd0c",
			1717 => x"040a2804",
			1718 => x"00001af1",
			1719 => x"0b06d204",
			1720 => x"011c1af1",
			1721 => x"00001af1",
			1722 => x"ffae1af1",
			1723 => x"fe841af1",
			1724 => x"01011108",
			1725 => x"0901b804",
			1726 => x"fe7e1b65",
			1727 => x"00001b65",
			1728 => x"0e095110",
			1729 => x"0409db08",
			1730 => x"0e08e104",
			1731 => x"00ba1b65",
			1732 => x"fec91b65",
			1733 => x"0c061304",
			1734 => x"016c1b65",
			1735 => x"00001b65",
			1736 => x"0901f008",
			1737 => x"05078104",
			1738 => x"00001b65",
			1739 => x"fe6d1b65",
			1740 => x"0b06cb0c",
			1741 => x"0c05fc08",
			1742 => x"06018d04",
			1743 => x"01041b65",
			1744 => x"00001b65",
			1745 => x"00001b65",
			1746 => x"01013a0c",
			1747 => x"07066e04",
			1748 => x"00001b65",
			1749 => x"0b06fc04",
			1750 => x"003f1b65",
			1751 => x"00001b65",
			1752 => x"ff231b65",
			1753 => x"0901bc14",
			1754 => x"00039a10",
			1755 => x"0901a904",
			1756 => x"ff121be9",
			1757 => x"0802ae08",
			1758 => x"00031a04",
			1759 => x"00001be9",
			1760 => x"fff31be9",
			1761 => x"003c1be9",
			1762 => x"fe6f1be9",
			1763 => x"0309c024",
			1764 => x"040a7b1c",
			1765 => x"0e095114",
			1766 => x"0c06110c",
			1767 => x"0901fc08",
			1768 => x"0507cc04",
			1769 => x"01601be9",
			1770 => x"00001be9",
			1771 => x"00001be9",
			1772 => x"0802a504",
			1773 => x"00001be9",
			1774 => x"ff9a1be9",
			1775 => x"0f09a304",
			1776 => x"00001be9",
			1777 => x"fe5b1be9",
			1778 => x"06018a04",
			1779 => x"019d1be9",
			1780 => x"00001be9",
			1781 => x"0507bc08",
			1782 => x"09020504",
			1783 => x"ff221be9",
			1784 => x"00901be9",
			1785 => x"feb31be9",
			1786 => x"01010604",
			1787 => x"fe5c1c55",
			1788 => x"0d082220",
			1789 => x"0e09c11c",
			1790 => x"01013c14",
			1791 => x"0d080e0c",
			1792 => x"08028704",
			1793 => x"058c1c55",
			1794 => x"0b06cc04",
			1795 => x"03471c55",
			1796 => x"04d41c55",
			1797 => x"040a2804",
			1798 => x"ff701c55",
			1799 => x"03541c55",
			1800 => x"0901fe04",
			1801 => x"05e91c55",
			1802 => x"032f1c55",
			1803 => x"fe821c55",
			1804 => x"0e098708",
			1805 => x"01013004",
			1806 => x"fe4c1c55",
			1807 => x"03201c55",
			1808 => x"0e09c108",
			1809 => x"0f0a0304",
			1810 => x"fe7c1c55",
			1811 => x"01231c55",
			1812 => x"fe5d1c55",
			1813 => x"01010b04",
			1814 => x"fe651ca1",
			1815 => x"0309d820",
			1816 => x"0e08e104",
			1817 => x"01b31ca1",
			1818 => x"040a0108",
			1819 => x"03092204",
			1820 => x"ffa41ca1",
			1821 => x"fdae1ca1",
			1822 => x"0901d204",
			1823 => x"ff061ca1",
			1824 => x"0e09a208",
			1825 => x"07065a04",
			1826 => x"019f1ca1",
			1827 => x"00341ca1",
			1828 => x"040acf04",
			1829 => x"fe7f1ca1",
			1830 => x"01a61ca1",
			1831 => x"fe6a1ca1",
			1832 => x"0802fb38",
			1833 => x"040adc28",
			1834 => x"0e092418",
			1835 => x"06015708",
			1836 => x"02090c04",
			1837 => x"ffad1d15",
			1838 => x"00001d15",
			1839 => x"0a02490c",
			1840 => x"0901f608",
			1841 => x"0901b804",
			1842 => x"00001d15",
			1843 => x"01031d15",
			1844 => x"00001d15",
			1845 => x"00001d15",
			1846 => x"0901ec0c",
			1847 => x"0507d908",
			1848 => x"0d07ee04",
			1849 => x"00001d15",
			1850 => x"feba1d15",
			1851 => x"00001d15",
			1852 => x"00001d15",
			1853 => x"0508040c",
			1854 => x"09019c04",
			1855 => x"00001d15",
			1856 => x"0e09e004",
			1857 => x"01411d15",
			1858 => x"00001d15",
			1859 => x"00001d15",
			1860 => x"fec41d15",
			1861 => x"0901bc14",
			1862 => x"00039a10",
			1863 => x"01010604",
			1864 => x"fef11dc1",
			1865 => x"00035308",
			1866 => x"01010f04",
			1867 => x"ffcb1dc1",
			1868 => x"00001dc1",
			1869 => x"00561dc1",
			1870 => x"fe6c1dc1",
			1871 => x"07065824",
			1872 => x"0309c018",
			1873 => x"0c061310",
			1874 => x"01013d08",
			1875 => x"0e09a204",
			1876 => x"01751dc1",
			1877 => x"00001dc1",
			1878 => x"01013f04",
			1879 => x"ffa41dc1",
			1880 => x"00931dc1",
			1881 => x"0c061404",
			1882 => x"ff761dc1",
			1883 => x"00001dc1",
			1884 => x"01014504",
			1885 => x"fe9c1dc1",
			1886 => x"0507d704",
			1887 => x"00a51dc1",
			1888 => x"00001dc1",
			1889 => x"0a02490c",
			1890 => x"03099608",
			1891 => x"00032c04",
			1892 => x"00001dc1",
			1893 => x"00b91dc1",
			1894 => x"00001dc1",
			1895 => x"040b1c04",
			1896 => x"fe321dc1",
			1897 => x"00039d08",
			1898 => x"09021804",
			1899 => x"00261dc1",
			1900 => x"00001dc1",
			1901 => x"0c05dc04",
			1902 => x"00001dc1",
			1903 => x"ff241dc1",
			1904 => x"0802f838",
			1905 => x"0e08e10c",
			1906 => x"06015204",
			1907 => x"ff4f1e35",
			1908 => x"01010604",
			1909 => x"00001e35",
			1910 => x"015e1e35",
			1911 => x"0c05f91c",
			1912 => x"040a150c",
			1913 => x"0802ae08",
			1914 => x"06016804",
			1915 => x"00001e35",
			1916 => x"fef31e35",
			1917 => x"00001e35",
			1918 => x"0e097704",
			1919 => x"01291e35",
			1920 => x"01013b04",
			1921 => x"feee1e35",
			1922 => x"040aa904",
			1923 => x"00001e35",
			1924 => x"00a71e35",
			1925 => x"07063f04",
			1926 => x"00001e35",
			1927 => x"040b4a08",
			1928 => x"06016c04",
			1929 => x"00001e35",
			1930 => x"fe811e35",
			1931 => x"00001e35",
			1932 => x"fe811e35",
			1933 => x"01010604",
			1934 => x"fea91ec9",
			1935 => x"07062e20",
			1936 => x"040a7b14",
			1937 => x"03094008",
			1938 => x"01013704",
			1939 => x"00bd1ec9",
			1940 => x"00001ec9",
			1941 => x"0c05f308",
			1942 => x"0d07e404",
			1943 => x"00001ec9",
			1944 => x"ff6c1ec9",
			1945 => x"00001ec9",
			1946 => x"0e09c108",
			1947 => x"0c057f04",
			1948 => x"00001ec9",
			1949 => x"016c1ec9",
			1950 => x"00001ec9",
			1951 => x"0c05f310",
			1952 => x"0802b308",
			1953 => x"03092e04",
			1954 => x"00001ec9",
			1955 => x"ffce1ec9",
			1956 => x"0802e804",
			1957 => x"00d21ec9",
			1958 => x"00001ec9",
			1959 => x"0e09150c",
			1960 => x"0d080a04",
			1961 => x"00491ec9",
			1962 => x"0a022b04",
			1963 => x"ffe31ec9",
			1964 => x"00001ec9",
			1965 => x"07064104",
			1966 => x"00001ec9",
			1967 => x"0802c304",
			1968 => x"00001ec9",
			1969 => x"fecb1ec9",
			1970 => x"01010b04",
			1971 => x"fe641f1d",
			1972 => x"0309d824",
			1973 => x"0e08e104",
			1974 => x"01c31f1d",
			1975 => x"040a010c",
			1976 => x"03092204",
			1977 => x"ff941f1d",
			1978 => x"03094f04",
			1979 => x"fd091f1d",
			1980 => x"fe961f1d",
			1981 => x"0901d204",
			1982 => x"fed21f1d",
			1983 => x"0e09a208",
			1984 => x"07065a04",
			1985 => x"01c01f1d",
			1986 => x"00741f1d",
			1987 => x"040acf04",
			1988 => x"fe7a1f1d",
			1989 => x"01f31f1d",
			1990 => x"fe671f1d",
			1991 => x"01010604",
			1992 => x"fe601f81",
			1993 => x"0d083024",
			1994 => x"0802f820",
			1995 => x"020a2d1c",
			1996 => x"0d081710",
			1997 => x"0c05fa08",
			1998 => x"040a2804",
			1999 => x"02261f81",
			2000 => x"026c1f81",
			2001 => x"02098e04",
			2002 => x"00601f81",
			2003 => x"01f21f81",
			2004 => x"00035304",
			2005 => x"fe741f81",
			2006 => x"06018104",
			2007 => x"026d1f81",
			2008 => x"fec31f81",
			2009 => x"04711f81",
			2010 => x"fe461f81",
			2011 => x"0309c008",
			2012 => x"01012e04",
			2013 => x"fe611f81",
			2014 => x"010e1f81",
			2015 => x"fe611f81",
			2016 => x"01010604",
			2017 => x"fe661fe5",
			2018 => x"0e09c12c",
			2019 => x"03091a08",
			2020 => x"01010f04",
			2021 => x"02c71fe5",
			2022 => x"01af1fe5",
			2023 => x"040a010c",
			2024 => x"0e08fd04",
			2025 => x"ff5c1fe5",
			2026 => x"07063d04",
			2027 => x"fcda1fe5",
			2028 => x"fe4a1fe5",
			2029 => x"0901d208",
			2030 => x"06016c04",
			2031 => x"00da1fe5",
			2032 => x"fe551fe5",
			2033 => x"040a5b08",
			2034 => x"0a024904",
			2035 => x"014f1fe5",
			2036 => x"fc6c1fe5",
			2037 => x"020a2d04",
			2038 => x"019f1fe5",
			2039 => x"02e91fe5",
			2040 => x"fe6c1fe5",
			2041 => x"01010604",
			2042 => x"fe642039",
			2043 => x"0e09c124",
			2044 => x"0802fb20",
			2045 => x"0e08e104",
			2046 => x"01d42039",
			2047 => x"02095d0c",
			2048 => x"03092204",
			2049 => x"ffd22039",
			2050 => x"0a021d04",
			2051 => x"fe962039",
			2052 => x"fd152039",
			2053 => x"0901d208",
			2054 => x"0c05f304",
			2055 => x"00e22039",
			2056 => x"fda12039",
			2057 => x"0901d404",
			2058 => x"08672039",
			2059 => x"01b02039",
			2060 => x"fe0b2039",
			2061 => x"fe672039",
			2062 => x"0802fb38",
			2063 => x"06015704",
			2064 => x"fead20ad",
			2065 => x"0d07f114",
			2066 => x"0705e80c",
			2067 => x"01010f08",
			2068 => x"02095704",
			2069 => x"ffc220ad",
			2070 => x"000020ad",
			2071 => x"00b320ad",
			2072 => x"06018104",
			2073 => x"017520ad",
			2074 => x"000020ad",
			2075 => x"040adc14",
			2076 => x"0e098710",
			2077 => x"02098108",
			2078 => x"0e090704",
			2079 => x"009520ad",
			2080 => x"fec520ad",
			2081 => x"0d082204",
			2082 => x"014320ad",
			2083 => x"ffa720ad",
			2084 => x"fe8820ad",
			2085 => x"05080408",
			2086 => x"0e09e004",
			2087 => x"01b320ad",
			2088 => x"000020ad",
			2089 => x"ff1e20ad",
			2090 => x"fe7020ad",
			2091 => x"0802fb34",
			2092 => x"06015704",
			2093 => x"fec02119",
			2094 => x"0d07f114",
			2095 => x"01010604",
			2096 => x"00002119",
			2097 => x"0601810c",
			2098 => x"0c05a008",
			2099 => x"0c059f04",
			2100 => x"00882119",
			2101 => x"00002119",
			2102 => x"01682119",
			2103 => x"00002119",
			2104 => x"0c05d604",
			2105 => x"febf2119",
			2106 => x"0901d20c",
			2107 => x"0c05fa04",
			2108 => x"00002119",
			2109 => x"02095d04",
			2110 => x"00002119",
			2111 => x"feea2119",
			2112 => x"0d086d08",
			2113 => x"040ac204",
			2114 => x"000e2119",
			2115 => x"01942119",
			2116 => x"ff2c2119",
			2117 => x"fe742119",
			2118 => x"01010604",
			2119 => x"fe682195",
			2120 => x"0e08e104",
			2121 => x"01b02195",
			2122 => x"0c05f91c",
			2123 => x"0409c704",
			2124 => x"fdfa2195",
			2125 => x"0e093308",
			2126 => x"02095104",
			2127 => x"00002195",
			2128 => x"019c2195",
			2129 => x"040a7b08",
			2130 => x"0c05f704",
			2131 => x"fe682195",
			2132 => x"000d2195",
			2133 => x"0e09c104",
			2134 => x"01752195",
			2135 => x"fedb2195",
			2136 => x"07063f08",
			2137 => x"0309b004",
			2138 => x"01042195",
			2139 => x"00002195",
			2140 => x"0c05fc08",
			2141 => x"01013404",
			2142 => x"fbc32195",
			2143 => x"00002195",
			2144 => x"0e098708",
			2145 => x"0901df04",
			2146 => x"fe632195",
			2147 => x"012b2195",
			2148 => x"fe7a2195",
			2149 => x"01010604",
			2150 => x"fe6e223b",
			2151 => x"0e08e108",
			2152 => x"06015704",
			2153 => x"0000223b",
			2154 => x"0190223b",
			2155 => x"0c05d714",
			2156 => x"0d07ee0c",
			2157 => x"01012304",
			2158 => x"ff2d223b",
			2159 => x"040b1604",
			2160 => x"0102223b",
			2161 => x"0000223b",
			2162 => x"01013b04",
			2163 => x"fe53223b",
			2164 => x"0000223b",
			2165 => x"0706581c",
			2166 => x"0a02390c",
			2167 => x"02093004",
			2168 => x"ff04223b",
			2169 => x"0d080a04",
			2170 => x"010d223b",
			2171 => x"ff93223b",
			2172 => x"06018808",
			2173 => x"040a1504",
			2174 => x"0000223b",
			2175 => x"01b7223b",
			2176 => x"0d081704",
			2177 => x"0000223b",
			2178 => x"ff28223b",
			2179 => x"0c05f40c",
			2180 => x"0a023904",
			2181 => x"0000223b",
			2182 => x"06018d04",
			2183 => x"011b223b",
			2184 => x"0000223b",
			2185 => x"0802be04",
			2186 => x"0000223b",
			2187 => x"040b1c04",
			2188 => x"fde3223b",
			2189 => x"ff4e223b",
			2190 => x"0000223d",
			2191 => x"00002241",
			2192 => x"00002245",
			2193 => x"00002249",
			2194 => x"0000224d",
			2195 => x"00002251",
			2196 => x"00002255",
			2197 => x"00002259",
			2198 => x"0000225d",
			2199 => x"00002261",
			2200 => x"00002265",
			2201 => x"00002269",
			2202 => x"0000226d",
			2203 => x"00002271",
			2204 => x"00002275",
			2205 => x"00002279",
			2206 => x"0000227d",
			2207 => x"00002281",
			2208 => x"00002285",
			2209 => x"00002289",
			2210 => x"0000228d",
			2211 => x"00002291",
			2212 => x"00002295",
			2213 => x"00002299",
			2214 => x"0000229d",
			2215 => x"000022a1",
			2216 => x"000022a5",
			2217 => x"0e093304",
			2218 => x"000022b1",
			2219 => x"fffc22b1",
			2220 => x"0802be04",
			2221 => x"000022bd",
			2222 => x"fff522bd",
			2223 => x"0901f004",
			2224 => x"fffd22c9",
			2225 => x"000022c9",
			2226 => x"0e08e108",
			2227 => x"0e081604",
			2228 => x"000022dd",
			2229 => x"002822dd",
			2230 => x"fffb22dd",
			2231 => x"01012408",
			2232 => x"0901d904",
			2233 => x"ffe422f1",
			2234 => x"000022f1",
			2235 => x"000022f1",
			2236 => x"01011104",
			2237 => x"00002305",
			2238 => x"09020804",
			2239 => x"00192305",
			2240 => x"00002305",
			2241 => x"0e08e10c",
			2242 => x"0e081604",
			2243 => x"00002321",
			2244 => x"03093704",
			2245 => x"00332321",
			2246 => x"00002321",
			2247 => x"fff32321",
			2248 => x"0101370c",
			2249 => x"0c060f08",
			2250 => x"0802a504",
			2251 => x"0000233d",
			2252 => x"ffcc233d",
			2253 => x"0000233d",
			2254 => x"0000233d",
			2255 => x"0e09330c",
			2256 => x"0f091f04",
			2257 => x"00002361",
			2258 => x"0f09a304",
			2259 => x"00052361",
			2260 => x"00002361",
			2261 => x"0f099504",
			2262 => x"00002361",
			2263 => x"fffb2361",
			2264 => x"0e08e10c",
			2265 => x"09019c04",
			2266 => x"0000238d",
			2267 => x"00030204",
			2268 => x"0000238d",
			2269 => x"0031238d",
			2270 => x"01013f08",
			2271 => x"0c059f04",
			2272 => x"0000238d",
			2273 => x"ffbb238d",
			2274 => x"0000238d",
			2275 => x"01011704",
			2276 => x"000023b1",
			2277 => x"0902080c",
			2278 => x"0802fb08",
			2279 => x"0802aa04",
			2280 => x"000023b1",
			2281 => x"002a23b1",
			2282 => x"000023b1",
			2283 => x"000023b1",
			2284 => x"0802e610",
			2285 => x"0d08220c",
			2286 => x"08026f04",
			2287 => x"000023d5",
			2288 => x"0d071604",
			2289 => x"000023d5",
			2290 => x"003123d5",
			2291 => x"000023d5",
			2292 => x"000023d5",
			2293 => x"0901f010",
			2294 => x"0e08e104",
			2295 => x"000023f9",
			2296 => x"020a6308",
			2297 => x"03092204",
			2298 => x"000023f9",
			2299 => x"ffdd23f9",
			2300 => x"000023f9",
			2301 => x"000023f9",
			2302 => x"0e08e110",
			2303 => x"0e081604",
			2304 => x"00002425",
			2305 => x"02089004",
			2306 => x"00002425",
			2307 => x"020a1004",
			2308 => x"00312425",
			2309 => x"00002425",
			2310 => x"040a5b04",
			2311 => x"ffc52425",
			2312 => x"00002425",
			2313 => x"0901d908",
			2314 => x"0b06ae04",
			2315 => x"00002459",
			2316 => x"ff962459",
			2317 => x"040a2804",
			2318 => x"00002459",
			2319 => x"0f0a190c",
			2320 => x"0c061708",
			2321 => x"0a026204",
			2322 => x"007b2459",
			2323 => x"00002459",
			2324 => x"00002459",
			2325 => x"00002459",
			2326 => x"0e08e104",
			2327 => x"00002485",
			2328 => x"0901f010",
			2329 => x"0c060f0c",
			2330 => x"0c059f04",
			2331 => x"00002485",
			2332 => x"01013704",
			2333 => x"ffc02485",
			2334 => x"00002485",
			2335 => x"00002485",
			2336 => x"00002485",
			2337 => x"0209a414",
			2338 => x"0e08e108",
			2339 => x"01011104",
			2340 => x"ffb724d1",
			2341 => x"006524d1",
			2342 => x"040a2808",
			2343 => x"0c061704",
			2344 => x"ff2d24d1",
			2345 => x"000024d1",
			2346 => x"000024d1",
			2347 => x"0e09870c",
			2348 => x"0003ea08",
			2349 => x"01010604",
			2350 => x"000024d1",
			2351 => x"00be24d1",
			2352 => x"000024d1",
			2353 => x"01013904",
			2354 => x"ffc324d1",
			2355 => x"000024d1",
			2356 => x"02097010",
			2357 => x"0c06140c",
			2358 => x"06017408",
			2359 => x"0e08cb04",
			2360 => x"0000251d",
			2361 => x"ffb7251d",
			2362 => x"0000251d",
			2363 => x"0000251d",
			2364 => x"0e093310",
			2365 => x"06016004",
			2366 => x"0000251d",
			2367 => x"0c061308",
			2368 => x"0a026d04",
			2369 => x"007e251d",
			2370 => x"0000251d",
			2371 => x"0000251d",
			2372 => x"040a7b04",
			2373 => x"ffc8251d",
			2374 => x"0000251d",
			2375 => x"0101170c",
			2376 => x"0901c308",
			2377 => x"04091d04",
			2378 => x"00002561",
			2379 => x"ffdc2561",
			2380 => x"00002561",
			2381 => x"0d086d14",
			2382 => x"040a3a04",
			2383 => x"00002561",
			2384 => x"0e09c10c",
			2385 => x"06018908",
			2386 => x"00034b04",
			2387 => x"00002561",
			2388 => x"009a2561",
			2389 => x"00002561",
			2390 => x"00002561",
			2391 => x"00002561",
			2392 => x"0c05b80c",
			2393 => x"0802a504",
			2394 => x"000025ad",
			2395 => x"01012104",
			2396 => x"ffd925ad",
			2397 => x"000025ad",
			2398 => x"040a5b08",
			2399 => x"0802be04",
			2400 => x"000025ad",
			2401 => x"ffd325ad",
			2402 => x"06018610",
			2403 => x"0802fb0c",
			2404 => x"020a6b08",
			2405 => x"0c063a04",
			2406 => x"00bb25ad",
			2407 => x"000025ad",
			2408 => x"000025ad",
			2409 => x"000025ad",
			2410 => x"000025ad",
			2411 => x"0c05d704",
			2412 => x"000025e1",
			2413 => x"0d083814",
			2414 => x"0c061310",
			2415 => x"0e09c10c",
			2416 => x"01011104",
			2417 => x"000025e1",
			2418 => x"0d083104",
			2419 => x"008725e1",
			2420 => x"000025e1",
			2421 => x"000025e1",
			2422 => x"000025e1",
			2423 => x"000025e1",
			2424 => x"01012410",
			2425 => x"0c05b80c",
			2426 => x"07061608",
			2427 => x"0409c704",
			2428 => x"00002635",
			2429 => x"ffb52635",
			2430 => x"00002635",
			2431 => x"00002635",
			2432 => x"040a3a08",
			2433 => x"01012804",
			2434 => x"00002635",
			2435 => x"fffb2635",
			2436 => x"0f0a5a10",
			2437 => x"0601860c",
			2438 => x"01014b08",
			2439 => x"0c061704",
			2440 => x"009d2635",
			2441 => x"00002635",
			2442 => x"00002635",
			2443 => x"00002635",
			2444 => x"00002635",
			2445 => x"01010b08",
			2446 => x"01010604",
			2447 => x"c8fc2691",
			2448 => x"cbf82691",
			2449 => x"03096814",
			2450 => x"0b06cb0c",
			2451 => x"08028704",
			2452 => x"e4a02691",
			2453 => x"01013c04",
			2454 => x"f6e42691",
			2455 => x"e6352691",
			2456 => x"00033504",
			2457 => x"c9462691",
			2458 => x"e7f92691",
			2459 => x"0e098708",
			2460 => x"040a5b04",
			2461 => x"c9092691",
			2462 => x"f40c2691",
			2463 => x"0e09c108",
			2464 => x"01013904",
			2465 => x"c9102691",
			2466 => x"d4e52691",
			2467 => x"c8fc2691",
			2468 => x"0209be20",
			2469 => x"0a024c18",
			2470 => x"0e092410",
			2471 => x"0901f20c",
			2472 => x"01011304",
			2473 => x"000026f5",
			2474 => x"0507bc04",
			2475 => x"00b926f5",
			2476 => x"000026f5",
			2477 => x"000026f5",
			2478 => x"01013a04",
			2479 => x"ffde26f5",
			2480 => x"000026f5",
			2481 => x"0209b704",
			2482 => x"fec326f5",
			2483 => x"000026f5",
			2484 => x"0309c00c",
			2485 => x"06018808",
			2486 => x"01010604",
			2487 => x"000026f5",
			2488 => x"011326f5",
			2489 => x"000026f5",
			2490 => x"01013904",
			2491 => x"ff9826f5",
			2492 => x"000026f5",
			2493 => x"0c05d70c",
			2494 => x"0802be04",
			2495 => x"00002759",
			2496 => x"0901ec04",
			2497 => x"fecc2759",
			2498 => x"00002759",
			2499 => x"07062c10",
			2500 => x"0409c704",
			2501 => x"00002759",
			2502 => x"0e09e008",
			2503 => x"01011104",
			2504 => x"00002759",
			2505 => x"00e42759",
			2506 => x"00002759",
			2507 => x"0c05f90c",
			2508 => x"0d081708",
			2509 => x"01011304",
			2510 => x"00002759",
			2511 => x"00652759",
			2512 => x"00002759",
			2513 => x"0802c304",
			2514 => x"00002759",
			2515 => x"040b1c04",
			2516 => x"ff1e2759",
			2517 => x"00002759",
			2518 => x"0c05b80c",
			2519 => x"01012108",
			2520 => x"00032c04",
			2521 => x"000027bd",
			2522 => x"ff8227bd",
			2523 => x"000027bd",
			2524 => x"07062a0c",
			2525 => x"06018908",
			2526 => x"01010604",
			2527 => x"000027bd",
			2528 => x"00b527bd",
			2529 => x"000027bd",
			2530 => x"0901f010",
			2531 => x"0e08fd04",
			2532 => x"000027bd",
			2533 => x"06016c04",
			2534 => x"000027bd",
			2535 => x"01013804",
			2536 => x"ff4327bd",
			2537 => x"000027bd",
			2538 => x"0c05f808",
			2539 => x"0e09c104",
			2540 => x"007827bd",
			2541 => x"000027bd",
			2542 => x"000027bd",
			2543 => x"01012420",
			2544 => x"0802c318",
			2545 => x"08027908",
			2546 => x"0a020804",
			2547 => x"ff802831",
			2548 => x"00002831",
			2549 => x"0e09330c",
			2550 => x"0901a904",
			2551 => x"00002831",
			2552 => x"0507c704",
			2553 => x"008e2831",
			2554 => x"00002831",
			2555 => x"00002831",
			2556 => x"01012104",
			2557 => x"fef12831",
			2558 => x"00002831",
			2559 => x"0e09a214",
			2560 => x"0a02390c",
			2561 => x"03094008",
			2562 => x"01013604",
			2563 => x"00762831",
			2564 => x"00002831",
			2565 => x"ff8b2831",
			2566 => x"0309b004",
			2567 => x"012a2831",
			2568 => x"00002831",
			2569 => x"0507b804",
			2570 => x"00002831",
			2571 => x"ff9f2831",
			2572 => x"0c05b810",
			2573 => x"0101210c",
			2574 => x"08029e04",
			2575 => x"0000289d",
			2576 => x"07061504",
			2577 => x"ff7f289d",
			2578 => x"0000289d",
			2579 => x"0000289d",
			2580 => x"07062a0c",
			2581 => x"0901f608",
			2582 => x"01010604",
			2583 => x"0000289d",
			2584 => x"00b7289d",
			2585 => x"0000289d",
			2586 => x"0f099510",
			2587 => x"0a022304",
			2588 => x"0000289d",
			2589 => x"0802c308",
			2590 => x"02093004",
			2591 => x"0000289d",
			2592 => x"007f289d",
			2593 => x"0000289d",
			2594 => x"01013408",
			2595 => x"0e092404",
			2596 => x"0000289d",
			2597 => x"ff7c289d",
			2598 => x"0000289d",
			2599 => x"0c05d71c",
			2600 => x"0209a410",
			2601 => x"0b06cf0c",
			2602 => x"0d081808",
			2603 => x"07062e04",
			2604 => x"fedf2919",
			2605 => x"00002919",
			2606 => x"00002919",
			2607 => x"00002919",
			2608 => x"0e097708",
			2609 => x"0d073004",
			2610 => x"00002919",
			2611 => x"00112919",
			2612 => x"00002919",
			2613 => x"0d081714",
			2614 => x"0c05f910",
			2615 => x"02093004",
			2616 => x"00002919",
			2617 => x"0e09c108",
			2618 => x"06016004",
			2619 => x"00002919",
			2620 => x"00d62919",
			2621 => x"00002919",
			2622 => x"00002919",
			2623 => x"040abb0c",
			2624 => x"0c05d904",
			2625 => x"00002919",
			2626 => x"0b06ae04",
			2627 => x"00002919",
			2628 => x"ff722919",
			2629 => x"00002919",
			2630 => x"0901bc04",
			2631 => x"00002955",
			2632 => x"05080418",
			2633 => x"00031a04",
			2634 => x"00002955",
			2635 => x"06018810",
			2636 => x"0e09c10c",
			2637 => x"0705ff04",
			2638 => x"00002955",
			2639 => x"0a022b04",
			2640 => x"00002955",
			2641 => x"00662955",
			2642 => x"00002955",
			2643 => x"00002955",
			2644 => x"00002955",
			2645 => x"02093004",
			2646 => x"00002991",
			2647 => x"0b06cf18",
			2648 => x"0802aa04",
			2649 => x"00002991",
			2650 => x"07065a10",
			2651 => x"040a0104",
			2652 => x"00002991",
			2653 => x"0802fb08",
			2654 => x"0e09c104",
			2655 => x"009b2991",
			2656 => x"00002991",
			2657 => x"00002991",
			2658 => x"00002991",
			2659 => x"00002991",
			2660 => x"0901a90c",
			2661 => x"09019c04",
			2662 => x"fe5a29fd",
			2663 => x"0901a104",
			2664 => x"fff629fd",
			2665 => x"fe8e29fd",
			2666 => x"0d082218",
			2667 => x"0e09c114",
			2668 => x"0f08e604",
			2669 => x"05df29fd",
			2670 => x"00031a04",
			2671 => x"016629fd",
			2672 => x"0f0a0308",
			2673 => x"0901fe04",
			2674 => x"041529fd",
			2675 => x"024329fd",
			2676 => x"06ab29fd",
			2677 => x"fe7b29fd",
			2678 => x"0e098708",
			2679 => x"0901e604",
			2680 => x"fe4729fd",
			2681 => x"039629fd",
			2682 => x"0e09c108",
			2683 => x"0c05f304",
			2684 => x"015d29fd",
			2685 => x"fe7929fd",
			2686 => x"fe5b29fd",
			2687 => x"0901a904",
			2688 => x"fe672a51",
			2689 => x"0e096214",
			2690 => x"0e08e104",
			2691 => x"01aa2a51",
			2692 => x"0409db04",
			2693 => x"fdaa2a51",
			2694 => x"0901d204",
			2695 => x"fea12a51",
			2696 => x"06018104",
			2697 => x"01af2a51",
			2698 => x"007c2a51",
			2699 => x"0c05f810",
			2700 => x"040a8804",
			2701 => x"fe562a51",
			2702 => x"0e09c108",
			2703 => x"020a1004",
			2704 => x"00892a51",
			2705 => x"020c2a51",
			2706 => x"febc2a51",
			2707 => x"fe712a51",
			2708 => x"0c05d720",
			2709 => x"0209a410",
			2710 => x"0b06cf0c",
			2711 => x"0d081808",
			2712 => x"07062e04",
			2713 => x"feb42ae5",
			2714 => x"00002ae5",
			2715 => x"00002ae5",
			2716 => x"00002ae5",
			2717 => x"0e09770c",
			2718 => x"0b062a04",
			2719 => x"00002ae5",
			2720 => x"020a1004",
			2721 => x"00262ae5",
			2722 => x"00002ae5",
			2723 => x"00002ae5",
			2724 => x"0901d90c",
			2725 => x"0c05f904",
			2726 => x"00002ae5",
			2727 => x"0c061404",
			2728 => x"ff542ae5",
			2729 => x"00002ae5",
			2730 => x"0d08170c",
			2731 => x"02093004",
			2732 => x"00002ae5",
			2733 => x"0e09c104",
			2734 => x"00fe2ae5",
			2735 => x"00002ae5",
			2736 => x"040abb0c",
			2737 => x"01012a04",
			2738 => x"00002ae5",
			2739 => x"07063f04",
			2740 => x"00002ae5",
			2741 => x"ffbb2ae5",
			2742 => x"0e09e004",
			2743 => x"000b2ae5",
			2744 => x"00002ae5",
			2745 => x"01010604",
			2746 => x"fe6d2b39",
			2747 => x"0e08e108",
			2748 => x"0b06bb04",
			2749 => x"01942b39",
			2750 => x"00002b39",
			2751 => x"040a150c",
			2752 => x"0409c704",
			2753 => x"fe3c2b39",
			2754 => x"03092e04",
			2755 => x"00672b39",
			2756 => x"febc2b39",
			2757 => x"0e09c110",
			2758 => x"01011f04",
			2759 => x"fee12b39",
			2760 => x"040a8808",
			2761 => x"0e096204",
			2762 => x"014a2b39",
			2763 => x"fe992b39",
			2764 => x"01ce2b39",
			2765 => x"fe9f2b39",
			2766 => x"01010604",
			2767 => x"fe5d2b95",
			2768 => x"0d082218",
			2769 => x"0802f814",
			2770 => x"020a2d10",
			2771 => x"0c06130c",
			2772 => x"020a1008",
			2773 => x"0309a304",
			2774 => x"02db2b95",
			2775 => x"01342b95",
			2776 => x"042a2b95",
			2777 => x"01342b95",
			2778 => x"075a2b95",
			2779 => x"fe362b95",
			2780 => x"0507bc08",
			2781 => x"0003c804",
			2782 => x"03e42b95",
			2783 => x"ff302b95",
			2784 => x"0e096208",
			2785 => x"01012304",
			2786 => x"fe4b2b95",
			2787 => x"02a82b95",
			2788 => x"fe5e2b95",
			2789 => x"0802fb2c",
			2790 => x"040adc1c",
			2791 => x"0e098718",
			2792 => x"01011108",
			2793 => x"0901b804",
			2794 => x"feb72bf1",
			2795 => x"00002bf1",
			2796 => x"040a3a0c",
			2797 => x"0507a004",
			2798 => x"011d2bf1",
			2799 => x"0e08e104",
			2800 => x"00ae2bf1",
			2801 => x"ff352bf1",
			2802 => x"014f2bf1",
			2803 => x"fe922bf1",
			2804 => x"0508040c",
			2805 => x"01010604",
			2806 => x"00002bf1",
			2807 => x"0e09e004",
			2808 => x"01b32bf1",
			2809 => x"00002bf1",
			2810 => x"ff2f2bf1",
			2811 => x"fe722bf1",
			2812 => x"0802f838",
			2813 => x"0e08fd18",
			2814 => x"0209130c",
			2815 => x"00033508",
			2816 => x"01011104",
			2817 => x"ffe82c65",
			2818 => x"00292c65",
			2819 => x"ff2a2c65",
			2820 => x"03092e08",
			2821 => x"01010604",
			2822 => x"00002c65",
			2823 => x"016a2c65",
			2824 => x"00002c65",
			2825 => x"01013410",
			2826 => x"0d07e404",
			2827 => x"00002c65",
			2828 => x"07065b08",
			2829 => x"06016c04",
			2830 => x"00002c65",
			2831 => x"fe912c65",
			2832 => x"00002c65",
			2833 => x"0d081708",
			2834 => x"02099504",
			2835 => x"00002c65",
			2836 => x"01202c65",
			2837 => x"0e098704",
			2838 => x"00002c65",
			2839 => x"ff392c65",
			2840 => x"fe7d2c65",
			2841 => x"01011108",
			2842 => x"0901b804",
			2843 => x"fe812ce9",
			2844 => x"00002ce9",
			2845 => x"0f09b11c",
			2846 => x"0409db0c",
			2847 => x"0308f704",
			2848 => x"00b42ce9",
			2849 => x"0c05f804",
			2850 => x"fec22ce9",
			2851 => x"00002ce9",
			2852 => x"0c061308",
			2853 => x"03097804",
			2854 => x"01622ce9",
			2855 => x"00002ce9",
			2856 => x"0901db04",
			2857 => x"ffb52ce9",
			2858 => x"00092ce9",
			2859 => x"0901f008",
			2860 => x"0b069c04",
			2861 => x"00002ce9",
			2862 => x"fe862ce9",
			2863 => x"0d081708",
			2864 => x"0003a704",
			2865 => x"01192ce9",
			2866 => x"00002ce9",
			2867 => x"0901f608",
			2868 => x"0b06f004",
			2869 => x"00002ce9",
			2870 => x"002e2ce9",
			2871 => x"0b06bb04",
			2872 => x"00002ce9",
			2873 => x"ff112ce9",
			2874 => x"0901a904",
			2875 => x"fe682d55",
			2876 => x"0e096218",
			2877 => x"0e08e104",
			2878 => x"01a32d55",
			2879 => x"0409db04",
			2880 => x"fdf22d55",
			2881 => x"0901d204",
			2882 => x"fecd2d55",
			2883 => x"06018108",
			2884 => x"0901d904",
			2885 => x"003e2d55",
			2886 => x"01b12d55",
			2887 => x"005b2d55",
			2888 => x"0c05f810",
			2889 => x"040a8804",
			2890 => x"fe6a2d55",
			2891 => x"0e09c108",
			2892 => x"020a1004",
			2893 => x"00612d55",
			2894 => x"01d92d55",
			2895 => x"feda2d55",
			2896 => x"0f09e108",
			2897 => x"06017804",
			2898 => x"ffed2d55",
			2899 => x"00002d55",
			2900 => x"fe6f2d55",
			2901 => x"0802fb30",
			2902 => x"040adc20",
			2903 => x"0e09771c",
			2904 => x"02098114",
			2905 => x"0e090710",
			2906 => x"06015708",
			2907 => x"02090c04",
			2908 => x"ff312db9",
			2909 => x"00002db9",
			2910 => x"0705e804",
			2911 => x"00002db9",
			2912 => x"00d42db9",
			2913 => x"fed32db9",
			2914 => x"0507ca04",
			2915 => x"013b2db9",
			2916 => x"00002db9",
			2917 => x"fee32db9",
			2918 => x"0d086d0c",
			2919 => x"06015c04",
			2920 => x"00002db9",
			2921 => x"0e09e004",
			2922 => x"01ba2db9",
			2923 => x"00002db9",
			2924 => x"ffdf2db9",
			2925 => x"fe8c2db9",
			2926 => x"0802fb38",
			2927 => x"040adc28",
			2928 => x"0802c31c",
			2929 => x"0d07ee08",
			2930 => x"0901a904",
			2931 => x"00002e2d",
			2932 => x"00b82e2d",
			2933 => x"0409db08",
			2934 => x"0e08c304",
			2935 => x"00002e2d",
			2936 => x"ff372e2d",
			2937 => x"03096804",
			2938 => x"00b72e2d",
			2939 => x"0a024504",
			2940 => x"ffa52e2d",
			2941 => x"00002e2d",
			2942 => x"0901ee08",
			2943 => x"0507d904",
			2944 => x"fec62e2d",
			2945 => x"00002e2d",
			2946 => x"00002e2d",
			2947 => x"0508040c",
			2948 => x"09019c04",
			2949 => x"00002e2d",
			2950 => x"0e09e004",
			2951 => x"01362e2d",
			2952 => x"00002e2d",
			2953 => x"00002e2d",
			2954 => x"fecc2e2d",
			2955 => x"0901a904",
			2956 => x"fe612e81",
			2957 => x"0e09c124",
			2958 => x"0d08311c",
			2959 => x"020a2d18",
			2960 => x"0d082210",
			2961 => x"03091a08",
			2962 => x"08028704",
			2963 => x"03062e81",
			2964 => x"02332e81",
			2965 => x"040a0104",
			2966 => x"fd642e81",
			2967 => x"021d2e81",
			2968 => x"01013204",
			2969 => x"fe6a2e81",
			2970 => x"014d2e81",
			2971 => x"04702e81",
			2972 => x"0f0a0304",
			2973 => x"fe6e2e81",
			2974 => x"026b2e81",
			2975 => x"fe622e81",
			2976 => x"01010604",
			2977 => x"feaf2efd",
			2978 => x"040a882c",
			2979 => x"0f09b120",
			2980 => x"0409db0c",
			2981 => x"0308f704",
			2982 => x"004b2efd",
			2983 => x"07065a04",
			2984 => x"ff352efd",
			2985 => x"00002efd",
			2986 => x"0c060f08",
			2987 => x"03099604",
			2988 => x"01092efd",
			2989 => x"00002efd",
			2990 => x"00035b08",
			2991 => x"03097804",
			2992 => x"00382efd",
			2993 => x"00002efd",
			2994 => x"ff9e2efd",
			2995 => x"040a7b08",
			2996 => x"09020204",
			2997 => x"fede2efd",
			2998 => x"00002efd",
			2999 => x"00002efd",
			3000 => x"0309d808",
			3001 => x"06018d04",
			3002 => x"01642efd",
			3003 => x"00002efd",
			3004 => x"0802d504",
			3005 => x"00002efd",
			3006 => x"ff852efd",
			3007 => x"01010f08",
			3008 => x"0901b804",
			3009 => x"fe902f89",
			3010 => x"00002f89",
			3011 => x"07062a10",
			3012 => x"0309c00c",
			3013 => x"0901f608",
			3014 => x"0c057204",
			3015 => x"00002f89",
			3016 => x"01a32f89",
			3017 => x"00002f89",
			3018 => x"00002f89",
			3019 => x"01012e10",
			3020 => x"0e08e104",
			3021 => x"004b2f89",
			3022 => x"0901df08",
			3023 => x"07066f04",
			3024 => x"feef2f89",
			3025 => x"00002f89",
			3026 => x"00002f89",
			3027 => x"0d08170c",
			3028 => x"02096004",
			3029 => x"00002f89",
			3030 => x"0e09c104",
			3031 => x"01272f89",
			3032 => x"00002f89",
			3033 => x"0c05f80c",
			3034 => x"0901f004",
			3035 => x"00002f89",
			3036 => x"06018504",
			3037 => x"00ae2f89",
			3038 => x"00002f89",
			3039 => x"0901e804",
			3040 => x"00002f89",
			3041 => x"ff392f89",
			3042 => x"0802fb3c",
			3043 => x"040a8828",
			3044 => x"0e095120",
			3045 => x"040a1514",
			3046 => x"0e08e10c",
			3047 => x"06015304",
			3048 => x"00003005",
			3049 => x"0d077004",
			3050 => x"00003005",
			3051 => x"00b03005",
			3052 => x"0f097d04",
			3053 => x"fefb3005",
			3054 => x"00003005",
			3055 => x"01011304",
			3056 => x"00003005",
			3057 => x"0802aa04",
			3058 => x"00003005",
			3059 => x"01263005",
			3060 => x"01013c04",
			3061 => x"fe9b3005",
			3062 => x"00003005",
			3063 => x"0d086d10",
			3064 => x"01010604",
			3065 => x"00003005",
			3066 => x"06018608",
			3067 => x"0e09c104",
			3068 => x"01aa3005",
			3069 => x"00003005",
			3070 => x"00003005",
			3071 => x"ffc93005",
			3072 => x"fe933005",
			3073 => x"01010604",
			3074 => x"fe6b3091",
			3075 => x"07062c18",
			3076 => x"040a280c",
			3077 => x"03092204",
			3078 => x"01763091",
			3079 => x"040a0104",
			3080 => x"fe793091",
			3081 => x"00003091",
			3082 => x"0e09c108",
			3083 => x"040b7d04",
			3084 => x"01893091",
			3085 => x"03063091",
			3086 => x"ff973091",
			3087 => x"0e095114",
			3088 => x"0a022b08",
			3089 => x"03091a04",
			3090 => x"00473091",
			3091 => x"fe773091",
			3092 => x"0901c804",
			3093 => x"ff173091",
			3094 => x"00034604",
			3095 => x"00033091",
			3096 => x"01933091",
			3097 => x"03098704",
			3098 => x"fdcb3091",
			3099 => x"0507e410",
			3100 => x"07064008",
			3101 => x"0309d804",
			3102 => x"00843091",
			3103 => x"00003091",
			3104 => x"07065804",
			3105 => x"ff3f3091",
			3106 => x"00003091",
			3107 => x"fe993091",
			3108 => x"01010604",
			3109 => x"fe6630ed",
			3110 => x"0e09c128",
			3111 => x"03091a04",
			3112 => x"01b430ed",
			3113 => x"040a010c",
			3114 => x"0f095608",
			3115 => x"0e08fd04",
			3116 => x"000d30ed",
			3117 => x"fec430ed",
			3118 => x"fd9030ed",
			3119 => x"01011f08",
			3120 => x"0e096204",
			3121 => x"ff8d30ed",
			3122 => x"fe1e30ed",
			3123 => x"040a5b08",
			3124 => x"0a024904",
			3125 => x"00e530ed",
			3126 => x"fc9b30ed",
			3127 => x"020a2d04",
			3128 => x"01a930ed",
			3129 => x"02b330ed",
			3130 => x"fe6d30ed",
			3131 => x"0901a904",
			3132 => x"fe623159",
			3133 => x"0e09c130",
			3134 => x"0c06131c",
			3135 => x"020a2d18",
			3136 => x"0d082210",
			3137 => x"0e095108",
			3138 => x"040a0104",
			3139 => x"01aa3159",
			3140 => x"02053159",
			3141 => x"040a5b04",
			3142 => x"fd9f3159",
			3143 => x"01963159",
			3144 => x"040a5b04",
			3145 => x"fe733159",
			3146 => x"00c63159",
			3147 => x"044c3159",
			3148 => x"0c061408",
			3149 => x"0901d404",
			3150 => x"fca93159",
			3151 => x"00723159",
			3152 => x"0d083004",
			3153 => x"02303159",
			3154 => x"01012e04",
			3155 => x"fe793159",
			3156 => x"00593159",
			3157 => x"fe643159",
			3158 => x"01010604",
			3159 => x"fe6a31f5",
			3160 => x"07062c1c",
			3161 => x"040b9d14",
			3162 => x"03092204",
			3163 => x"019331f5",
			3164 => x"040a0104",
			3165 => x"fe6131f5",
			3166 => x"0e09c108",
			3167 => x"040a2804",
			3168 => x"000031f5",
			3169 => x"017a31f5",
			3170 => x"ffc831f5",
			3171 => x"0f0ac904",
			3172 => x"03a131f5",
			3173 => x"000031f5",
			3174 => x"0e095110",
			3175 => x"0a022b08",
			3176 => x"03091a04",
			3177 => x"005431f5",
			3178 => x"fe6b31f5",
			3179 => x"01012104",
			3180 => x"ffdd31f5",
			3181 => x"018131f5",
			3182 => x"0c05f810",
			3183 => x"07064008",
			3184 => x"0309d804",
			3185 => x"00a531f5",
			3186 => x"000031f5",
			3187 => x"0c05f704",
			3188 => x"fef031f5",
			3189 => x"000031f5",
			3190 => x"0b06bd04",
			3191 => x"fdaa31f5",
			3192 => x"0309a308",
			3193 => x"0507e404",
			3194 => x"003c31f5",
			3195 => x"000031f5",
			3196 => x"fe9631f5",
			3197 => x"0802f83c",
			3198 => x"06015704",
			3199 => x"fea73271",
			3200 => x"0e092418",
			3201 => x"0e08e108",
			3202 => x"0e081604",
			3203 => x"00003271",
			3204 => x"01ab3271",
			3205 => x"0209700c",
			3206 => x"03092208",
			3207 => x"0a023304",
			3208 => x"012b3271",
			3209 => x"00003271",
			3210 => x"feba3271",
			3211 => x"01943271",
			3212 => x"040a5b10",
			3213 => x"0a024c0c",
			3214 => x"0a023904",
			3215 => x"fe523271",
			3216 => x"0802be04",
			3217 => x"009b3271",
			3218 => x"ff173271",
			3219 => x"fd0f3271",
			3220 => x"0e09c10c",
			3221 => x"040a8808",
			3222 => x"03098704",
			3223 => x"014e3271",
			3224 => x"fef53271",
			3225 => x"017f3271",
			3226 => x"fe8e3271",
			3227 => x"fe693271",
			3228 => x"01010604",
			3229 => x"fed532fd",
			3230 => x"0e08e108",
			3231 => x"0f099504",
			3232 => x"00ed32fd",
			3233 => x"000032fd",
			3234 => x"0101240c",
			3235 => x"0d07ca04",
			3236 => x"000032fd",
			3237 => x"0901d904",
			3238 => x"fef232fd",
			3239 => x"000032fd",
			3240 => x"07064318",
			3241 => x"0c05d70c",
			3242 => x"03094004",
			3243 => x"000032fd",
			3244 => x"0d07ee04",
			3245 => x"000032fd",
			3246 => x"ffbb32fd",
			3247 => x"06018808",
			3248 => x"0309c004",
			3249 => x"010232fd",
			3250 => x"000032fd",
			3251 => x"000032fd",
			3252 => x"07065b0c",
			3253 => x"0c05dc04",
			3254 => x"000032fd",
			3255 => x"0b06f004",
			3256 => x"ff0432fd",
			3257 => x"000032fd",
			3258 => x"0f0a1908",
			3259 => x"07067004",
			3260 => x"003b32fd",
			3261 => x"000032fd",
			3262 => x"000032fd",
			3263 => x"01010604",
			3264 => x"fe7033b3",
			3265 => x"0e08e108",
			3266 => x"0b06bb04",
			3267 => x"018333b3",
			3268 => x"000033b3",
			3269 => x"0c05d71c",
			3270 => x"05079c0c",
			3271 => x"01011f04",
			3272 => x"ff9733b3",
			3273 => x"08030804",
			3274 => x"00d433b3",
			3275 => x"000033b3",
			3276 => x"01012e08",
			3277 => x"0d081804",
			3278 => x"fe5633b3",
			3279 => x"000033b3",
			3280 => x"0901f004",
			3281 => x"000033b3",
			3282 => x"ffb233b3",
			3283 => x"07065820",
			3284 => x"0a023910",
			3285 => x"0d080a08",
			3286 => x"07062904",
			3287 => x"000033b3",
			3288 => x"00c233b3",
			3289 => x"0b06ce04",
			3290 => x"ff5033b3",
			3291 => x"000033b3",
			3292 => x"0c061308",
			3293 => x"0e09a204",
			3294 => x"019533b3",
			3295 => x"000033b3",
			3296 => x"0c061504",
			3297 => x"ff6e33b3",
			3298 => x"000033b3",
			3299 => x"0c05f40c",
			3300 => x"0a023904",
			3301 => x"000033b3",
			3302 => x"0802e804",
			3303 => x"010033b3",
			3304 => x"000033b3",
			3305 => x"0802be04",
			3306 => x"000033b3",
			3307 => x"fe7a33b3",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1096, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(2190, initial_addr_3'length));
	end generate gen_rom_11;

	gen_rom_12: if SELECT_ROM = 12 generate
		bank <= (
			0 => x"00000005",
			1 => x"00000009",
			2 => x"0000000d",
			3 => x"00000011",
			4 => x"00000015",
			5 => x"00000019",
			6 => x"0000001d",
			7 => x"00000021",
			8 => x"00000025",
			9 => x"00000029",
			10 => x"0000002d",
			11 => x"00000031",
			12 => x"00000035",
			13 => x"00000039",
			14 => x"0000003d",
			15 => x"00000041",
			16 => x"00000045",
			17 => x"00000049",
			18 => x"0000004d",
			19 => x"00000051",
			20 => x"00000055",
			21 => x"00000059",
			22 => x"0000005d",
			23 => x"00000061",
			24 => x"00000065",
			25 => x"00000069",
			26 => x"0000006d",
			27 => x"00000071",
			28 => x"00000075",
			29 => x"040f0204",
			30 => x"fffa0081",
			31 => x"00000081",
			32 => x"040d5504",
			33 => x"fffb008d",
			34 => x"0000008d",
			35 => x"0410bb04",
			36 => x"ffe70099",
			37 => x"00000099",
			38 => x"040fc604",
			39 => x"ffec00a5",
			40 => x"000000a5",
			41 => x"0410bb04",
			42 => x"ffe200b1",
			43 => x"000000b1",
			44 => x"0100ca04",
			45 => x"ffed00bd",
			46 => x"000000bd",
			47 => x"040fc604",
			48 => x"fff800c9",
			49 => x"000000c9",
			50 => x"040c4404",
			51 => x"fff000dd",
			52 => x"04120c04",
			53 => x"000500dd",
			54 => x"000000dd",
			55 => x"04112a08",
			56 => x"09015804",
			57 => x"ffae00f1",
			58 => x"000000f1",
			59 => x"000000f1",
			60 => x"0209ce04",
			61 => x"fff60105",
			62 => x"020a2d04",
			63 => x"000b0105",
			64 => x"00000105",
			65 => x"0209c104",
			66 => x"00000119",
			67 => x"020a2d04",
			68 => x"00350119",
			69 => x"00000119",
			70 => x"0209ce04",
			71 => x"ffef012d",
			72 => x"020a6b04",
			73 => x"0036012d",
			74 => x"0000012d",
			75 => x"0410bb08",
			76 => x"09015804",
			77 => x"ffd60141",
			78 => x"00000141",
			79 => x"00000141",
			80 => x"0100dc08",
			81 => x"020a0604",
			82 => x"ffda0155",
			83 => x"00000155",
			84 => x"00000155",
			85 => x"0209c10c",
			86 => x"06017408",
			87 => x"0100f304",
			88 => x"ffb10171",
			89 => x"00000171",
			90 => x"00000171",
			91 => x"00000171",
			92 => x"0e073b0c",
			93 => x"040d1b04",
			94 => x"0000018d",
			95 => x"04120c04",
			96 => x"0011018d",
			97 => x"0000018d",
			98 => x"fffd018d",
			99 => x"040cbf04",
			100 => x"fff601a9",
			101 => x"0209b104",
			102 => x"000001a9",
			103 => x"020a6b04",
			104 => x"001401a9",
			105 => x"000001a9",
			106 => x"0100dc0c",
			107 => x"020a0608",
			108 => x"09016304",
			109 => x"ffcc01c5",
			110 => x"000001c5",
			111 => x"000001c5",
			112 => x"000001c5",
			113 => x"0100de08",
			114 => x"020a0604",
			115 => x"ffb301e9",
			116 => x"000001e9",
			117 => x"05073908",
			118 => x"040c3204",
			119 => x"000001e9",
			120 => x"002701e9",
			121 => x"000001e9",
			122 => x"0100ad04",
			123 => x"ffb1020d",
			124 => x"0e078e0c",
			125 => x"06016f08",
			126 => x"0705d004",
			127 => x"002f020d",
			128 => x"0000020d",
			129 => x"0000020d",
			130 => x"0000020d",
			131 => x"040c8504",
			132 => x"fff40231",
			133 => x"0209ce04",
			134 => x"00000231",
			135 => x"020a6308",
			136 => x"04120c04",
			137 => x"00460231",
			138 => x"00000231",
			139 => x"00000231",
			140 => x"040d5504",
			141 => x"ffde0255",
			142 => x"0d07080c",
			143 => x"0e054b04",
			144 => x"00000255",
			145 => x"0d066a04",
			146 => x"00000255",
			147 => x"00250255",
			148 => x"00000255",
			149 => x"0100c508",
			150 => x"040fc604",
			151 => x"ff870281",
			152 => x"00000281",
			153 => x"0e07580c",
			154 => x"07057504",
			155 => x"00000281",
			156 => x"0100ca04",
			157 => x"00000281",
			158 => x"00710281",
			159 => x"00000281",
			160 => x"0100ca08",
			161 => x"0410bb04",
			162 => x"ff9902ad",
			163 => x"000002ad",
			164 => x"0e073b0c",
			165 => x"07057504",
			166 => x"000002ad",
			167 => x"06017304",
			168 => x"004d02ad",
			169 => x"000002ad",
			170 => x"000002ad",
			171 => x"0209c90c",
			172 => x"00041004",
			173 => x"000002e1",
			174 => x"0c056404",
			175 => x"ff5e02e1",
			176 => x"000002e1",
			177 => x"0f09150c",
			178 => x"0a02f308",
			179 => x"0c051104",
			180 => x"000002e1",
			181 => x"009a02e1",
			182 => x"000002e1",
			183 => x"000002e1",
			184 => x"040caf04",
			185 => x"ff5d0315",
			186 => x"0b06090c",
			187 => x"0100ca04",
			188 => x"00000315",
			189 => x"07057504",
			190 => x"00000315",
			191 => x"00a80315",
			192 => x"08033a04",
			193 => x"00000315",
			194 => x"0e073b04",
			195 => x"00000315",
			196 => x"ff8c0315",
			197 => x"09012708",
			198 => x"020a0604",
			199 => x"ff8f0349",
			200 => x"00000349",
			201 => x"0e075810",
			202 => x"0c052804",
			203 => x"00000349",
			204 => x"02094304",
			205 => x"00000349",
			206 => x"06017c04",
			207 => x"00580349",
			208 => x"00000349",
			209 => x"00000349",
			210 => x"09010f04",
			211 => x"ffae0375",
			212 => x"0e078e10",
			213 => x"06016f0c",
			214 => x"0b05a704",
			215 => x"00000375",
			216 => x"0f080504",
			217 => x"00000375",
			218 => x"00320375",
			219 => x"00000375",
			220 => x"00000375",
			221 => x"02099a0c",
			222 => x"07058c08",
			223 => x"0c056304",
			224 => x"fec703b9",
			225 => x"000003b9",
			226 => x"000003b9",
			227 => x"0f08cd10",
			228 => x"0803960c",
			229 => x"0e073b08",
			230 => x"0100bb04",
			231 => x"000003b9",
			232 => x"00fd03b9",
			233 => x"000003b9",
			234 => x"000003b9",
			235 => x"0e078e04",
			236 => x"000003b9",
			237 => x"ff9803b9",
			238 => x"040c8504",
			239 => x"ff0803f5",
			240 => x"0100ca08",
			241 => x"04112a04",
			242 => x"ff8c03f5",
			243 => x"000003f5",
			244 => x"0601700c",
			245 => x"0307c408",
			246 => x"0a02a504",
			247 => x"005d03f5",
			248 => x"000003f5",
			249 => x"fff803f5",
			250 => x"0e07dc04",
			251 => x"00cd03f5",
			252 => x"000003f5",
			253 => x"040c8504",
			254 => x"00000429",
			255 => x"06017814",
			256 => x"01009204",
			257 => x"00000429",
			258 => x"0307c40c",
			259 => x"0f08cd08",
			260 => x"07054904",
			261 => x"00000429",
			262 => x"00600429",
			263 => x"00000429",
			264 => x"00000429",
			265 => x"00000429",
			266 => x"040c8504",
			267 => x"ff14046d",
			268 => x"0100ca08",
			269 => x"04112a04",
			270 => x"ff97046d",
			271 => x"0000046d",
			272 => x"06017010",
			273 => x"0f08aa08",
			274 => x"0a02a004",
			275 => x"002f046d",
			276 => x"0000046d",
			277 => x"0a028d04",
			278 => x"0000046d",
			279 => x"ffe9046d",
			280 => x"0f093d04",
			281 => x"00bb046d",
			282 => x"0000046d",
			283 => x"02094304",
			284 => x"fe8e04b9",
			285 => x"06016f0c",
			286 => x"01009204",
			287 => x"000004b9",
			288 => x"0f08f904",
			289 => x"013004b9",
			290 => x"000004b9",
			291 => x"0100de0c",
			292 => x"07060008",
			293 => x"0a029d04",
			294 => x"000004b9",
			295 => x"fefc04b9",
			296 => x"000004b9",
			297 => x"0e07dc08",
			298 => x"0a029204",
			299 => x"000004b9",
			300 => x"00fc04b9",
			301 => x"ff7604b9",
			302 => x"040cc608",
			303 => x"040cb604",
			304 => x"fe950505",
			305 => x"00000505",
			306 => x"01009204",
			307 => x"ff0f0505",
			308 => x"0506d20c",
			309 => x"06017d08",
			310 => x"0a030404",
			311 => x"01590505",
			312 => x"00000505",
			313 => x"00000505",
			314 => x"0100df04",
			315 => x"ff1e0505",
			316 => x"0f094508",
			317 => x"0209c104",
			318 => x"00000505",
			319 => x"01100505",
			320 => x"00000505",
			321 => x"0209b114",
			322 => x"0100cd04",
			323 => x"fe780569",
			324 => x"0506e20c",
			325 => x"0209ab08",
			326 => x"0e078e04",
			327 => x"00eb0569",
			328 => x"00000569",
			329 => x"00000569",
			330 => x"fe9c0569",
			331 => x"06016b0c",
			332 => x"01009204",
			333 => x"00000569",
			334 => x"03089d04",
			335 => x"022a0569",
			336 => x"00000569",
			337 => x"0f092a10",
			338 => x"09015804",
			339 => x"ff380569",
			340 => x"0209c108",
			341 => x"0307c404",
			342 => x"00000569",
			343 => x"ffd40569",
			344 => x"01470569",
			345 => x"fed00569",
			346 => x"0209b10c",
			347 => x"0c056308",
			348 => x"0705a304",
			349 => x"fef205b5",
			350 => x"000005b5",
			351 => x"000005b5",
			352 => x"0c059d18",
			353 => x"0c052804",
			354 => x"000005b5",
			355 => x"020a2d10",
			356 => x"0209c104",
			357 => x"000005b5",
			358 => x"040caf04",
			359 => x"000005b5",
			360 => x"00055404",
			361 => x"00eb05b5",
			362 => x"000005b5",
			363 => x"000005b5",
			364 => x"000005b5",
			365 => x"02094304",
			366 => x"fe8a05f9",
			367 => x"0f09331c",
			368 => x"0209ce10",
			369 => x"0a029d0c",
			370 => x"0e078e08",
			371 => x"0100cf04",
			372 => x"000005f9",
			373 => x"00fd05f9",
			374 => x"000005f9",
			375 => x"ff3105f9",
			376 => x"0a030408",
			377 => x"0c051104",
			378 => x"000005f9",
			379 => x"010b05f9",
			380 => x"000005f9",
			381 => x"fefc05f9",
			382 => x"0209b118",
			383 => x"0100cd04",
			384 => x"fe7a065d",
			385 => x"0b06060c",
			386 => x"0209ab08",
			387 => x"0e07dc04",
			388 => x"00d3065d",
			389 => x"0000065d",
			390 => x"0000065d",
			391 => x"0e073b04",
			392 => x"0000065d",
			393 => x"feac065d",
			394 => x"0f092a18",
			395 => x"06016b08",
			396 => x"01009204",
			397 => x"0000065d",
			398 => x"01fb065d",
			399 => x"09015804",
			400 => x"ff4b065d",
			401 => x"0209c108",
			402 => x"0d071604",
			403 => x"0000065d",
			404 => x"ffea065d",
			405 => x"013c065d",
			406 => x"fed9065d",
			407 => x"040c4404",
			408 => x"ffe10699",
			409 => x"01009204",
			410 => x"00000699",
			411 => x"020a2d14",
			412 => x"06017c10",
			413 => x"0c059d0c",
			414 => x"07054704",
			415 => x"00000699",
			416 => x"0c052504",
			417 => x"00000699",
			418 => x"00660699",
			419 => x"00000699",
			420 => x"00000699",
			421 => x"00000699",
			422 => x"01009204",
			423 => x"ff1906ed",
			424 => x"06016f0c",
			425 => x"040c3204",
			426 => x"000006ed",
			427 => x"06016a04",
			428 => x"009006ed",
			429 => x"000006ed",
			430 => x"08034814",
			431 => x"0c059910",
			432 => x"06017004",
			433 => x"000006ed",
			434 => x"06017908",
			435 => x"0003fb04",
			436 => x"000006ed",
			437 => x"003a06ed",
			438 => x"000006ed",
			439 => x"000006ed",
			440 => x"0100df04",
			441 => x"ff8306ed",
			442 => x"000006ed",
			443 => x"0100b004",
			444 => x"fe6d0749",
			445 => x"0c059b24",
			446 => x"0e075814",
			447 => x"0d06f90c",
			448 => x"0f082b04",
			449 => x"00000749",
			450 => x"0b05a704",
			451 => x"00000749",
			452 => x"01d40749",
			453 => x"09015a04",
			454 => x"fecc0749",
			455 => x"01690749",
			456 => x"0c056308",
			457 => x"0a028d04",
			458 => x"00000749",
			459 => x"fe4c0749",
			460 => x"0e07dc04",
			461 => x"01420749",
			462 => x"00000749",
			463 => x"0e073b04",
			464 => x"00000749",
			465 => x"fe840749",
			466 => x"09011304",
			467 => x"fe6e07a5",
			468 => x"0307b014",
			469 => x"040c4404",
			470 => x"ffc307a5",
			471 => x"0803b40c",
			472 => x"0c052804",
			473 => x"000007a5",
			474 => x"0209dd04",
			475 => x"00fb07a5",
			476 => x"01fa07a5",
			477 => x"000007a5",
			478 => x"0d077014",
			479 => x"0209c10c",
			480 => x"0a028d08",
			481 => x"040c3204",
			482 => x"000007a5",
			483 => x"009407a5",
			484 => x"fe5107a5",
			485 => x"0f093d04",
			486 => x"016d07a5",
			487 => x"000007a5",
			488 => x"fe8007a5",
			489 => x"040cbf08",
			490 => x"040cb604",
			491 => x"fe8d0819",
			492 => x"00000819",
			493 => x"0209c914",
			494 => x"08033a0c",
			495 => x"0f08b808",
			496 => x"0100cf04",
			497 => x"00000819",
			498 => x"00b90819",
			499 => x"00000819",
			500 => x"0a028804",
			501 => x"00000819",
			502 => x"fee00819",
			503 => x"03079c14",
			504 => x"0a030410",
			505 => x"0209ce04",
			506 => x"00000819",
			507 => x"020a2d08",
			508 => x"07054704",
			509 => x"00000819",
			510 => x"01d80819",
			511 => x"00000819",
			512 => x"00000819",
			513 => x"0100dc04",
			514 => x"ff260819",
			515 => x"0d078804",
			516 => x"00bb0819",
			517 => x"00000819",
			518 => x"0100b404",
			519 => x"fe690865",
			520 => x"0d077020",
			521 => x"040c3204",
			522 => x"feeb0865",
			523 => x"0506d20c",
			524 => x"0c052804",
			525 => x"002a0865",
			526 => x"0004bc04",
			527 => x"01900865",
			528 => x"02b20865",
			529 => x"09015a04",
			530 => x"fe6f0865",
			531 => x"0c054804",
			532 => x"00000865",
			533 => x"0100df04",
			534 => x"00000865",
			535 => x"017b0865",
			536 => x"fe680865",
			537 => x"0100ad04",
			538 => x"fe6b08c1",
			539 => x"0d077028",
			540 => x"0209c11c",
			541 => x"0e07580c",
			542 => x"0a02b008",
			543 => x"02094304",
			544 => x"000008c1",
			545 => x"017a08c1",
			546 => x"ff0d08c1",
			547 => x"0c056508",
			548 => x"0a028d04",
			549 => x"000008c1",
			550 => x"fe0b08c1",
			551 => x"0307f404",
			552 => x"002608c1",
			553 => x"000008c1",
			554 => x"06018508",
			555 => x"0a02e404",
			556 => x"01b008c1",
			557 => x"000008c1",
			558 => x"000008c1",
			559 => x"fe7208c1",
			560 => x"02096c08",
			561 => x"02094904",
			562 => x"fe730935",
			563 => x"00000935",
			564 => x"0e05e010",
			565 => x"01009204",
			566 => x"00000935",
			567 => x"0b058704",
			568 => x"06280935",
			569 => x"0100a104",
			570 => x"00000935",
			571 => x"02050935",
			572 => x"0e07dc20",
			573 => x"08033f0c",
			574 => x"0705ba04",
			575 => x"01600935",
			576 => x"0705ce04",
			577 => x"00000935",
			578 => x"00790935",
			579 => x"0209ce0c",
			580 => x"0b05d908",
			581 => x"0100b404",
			582 => x"00000935",
			583 => x"003a0935",
			584 => x"febd0935",
			585 => x"08037e04",
			586 => x"01300935",
			587 => x"ff6a0935",
			588 => x"fea80935",
			589 => x"02094304",
			590 => x"fe970991",
			591 => x"0f092a28",
			592 => x"08033f0c",
			593 => x"040c3204",
			594 => x"00000991",
			595 => x"0100cf04",
			596 => x"00000991",
			597 => x"01190991",
			598 => x"06016608",
			599 => x"01009204",
			600 => x"00000991",
			601 => x"00e40991",
			602 => x"0209e808",
			603 => x"06016a04",
			604 => x"00000991",
			605 => x"ff3c0991",
			606 => x"09015a08",
			607 => x"06016c04",
			608 => x"00000991",
			609 => x"ffd20991",
			610 => x"00a80991",
			611 => x"ff240991",
			612 => x"02096008",
			613 => x"02094304",
			614 => x"fe620a15",
			615 => x"fece0a15",
			616 => x"0c059c28",
			617 => x"0100ad0c",
			618 => x"0c054804",
			619 => x"fe740a15",
			620 => x"00055404",
			621 => x"06370a15",
			622 => x"feb30a15",
			623 => x"0306c504",
			624 => x"15610a15",
			625 => x"03073b08",
			626 => x"0a02db04",
			627 => x"051f0a15",
			628 => x"fff50a15",
			629 => x"09015808",
			630 => x"0a029904",
			631 => x"004f0a15",
			632 => x"fd210a15",
			633 => x"03087504",
			634 => x"01bc0a15",
			635 => x"fea10a15",
			636 => x"0705d10c",
			637 => x"0506d504",
			638 => x"ff0c0a15",
			639 => x"0c05a004",
			640 => x"ff7f0a15",
			641 => x"014f0a15",
			642 => x"0c059d04",
			643 => x"00000a15",
			644 => x"fe650a15",
			645 => x"02096c0c",
			646 => x"02094904",
			647 => x"fe680a81",
			648 => x"02094d04",
			649 => x"00000a81",
			650 => x"ff100a81",
			651 => x"0f093328",
			652 => x"09011304",
			653 => x"fe910a81",
			654 => x"0506d20c",
			655 => x"0c051104",
			656 => x"00000a81",
			657 => x"0a02e404",
			658 => x"01bd0a81",
			659 => x"00000a81",
			660 => x"0209c90c",
			661 => x"08033a08",
			662 => x"0307f404",
			663 => x"015a0a81",
			664 => x"ff270a81",
			665 => x"fe140a81",
			666 => x"09015a04",
			667 => x"ff6e0a81",
			668 => x"0705a104",
			669 => x"00000a81",
			670 => x"01ac0a81",
			671 => x"fe640a81",
			672 => x"0100b404",
			673 => x"fe680add",
			674 => x"0d077028",
			675 => x"040c3204",
			676 => x"feda0add",
			677 => x"0506d20c",
			678 => x"0004c908",
			679 => x"0a02c704",
			680 => x"01970add",
			681 => x"00000add",
			682 => x"036c0add",
			683 => x"0100df0c",
			684 => x"0a02a904",
			685 => x"00d20add",
			686 => x"0f08c604",
			687 => x"fe460add",
			688 => x"00000add",
			689 => x"0c056308",
			690 => x"0209c104",
			691 => x"00000add",
			692 => x"00de0add",
			693 => x"01a80add",
			694 => x"fe660add",
			695 => x"02096004",
			696 => x"fe670b5b",
			697 => x"0c059d2c",
			698 => x"0100ad04",
			699 => x"fe7b0b5b",
			700 => x"0e075810",
			701 => x"0803b40c",
			702 => x"0100d404",
			703 => x"034d0b5b",
			704 => x"0100da04",
			705 => x"00250b5b",
			706 => x"01ae0b5b",
			707 => x"fea50b5b",
			708 => x"0100e80c",
			709 => x"040d8808",
			710 => x"040c5204",
			711 => x"fef10b5b",
			712 => x"00000b5b",
			713 => x"fbf10b5b",
			714 => x"0e07dc08",
			715 => x"0209ce04",
			716 => x"009f0b5b",
			717 => x"03610b5b",
			718 => x"febf0b5b",
			719 => x"0705d10c",
			720 => x"0e073b08",
			721 => x"0e03bd04",
			722 => x"ff930b5b",
			723 => x"00f00b5b",
			724 => x"fe7a0b5b",
			725 => x"fe660b5b",
			726 => x"00000b5d",
			727 => x"00000b61",
			728 => x"00000b65",
			729 => x"00000b69",
			730 => x"00000b6d",
			731 => x"00000b71",
			732 => x"00000b75",
			733 => x"00000b79",
			734 => x"00000b7d",
			735 => x"00000b81",
			736 => x"00000b85",
			737 => x"00000b89",
			738 => x"00000b8d",
			739 => x"00000b91",
			740 => x"00000b95",
			741 => x"00000b99",
			742 => x"00000b9d",
			743 => x"00000ba1",
			744 => x"00000ba5",
			745 => x"00000ba9",
			746 => x"00000bad",
			747 => x"00000bb1",
			748 => x"00000bb5",
			749 => x"00000bb9",
			750 => x"00000bbd",
			751 => x"00000bc1",
			752 => x"00000bc5",
			753 => x"00000bc9",
			754 => x"00000bcd",
			755 => x"0410bb04",
			756 => x"fffb0bd9",
			757 => x"00000bd9",
			758 => x"040d5504",
			759 => x"fff90be5",
			760 => x"00000be5",
			761 => x"0209ce04",
			762 => x"ffe90bf1",
			763 => x"00000bf1",
			764 => x"040fc604",
			765 => x"ffee0bfd",
			766 => x"00000bfd",
			767 => x"0100ca04",
			768 => x"ffe70c09",
			769 => x"00000c09",
			770 => x"020a0604",
			771 => x"fffd0c15",
			772 => x"00000c15",
			773 => x"040fc604",
			774 => x"fffb0c21",
			775 => x"00000c21",
			776 => x"040c4404",
			777 => x"fff20c35",
			778 => x"04120c04",
			779 => x"00060c35",
			780 => x"00000c35",
			781 => x"040c8504",
			782 => x"00000c49",
			783 => x"04120c04",
			784 => x"000b0c49",
			785 => x"00000c49",
			786 => x"040cbf04",
			787 => x"00000c5d",
			788 => x"04120c04",
			789 => x"000f0c5d",
			790 => x"00000c5d",
			791 => x"0209c104",
			792 => x"ffff0c71",
			793 => x"020a2d04",
			794 => x"00300c71",
			795 => x"00000c71",
			796 => x"0209ce04",
			797 => x"fff50c85",
			798 => x"020a6b04",
			799 => x"00290c85",
			800 => x"00000c85",
			801 => x"040d5508",
			802 => x"0a028b04",
			803 => x"00000c99",
			804 => x"ffdf0c99",
			805 => x"00000c99",
			806 => x"0100ca04",
			807 => x"ff960cb5",
			808 => x"0e075808",
			809 => x"07057504",
			810 => x"00000cb5",
			811 => x"00800cb5",
			812 => x"00000cb5",
			813 => x"04112a0c",
			814 => x"0100dc08",
			815 => x"09016104",
			816 => x"ff910cd1",
			817 => x"00000cd1",
			818 => x"00000cd1",
			819 => x"00000cd1",
			820 => x"040c8504",
			821 => x"fff20ced",
			822 => x"0209b104",
			823 => x"00000ced",
			824 => x"020a6b04",
			825 => x"00190ced",
			826 => x"00000ced",
			827 => x"0901630c",
			828 => x"0410bb08",
			829 => x"0100dc04",
			830 => x"ffb20d09",
			831 => x"00000d09",
			832 => x"00000d09",
			833 => x"00000d09",
			834 => x"0100dc0c",
			835 => x"020a0608",
			836 => x"09016304",
			837 => x"ffd40d25",
			838 => x"00000d25",
			839 => x"00000d25",
			840 => x"00000d25",
			841 => x"0100ca04",
			842 => x"ff4d0d49",
			843 => x"0d07550c",
			844 => x"0c058008",
			845 => x"0e07dc04",
			846 => x"00990d49",
			847 => x"00000d49",
			848 => x"00000d49",
			849 => x"00000d49",
			850 => x"040c4404",
			851 => x"ffe20d6d",
			852 => x"09010f04",
			853 => x"00000d6d",
			854 => x"020a6b08",
			855 => x"07055f04",
			856 => x"00000d6d",
			857 => x"00230d6d",
			858 => x"00000d6d",
			859 => x"040c8504",
			860 => x"fff60d91",
			861 => x"0209ce04",
			862 => x"00000d91",
			863 => x"020a6308",
			864 => x"04120c04",
			865 => x"003d0d91",
			866 => x"00000d91",
			867 => x"00000d91",
			868 => x"040d5504",
			869 => x"ffe50db5",
			870 => x"0d07080c",
			871 => x"0d066a04",
			872 => x"00000db5",
			873 => x"0b061b04",
			874 => x"001d0db5",
			875 => x"00000db5",
			876 => x"00000db5",
			877 => x"0100ca08",
			878 => x"0410bb04",
			879 => x"ff840de1",
			880 => x"00000de1",
			881 => x"0e073b0c",
			882 => x"07057504",
			883 => x"00000de1",
			884 => x"06017304",
			885 => x"005d0de1",
			886 => x"00000de1",
			887 => x"00000de1",
			888 => x"0100de08",
			889 => x"020a0604",
			890 => x"ffaa0e0d",
			891 => x"00000e0d",
			892 => x"0b065b0c",
			893 => x"07058c04",
			894 => x"00000e0d",
			895 => x"040c3204",
			896 => x"00000e0d",
			897 => x"00400e0d",
			898 => x"00000e0d",
			899 => x"0209c90c",
			900 => x"00041004",
			901 => x"00000e41",
			902 => x"06017404",
			903 => x"ff7c0e41",
			904 => x"00000e41",
			905 => x"0f09150c",
			906 => x"0100ca04",
			907 => x"00000e41",
			908 => x"020a3a04",
			909 => x"009d0e41",
			910 => x"00000e41",
			911 => x"00000e41",
			912 => x"040caf04",
			913 => x"ff670e75",
			914 => x"0b06090c",
			915 => x"0100ca04",
			916 => x"00000e75",
			917 => x"07057504",
			918 => x"00000e75",
			919 => x"00990e75",
			920 => x"08033a04",
			921 => x"00000e75",
			922 => x"0d071604",
			923 => x"00000e75",
			924 => x"ffa90e75",
			925 => x"09014004",
			926 => x"ff6c0ea1",
			927 => x"0d075510",
			928 => x"0c05800c",
			929 => x"07055f04",
			930 => x"00000ea1",
			931 => x"0e07dc04",
			932 => x"00710ea1",
			933 => x"00000ea1",
			934 => x"00000ea1",
			935 => x"00000ea1",
			936 => x"040c4404",
			937 => x"ffe90ecd",
			938 => x"0c052504",
			939 => x"00000ecd",
			940 => x"020a2d0c",
			941 => x"04120c08",
			942 => x"0c059d04",
			943 => x"00460ecd",
			944 => x"00000ecd",
			945 => x"00000ecd",
			946 => x"00000ecd",
			947 => x"07054908",
			948 => x"0100d404",
			949 => x"fedf0f11",
			950 => x"00000f11",
			951 => x"0307c410",
			952 => x"0100ca04",
			953 => x"00000f11",
			954 => x"07057504",
			955 => x"00000f11",
			956 => x"0c058004",
			957 => x"01060f11",
			958 => x"00000f11",
			959 => x"0506d504",
			960 => x"00000f11",
			961 => x"0a029204",
			962 => x"ff3c0f11",
			963 => x"00000f11",
			964 => x"040fc618",
			965 => x"09014d04",
			966 => x"fe7f0f5d",
			967 => x"0e073b08",
			968 => x"09015804",
			969 => x"00000f5d",
			970 => x"01370f5d",
			971 => x"0b060904",
			972 => x"00000f5d",
			973 => x"0c054504",
			974 => x"00000f5d",
			975 => x"fee00f5d",
			976 => x"0a03040c",
			977 => x"0d06c708",
			978 => x"0209d404",
			979 => x"00000f5d",
			980 => x"02360f5d",
			981 => x"00000f5d",
			982 => x"ff420f5d",
			983 => x"040c4404",
			984 => x"ff480f99",
			985 => x"0209ce08",
			986 => x"08033a04",
			987 => x"00230f99",
			988 => x"ff970f99",
			989 => x"06018310",
			990 => x"0c051104",
			991 => x"00000f99",
			992 => x"0a030408",
			993 => x"0c059d04",
			994 => x"00bc0f99",
			995 => x"00000f99",
			996 => x"00000f99",
			997 => x"00000f99",
			998 => x"02099a0c",
			999 => x"0c056308",
			1000 => x"07058c04",
			1001 => x"fea10fe5",
			1002 => x"00000fe5",
			1003 => x"00000fe5",
			1004 => x"0f093318",
			1005 => x"0100ca10",
			1006 => x"0f080e0c",
			1007 => x"00055408",
			1008 => x"00050804",
			1009 => x"00000fe5",
			1010 => x"00640fe5",
			1011 => x"00000fe5",
			1012 => x"ffba0fe5",
			1013 => x"0209be04",
			1014 => x"00000fe5",
			1015 => x"00fa0fe5",
			1016 => x"ff670fe5",
			1017 => x"0100d420",
			1018 => x"0100ca18",
			1019 => x"0209c104",
			1020 => x"bd1c1039",
			1021 => x"0209c908",
			1022 => x"01004104",
			1023 => x"be031039",
			1024 => x"cb891039",
			1025 => x"06016b08",
			1026 => x"01009004",
			1027 => x"bd301039",
			1028 => x"cb891039",
			1029 => x"bd1e1039",
			1030 => x"0e071504",
			1031 => x"e5f91039",
			1032 => x"bd241039",
			1033 => x"0e078e04",
			1034 => x"19911039",
			1035 => x"0e07dc04",
			1036 => x"d83d1039",
			1037 => x"bd1c1039",
			1038 => x"040cc608",
			1039 => x"040cb604",
			1040 => x"fe9b1085",
			1041 => x"00001085",
			1042 => x"01009204",
			1043 => x"ff1e1085",
			1044 => x"0d07160c",
			1045 => x"06017d08",
			1046 => x"0a030404",
			1047 => x"011d1085",
			1048 => x"00001085",
			1049 => x"00001085",
			1050 => x"0100df04",
			1051 => x"ff2f1085",
			1052 => x"06018808",
			1053 => x"0209c104",
			1054 => x"00001085",
			1055 => x"00e31085",
			1056 => x"00001085",
			1057 => x"0209b10c",
			1058 => x"09017a08",
			1059 => x"0c056304",
			1060 => x"fe9c10d9",
			1061 => x"000010d9",
			1062 => x"000010d9",
			1063 => x"0f090d18",
			1064 => x"0209ce04",
			1065 => x"000010d9",
			1066 => x"0c052804",
			1067 => x"000010d9",
			1068 => x"0a03040c",
			1069 => x"020a3a08",
			1070 => x"06017c04",
			1071 => x"012710d9",
			1072 => x"000010d9",
			1073 => x"000010d9",
			1074 => x"000010d9",
			1075 => x"0f093304",
			1076 => x"000010d9",
			1077 => x"ff4c10d9",
			1078 => x"02099a0c",
			1079 => x"07058c08",
			1080 => x"0c056304",
			1081 => x"feed1125",
			1082 => x"00001125",
			1083 => x"00001125",
			1084 => x"0c059b18",
			1085 => x"0c052804",
			1086 => x"00001125",
			1087 => x"0209c104",
			1088 => x"00001125",
			1089 => x"020a2d0c",
			1090 => x"040caf04",
			1091 => x"00001125",
			1092 => x"00055404",
			1093 => x"00db1125",
			1094 => x"00001125",
			1095 => x"00001125",
			1096 => x"00001125",
			1097 => x"02099a08",
			1098 => x"0c056304",
			1099 => x"ff061169",
			1100 => x"00001169",
			1101 => x"0c059d18",
			1102 => x"0c052804",
			1103 => x"00001169",
			1104 => x"0209c104",
			1105 => x"00001169",
			1106 => x"020a2d0c",
			1107 => x"040caf04",
			1108 => x"00001169",
			1109 => x"00055404",
			1110 => x"00cb1169",
			1111 => x"00001169",
			1112 => x"00001169",
			1113 => x"00001169",
			1114 => x"07054904",
			1115 => x"ff1111bd",
			1116 => x"0307c414",
			1117 => x"0a02d710",
			1118 => x"09011304",
			1119 => x"000011bd",
			1120 => x"0c052804",
			1121 => x"000011bd",
			1122 => x"040c5204",
			1123 => x"000011bd",
			1124 => x"00ab11bd",
			1125 => x"000011bd",
			1126 => x"06017308",
			1127 => x"0b060904",
			1128 => x"000011bd",
			1129 => x"ffa011bd",
			1130 => x"06017908",
			1131 => x"0b064b04",
			1132 => x"003611bd",
			1133 => x"000011bd",
			1134 => x"000011bd",
			1135 => x"040c4404",
			1136 => x"ffe611f9",
			1137 => x"01009204",
			1138 => x"000011f9",
			1139 => x"020a2d14",
			1140 => x"06017c10",
			1141 => x"0c059d0c",
			1142 => x"07054704",
			1143 => x"000011f9",
			1144 => x"0c052504",
			1145 => x"000011f9",
			1146 => x"005a11f9",
			1147 => x"000011f9",
			1148 => x"000011f9",
			1149 => x"000011f9",
			1150 => x"07054908",
			1151 => x"0100d204",
			1152 => x"fe92125d",
			1153 => x"0000125d",
			1154 => x"0c059b24",
			1155 => x"0100dc18",
			1156 => x"06016a0c",
			1157 => x"0f07d504",
			1158 => x"0000125d",
			1159 => x"0003d804",
			1160 => x"0000125d",
			1161 => x"010a125d",
			1162 => x"0506f108",
			1163 => x"09016304",
			1164 => x"ff0b125d",
			1165 => x"0000125d",
			1166 => x"0000125d",
			1167 => x"0e07dc08",
			1168 => x"08034804",
			1169 => x"0120125d",
			1170 => x"0000125d",
			1171 => x"0000125d",
			1172 => x"0705ba04",
			1173 => x"0000125d",
			1174 => x"ff21125d",
			1175 => x"0100b404",
			1176 => x"fe6912a1",
			1177 => x"0d07701c",
			1178 => x"040c3204",
			1179 => x"fefb12a1",
			1180 => x"0506d208",
			1181 => x"0c052804",
			1182 => x"001c12a1",
			1183 => x"01d012a1",
			1184 => x"09015a04",
			1185 => x"fe8812a1",
			1186 => x"0c054804",
			1187 => x"000012a1",
			1188 => x"0100df04",
			1189 => x"000012a1",
			1190 => x"016f12a1",
			1191 => x"fe6a12a1",
			1192 => x"0100ad04",
			1193 => x"fe6f12fd",
			1194 => x"0e073b14",
			1195 => x"0803b410",
			1196 => x"02094304",
			1197 => x"000012fd",
			1198 => x"020a0608",
			1199 => x"0f08c604",
			1200 => x"010b12fd",
			1201 => x"000012fd",
			1202 => x"01f912fd",
			1203 => x"000012fd",
			1204 => x"0d077014",
			1205 => x"0209c10c",
			1206 => x"0a028d08",
			1207 => x"040c3204",
			1208 => x"000012fd",
			1209 => x"008812fd",
			1210 => x"fe7012fd",
			1211 => x"0f093d04",
			1212 => x"016112fd",
			1213 => x"000012fd",
			1214 => x"fe8512fd",
			1215 => x"040cbf04",
			1216 => x"feb51361",
			1217 => x"0e073b1c",
			1218 => x"01009204",
			1219 => x"ff8b1361",
			1220 => x"0d06c70c",
			1221 => x"06017308",
			1222 => x"0c052804",
			1223 => x"00001361",
			1224 => x"01231361",
			1225 => x"00001361",
			1226 => x"0a02bf08",
			1227 => x"0f087204",
			1228 => x"00001361",
			1229 => x"00d11361",
			1230 => x"ffb01361",
			1231 => x"08033a08",
			1232 => x"0705ba04",
			1233 => x"003d1361",
			1234 => x"00001361",
			1235 => x"0d071604",
			1236 => x"00001361",
			1237 => x"0b061b04",
			1238 => x"fee81361",
			1239 => x"00001361",
			1240 => x"02094304",
			1241 => x"fe6a13ad",
			1242 => x"0f093320",
			1243 => x"09011304",
			1244 => x"fe9c13ad",
			1245 => x"0209c114",
			1246 => x"08033a08",
			1247 => x"0e078e04",
			1248 => x"018813ad",
			1249 => x"ff3413ad",
			1250 => x"0506d208",
			1251 => x"09014404",
			1252 => x"000013ad",
			1253 => x"006013ad",
			1254 => x"fe0813ad",
			1255 => x"0a02e404",
			1256 => x"01be13ad",
			1257 => x"000013ad",
			1258 => x"fe6e13ad",
			1259 => x"0100ad04",
			1260 => x"fe711411",
			1261 => x"0d077028",
			1262 => x"0209c118",
			1263 => x"08033910",
			1264 => x"0003c404",
			1265 => x"ffb41411",
			1266 => x"0f08cd08",
			1267 => x"0100cf04",
			1268 => x"00001411",
			1269 => x"014e1411",
			1270 => x"00001411",
			1271 => x"0506d204",
			1272 => x"00001411",
			1273 => x"fe931411",
			1274 => x"0c052804",
			1275 => x"00001411",
			1276 => x"0803b408",
			1277 => x"0f093d04",
			1278 => x"019f1411",
			1279 => x"00001411",
			1280 => x"00001411",
			1281 => x"05072904",
			1282 => x"00001411",
			1283 => x"fe8c1411",
			1284 => x"02096c08",
			1285 => x"02094904",
			1286 => x"fe751485",
			1287 => x"00001485",
			1288 => x"06016a10",
			1289 => x"0705be0c",
			1290 => x"01009204",
			1291 => x"00001485",
			1292 => x"0c052804",
			1293 => x"00001485",
			1294 => x"026d1485",
			1295 => x"00001485",
			1296 => x"0f093320",
			1297 => x"0100de10",
			1298 => x"0f08b808",
			1299 => x"0a029d04",
			1300 => x"00001485",
			1301 => x"fed51485",
			1302 => x"09015a04",
			1303 => x"00001485",
			1304 => x"00541485",
			1305 => x"0209c10c",
			1306 => x"0307c404",
			1307 => x"006d1485",
			1308 => x"0c056604",
			1309 => x"ff701485",
			1310 => x"00001485",
			1311 => x"01561485",
			1312 => x"feb41485",
			1313 => x"02094304",
			1314 => x"fe6a14f1",
			1315 => x"0c05b42c",
			1316 => x"0209c11c",
			1317 => x"08033a0c",
			1318 => x"0e078e08",
			1319 => x"0100cf04",
			1320 => x"000014f1",
			1321 => x"018114f1",
			1322 => x"ff2414f1",
			1323 => x"0c056508",
			1324 => x"0a028804",
			1325 => x"000014f1",
			1326 => x"fe4814f1",
			1327 => x"0306ff04",
			1328 => x"000014f1",
			1329 => x"000414f1",
			1330 => x"0a02e40c",
			1331 => x"040caf04",
			1332 => x"ff8614f1",
			1333 => x"0c051104",
			1334 => x"000014f1",
			1335 => x"01b714f1",
			1336 => x"ff4414f1",
			1337 => x"0c05b804",
			1338 => x"000014f1",
			1339 => x"fe7214f1",
			1340 => x"040caf0c",
			1341 => x"040c8504",
			1342 => x"fe6a1575",
			1343 => x"040c8c04",
			1344 => x"ffe01575",
			1345 => x"fee31575",
			1346 => x"08038524",
			1347 => x"09011304",
			1348 => x"fe8f1575",
			1349 => x"0e073b0c",
			1350 => x"0506d204",
			1351 => x"01ce1575",
			1352 => x"0506d504",
			1353 => x"ffcc1575",
			1354 => x"01ad1575",
			1355 => x"08033a08",
			1356 => x"06017004",
			1357 => x"00aa1575",
			1358 => x"02331575",
			1359 => x"06017404",
			1360 => x"fd781575",
			1361 => x"0e078e04",
			1362 => x"01571575",
			1363 => x"ff131575",
			1364 => x"0a02f310",
			1365 => x"09010f04",
			1366 => x"fe761575",
			1367 => x"07057504",
			1368 => x"04691575",
			1369 => x"0a02db04",
			1370 => x"00001575",
			1371 => x"ff821575",
			1372 => x"fe681575",
			1373 => x"02095704",
			1374 => x"fe6515e9",
			1375 => x"0c059c24",
			1376 => x"0c051108",
			1377 => x"07057504",
			1378 => x"fe7915e9",
			1379 => x"000015e9",
			1380 => x"0a030418",
			1381 => x"0e065a08",
			1382 => x"0209ce04",
			1383 => x"02af15e9",
			1384 => x"07b915e9",
			1385 => x"0506d208",
			1386 => x"0100ca04",
			1387 => x"ff3315e9",
			1388 => x"01de15e9",
			1389 => x"09015a04",
			1390 => x"fd2b15e9",
			1391 => x"011d15e9",
			1392 => x"fe9815e9",
			1393 => x"0705d10c",
			1394 => x"0506d504",
			1395 => x"ff2115e9",
			1396 => x"0c05a004",
			1397 => x"ffa015e9",
			1398 => x"012a15e9",
			1399 => x"0c059d04",
			1400 => x"000015e9",
			1401 => x"fe6615e9",
			1402 => x"0100ad04",
			1403 => x"fe661675",
			1404 => x"0e075820",
			1405 => x"0506d210",
			1406 => x"0e062e04",
			1407 => x"03841675",
			1408 => x"040c4404",
			1409 => x"ff641675",
			1410 => x"0a02c704",
			1411 => x"01b81675",
			1412 => x"00001675",
			1413 => x"0100df0c",
			1414 => x"0f08aa08",
			1415 => x"0e06e204",
			1416 => x"00001675",
			1417 => x"fe571675",
			1418 => x"00651675",
			1419 => x"01951675",
			1420 => x"0d077020",
			1421 => x"0c056514",
			1422 => x"08033708",
			1423 => x"040b4204",
			1424 => x"ff231675",
			1425 => x"004a1675",
			1426 => x"0d070808",
			1427 => x"0506a604",
			1428 => x"ff841675",
			1429 => x"00011675",
			1430 => x"fd561675",
			1431 => x"040c5204",
			1432 => x"ff2a1675",
			1433 => x"09018004",
			1434 => x"004d1675",
			1435 => x"02361675",
			1436 => x"fe621675",
			1437 => x"02096004",
			1438 => x"fe6816fb",
			1439 => x"0c059d30",
			1440 => x"09011304",
			1441 => x"fe7f16fb",
			1442 => x"0e075814",
			1443 => x"0803b410",
			1444 => x"0100d408",
			1445 => x"0f088b04",
			1446 => x"031316fb",
			1447 => x"011516fb",
			1448 => x"0100da04",
			1449 => x"001d16fb",
			1450 => x"01aa16fb",
			1451 => x"fec816fb",
			1452 => x"0100e80c",
			1453 => x"08031404",
			1454 => x"000016fb",
			1455 => x"0b05fa04",
			1456 => x"fef916fb",
			1457 => x"fcc716fb",
			1458 => x"0e07dc08",
			1459 => x"0c056604",
			1460 => x"007716fb",
			1461 => x"02f716fb",
			1462 => x"fecd16fb",
			1463 => x"0705d10c",
			1464 => x"0e073b08",
			1465 => x"0e03bd04",
			1466 => x"ffaa16fb",
			1467 => x"00d416fb",
			1468 => x"febc16fb",
			1469 => x"fe6716fb",
			1470 => x"000016fd",
			1471 => x"00001701",
			1472 => x"00001705",
			1473 => x"00001709",
			1474 => x"0000170d",
			1475 => x"00001711",
			1476 => x"00001715",
			1477 => x"00001719",
			1478 => x"0000171d",
			1479 => x"00001721",
			1480 => x"00001725",
			1481 => x"00001729",
			1482 => x"0000172d",
			1483 => x"00001731",
			1484 => x"00001735",
			1485 => x"00001739",
			1486 => x"0000173d",
			1487 => x"00001741",
			1488 => x"00001745",
			1489 => x"00001749",
			1490 => x"0000174d",
			1491 => x"00001751",
			1492 => x"00001755",
			1493 => x"00001759",
			1494 => x"0000175d",
			1495 => x"00001761",
			1496 => x"00001765",
			1497 => x"00001769",
			1498 => x"0000176d",
			1499 => x"0410bb04",
			1500 => x"ffff1779",
			1501 => x"00001779",
			1502 => x"040d5504",
			1503 => x"fff61785",
			1504 => x"00001785",
			1505 => x"0209ce04",
			1506 => x"ffef1791",
			1507 => x"00001791",
			1508 => x"0004bc04",
			1509 => x"fffd179d",
			1510 => x"0000179d",
			1511 => x"0100ca04",
			1512 => x"ffe917a9",
			1513 => x"000017a9",
			1514 => x"040fc604",
			1515 => x"fff117b5",
			1516 => x"000017b5",
			1517 => x"0209c108",
			1518 => x"0100f304",
			1519 => x"ffa217c9",
			1520 => x"000017c9",
			1521 => x"000017c9",
			1522 => x"040c4404",
			1523 => x"fff417dd",
			1524 => x"04120c04",
			1525 => x"000317dd",
			1526 => x"000017dd",
			1527 => x"0209ce04",
			1528 => x"fff117f1",
			1529 => x"020a2d04",
			1530 => x"000a17f1",
			1531 => x"000017f1",
			1532 => x"040cbf04",
			1533 => x"00001805",
			1534 => x"04120c04",
			1535 => x"000c1805",
			1536 => x"00001805",
			1537 => x"0209c104",
			1538 => x"ffff1819",
			1539 => x"020a2004",
			1540 => x"00281819",
			1541 => x"00001819",
			1542 => x"0209ce04",
			1543 => x"fffc182d",
			1544 => x"020a6b04",
			1545 => x"001d182d",
			1546 => x"0000182d",
			1547 => x"0100dc08",
			1548 => x"0410bb04",
			1549 => x"ffcc1841",
			1550 => x"00001841",
			1551 => x"00001841",
			1552 => x"040fc60c",
			1553 => x"0100dc08",
			1554 => x"09016304",
			1555 => x"ff6b185d",
			1556 => x"0000185d",
			1557 => x"0000185d",
			1558 => x"0000185d",
			1559 => x"04112a0c",
			1560 => x"0100dc08",
			1561 => x"09016104",
			1562 => x"ff9d1879",
			1563 => x"00001879",
			1564 => x"00001879",
			1565 => x"00001879",
			1566 => x"040cbf04",
			1567 => x"fff51895",
			1568 => x"0209b104",
			1569 => x"00001895",
			1570 => x"020a6b04",
			1571 => x"00181895",
			1572 => x"00001895",
			1573 => x"0901630c",
			1574 => x"0410bb08",
			1575 => x"0100dc04",
			1576 => x"ffb918b1",
			1577 => x"000018b1",
			1578 => x"000018b1",
			1579 => x"000018b1",
			1580 => x"09015808",
			1581 => x"0410bb04",
			1582 => x"ff0b18d5",
			1583 => x"000018d5",
			1584 => x"0e075808",
			1585 => x"05070d04",
			1586 => x"008618d5",
			1587 => x"000018d5",
			1588 => x"000018d5",
			1589 => x"0100ca04",
			1590 => x"ff5718f9",
			1591 => x"0705ba0c",
			1592 => x"0e07dc08",
			1593 => x"0c058004",
			1594 => x"008018f9",
			1595 => x"000018f9",
			1596 => x"000018f9",
			1597 => x"000018f9",
			1598 => x"040c8504",
			1599 => x"fff1191d",
			1600 => x"0209ce04",
			1601 => x"0000191d",
			1602 => x"020a6308",
			1603 => x"04120c04",
			1604 => x"004e191d",
			1605 => x"0000191d",
			1606 => x"0000191d",
			1607 => x"040cbf04",
			1608 => x"00001941",
			1609 => x"020a200c",
			1610 => x"0209b104",
			1611 => x"00001941",
			1612 => x"04120c04",
			1613 => x"00371941",
			1614 => x"00001941",
			1615 => x"00001941",
			1616 => x"09015a08",
			1617 => x"0410bb04",
			1618 => x"ff35196d",
			1619 => x"0000196d",
			1620 => x"0e07dc0c",
			1621 => x"0209be04",
			1622 => x"0000196d",
			1623 => x"0c059b04",
			1624 => x"008c196d",
			1625 => x"0000196d",
			1626 => x"0000196d",
			1627 => x"0100ca08",
			1628 => x"0410bb04",
			1629 => x"ff8e1999",
			1630 => x"00001999",
			1631 => x"0e073b0c",
			1632 => x"07057504",
			1633 => x"00001999",
			1634 => x"06017304",
			1635 => x"00551999",
			1636 => x"00001999",
			1637 => x"00001999",
			1638 => x"040caf04",
			1639 => x"ff7019c5",
			1640 => x"0b060908",
			1641 => x"0100ca04",
			1642 => x"000019c5",
			1643 => x"008219c5",
			1644 => x"08033a04",
			1645 => x"000019c5",
			1646 => x"0f089c04",
			1647 => x"000019c5",
			1648 => x"ffcb19c5",
			1649 => x"0209c910",
			1650 => x"00041004",
			1651 => x"00001a01",
			1652 => x"06017408",
			1653 => x"0c058304",
			1654 => x"ff531a01",
			1655 => x"00001a01",
			1656 => x"00001a01",
			1657 => x"0f09150c",
			1658 => x"0a02f308",
			1659 => x"07055f04",
			1660 => x"00001a01",
			1661 => x"00a81a01",
			1662 => x"00001a01",
			1663 => x"00001a01",
			1664 => x"0209be08",
			1665 => x"08033904",
			1666 => x"00001a35",
			1667 => x"ff611a35",
			1668 => x"0f093310",
			1669 => x"07054904",
			1670 => x"00001a35",
			1671 => x"0a030408",
			1672 => x"0209c904",
			1673 => x"00001a35",
			1674 => x"00701a35",
			1675 => x"00001a35",
			1676 => x"00001a35",
			1677 => x"0100ad04",
			1678 => x"ffa51a61",
			1679 => x"0e078e10",
			1680 => x"0c059d0c",
			1681 => x"0f082204",
			1682 => x"00001a61",
			1683 => x"0c054604",
			1684 => x"00001a61",
			1685 => x"00211a61",
			1686 => x"00001a61",
			1687 => x"00001a61",
			1688 => x"02099a0c",
			1689 => x"07058c08",
			1690 => x"0c056304",
			1691 => x"fed51aa5",
			1692 => x"00001aa5",
			1693 => x"00001aa5",
			1694 => x"0f08a30c",
			1695 => x"08039608",
			1696 => x"0100bb04",
			1697 => x"00001aa5",
			1698 => x"00e61aa5",
			1699 => x"00001aa5",
			1700 => x"0e078e08",
			1701 => x"0100dc04",
			1702 => x"ffea1aa5",
			1703 => x"004c1aa5",
			1704 => x"ffa21aa5",
			1705 => x"02094304",
			1706 => x"fec11ae1",
			1707 => x"06016b0c",
			1708 => x"01009204",
			1709 => x"00001ae1",
			1710 => x"0e078e04",
			1711 => x"00db1ae1",
			1712 => x"00001ae1",
			1713 => x"09015a04",
			1714 => x"ff161ae1",
			1715 => x"0e075804",
			1716 => x"00771ae1",
			1717 => x"06016f04",
			1718 => x"00001ae1",
			1719 => x"ffaf1ae1",
			1720 => x"0209be0c",
			1721 => x"08033904",
			1722 => x"00001b25",
			1723 => x"0c058304",
			1724 => x"ff4c1b25",
			1725 => x"00001b25",
			1726 => x"0f093314",
			1727 => x"0c054804",
			1728 => x"00001b25",
			1729 => x"0c059c0c",
			1730 => x"06017808",
			1731 => x"01009204",
			1732 => x"00001b25",
			1733 => x"00ab1b25",
			1734 => x"00001b25",
			1735 => x"00001b25",
			1736 => x"00001b25",
			1737 => x"040ceb04",
			1738 => x"feeb1b69",
			1739 => x"0209ce10",
			1740 => x"08033f0c",
			1741 => x"0f08cd08",
			1742 => x"0100cf04",
			1743 => x"00001b69",
			1744 => x"003b1b69",
			1745 => x"00001b69",
			1746 => x"ff881b69",
			1747 => x"0601830c",
			1748 => x"0a030408",
			1749 => x"01009204",
			1750 => x"00001b69",
			1751 => x"00651b69",
			1752 => x"00001b69",
			1753 => x"00001b69",
			1754 => x"02099a0c",
			1755 => x"0c056308",
			1756 => x"07058c04",
			1757 => x"feaa1bb5",
			1758 => x"00001bb5",
			1759 => x"00001bb5",
			1760 => x"0f093318",
			1761 => x"0100ca10",
			1762 => x"0601660c",
			1763 => x"04128208",
			1764 => x"040fc604",
			1765 => x"00001bb5",
			1766 => x"006b1bb5",
			1767 => x"00001bb5",
			1768 => x"ffa51bb5",
			1769 => x"0209be04",
			1770 => x"00001bb5",
			1771 => x"00eb1bb5",
			1772 => x"ff721bb5",
			1773 => x"040d1b08",
			1774 => x"09015a04",
			1775 => x"feb71c11",
			1776 => x"00001c11",
			1777 => x"0209ce10",
			1778 => x"08033f0c",
			1779 => x"0f08cd08",
			1780 => x"0f084f04",
			1781 => x"00001c11",
			1782 => x"002a1c11",
			1783 => x"00001c11",
			1784 => x"ff731c11",
			1785 => x"0c05480c",
			1786 => x"0100dc08",
			1787 => x"0100b004",
			1788 => x"00001c11",
			1789 => x"ffd91c11",
			1790 => x"00001c11",
			1791 => x"0f093d08",
			1792 => x"0a030404",
			1793 => x"00b91c11",
			1794 => x"00001c11",
			1795 => x"00001c11",
			1796 => x"01009204",
			1797 => x"ff351c5d",
			1798 => x"0307c414",
			1799 => x"0c059d10",
			1800 => x"07054904",
			1801 => x"00001c5d",
			1802 => x"040c4404",
			1803 => x"00001c5d",
			1804 => x"0a030404",
			1805 => x"00c31c5d",
			1806 => x"00001c5d",
			1807 => x"00001c5d",
			1808 => x"09017a08",
			1809 => x"0d071604",
			1810 => x"00001c5d",
			1811 => x"ffc51c5d",
			1812 => x"0b064b04",
			1813 => x"00031c5d",
			1814 => x"00001c5d",
			1815 => x"0209b10c",
			1816 => x"09017a08",
			1817 => x"0c056304",
			1818 => x"fea91cb1",
			1819 => x"00001cb1",
			1820 => x"00001cb1",
			1821 => x"0f090d18",
			1822 => x"0209ce04",
			1823 => x"00001cb1",
			1824 => x"0c052804",
			1825 => x"00001cb1",
			1826 => x"0a03040c",
			1827 => x"0e075808",
			1828 => x"06017804",
			1829 => x"012d1cb1",
			1830 => x"00001cb1",
			1831 => x"00001cb1",
			1832 => x"00001cb1",
			1833 => x"0f093304",
			1834 => x"00001cb1",
			1835 => x"ff5a1cb1",
			1836 => x"0b06091c",
			1837 => x"0c050b04",
			1838 => x"00001cfd",
			1839 => x"0f08f014",
			1840 => x"02094304",
			1841 => x"00001cfd",
			1842 => x"04120c0c",
			1843 => x"0d066a04",
			1844 => x"00001cfd",
			1845 => x"020a5004",
			1846 => x"004f1cfd",
			1847 => x"00001cfd",
			1848 => x"00001cfd",
			1849 => x"00001cfd",
			1850 => x"0f089c04",
			1851 => x"00001cfd",
			1852 => x"0d071604",
			1853 => x"00001cfd",
			1854 => x"ffc11cfd",
			1855 => x"01009204",
			1856 => x"ff2e1d41",
			1857 => x"0f09151c",
			1858 => x"08034808",
			1859 => x"040c3204",
			1860 => x"00001d41",
			1861 => x"00911d41",
			1862 => x"0410bb0c",
			1863 => x"0b061908",
			1864 => x"020a2004",
			1865 => x"ff9e1d41",
			1866 => x"00001d41",
			1867 => x"00001d41",
			1868 => x"0b05b804",
			1869 => x"00021d41",
			1870 => x"00001d41",
			1871 => x"ffee1d41",
			1872 => x"0209b114",
			1873 => x"0100cd04",
			1874 => x"fe761dad",
			1875 => x"0b06060c",
			1876 => x"0209ab08",
			1877 => x"0c050c04",
			1878 => x"00001dad",
			1879 => x"00fc1dad",
			1880 => x"00001dad",
			1881 => x"fe891dad",
			1882 => x"06016b10",
			1883 => x"01009204",
			1884 => x"00001dad",
			1885 => x"03089d08",
			1886 => x"0c054304",
			1887 => x"00001dad",
			1888 => x"02601dad",
			1889 => x"00001dad",
			1890 => x"03087510",
			1891 => x"09015804",
			1892 => x"ff141dad",
			1893 => x"0209c108",
			1894 => x"0d071604",
			1895 => x"00001dad",
			1896 => x"ffb51dad",
			1897 => x"01521dad",
			1898 => x"fec91dad",
			1899 => x"07054908",
			1900 => x"0c054304",
			1901 => x"ff3e1e09",
			1902 => x"00001e09",
			1903 => x"0307c418",
			1904 => x"0c059d14",
			1905 => x"0900e004",
			1906 => x"00001e09",
			1907 => x"040c4404",
			1908 => x"00001e09",
			1909 => x"00055408",
			1910 => x"020a5004",
			1911 => x"00b21e09",
			1912 => x"00001e09",
			1913 => x"00001e09",
			1914 => x"00001e09",
			1915 => x"0b060904",
			1916 => x"00001e09",
			1917 => x"06017308",
			1918 => x"09018b04",
			1919 => x"ffc51e09",
			1920 => x"00001e09",
			1921 => x"00001e09",
			1922 => x"040caf04",
			1923 => x"fe6d1e65",
			1924 => x"0100ca0c",
			1925 => x"0100ad04",
			1926 => x"fe6b1e65",
			1927 => x"06017004",
			1928 => x"02301e65",
			1929 => x"fe7c1e65",
			1930 => x"0e075810",
			1931 => x"00046b04",
			1932 => x"01ab1e65",
			1933 => x"020a0604",
			1934 => x"ffa51e65",
			1935 => x"020a3a04",
			1936 => x"025c1e65",
			1937 => x"002b1e65",
			1938 => x"08033704",
			1939 => x"01291e65",
			1940 => x"0100ed04",
			1941 => x"fe1c1e65",
			1942 => x"0100f804",
			1943 => x"00141e65",
			1944 => x"ff121e65",
			1945 => x"040cbf08",
			1946 => x"040cb604",
			1947 => x"fe931ee1",
			1948 => x"00001ee1",
			1949 => x"0209c91c",
			1950 => x"08033a0c",
			1951 => x"0100cf04",
			1952 => x"00001ee1",
			1953 => x"0f08b804",
			1954 => x"00af1ee1",
			1955 => x"00001ee1",
			1956 => x"0601740c",
			1957 => x"0b061b08",
			1958 => x"0a028804",
			1959 => x"00001ee1",
			1960 => x"fef21ee1",
			1961 => x"00001ee1",
			1962 => x"00001ee1",
			1963 => x"0d06c70c",
			1964 => x"0a030408",
			1965 => x"0c052804",
			1966 => x"00001ee1",
			1967 => x"01c81ee1",
			1968 => x"00001ee1",
			1969 => x"0100dc08",
			1970 => x"0e071504",
			1971 => x"00001ee1",
			1972 => x"ff451ee1",
			1973 => x"0d078804",
			1974 => x"00ee1ee1",
			1975 => x"00001ee1",
			1976 => x"040cbf04",
			1977 => x"fed11f3d",
			1978 => x"0e07581c",
			1979 => x"0100ca18",
			1980 => x"0410bb08",
			1981 => x"0c056304",
			1982 => x"ff7a1f3d",
			1983 => x"00001f3d",
			1984 => x"0a03040c",
			1985 => x"0d069408",
			1986 => x"0f073b04",
			1987 => x"00001f3d",
			1988 => x"004c1f3d",
			1989 => x"00001f3d",
			1990 => x"00001f3d",
			1991 => x"00e51f3d",
			1992 => x"0c056508",
			1993 => x"0c052e04",
			1994 => x"00001f3d",
			1995 => x"ff2c1f3d",
			1996 => x"0f093d04",
			1997 => x"002d1f3d",
			1998 => x"00001f3d",
			1999 => x"02096c0c",
			2000 => x"02094904",
			2001 => x"fe6d1fc9",
			2002 => x"02094d04",
			2003 => x"00001fc9",
			2004 => x"ff981fc9",
			2005 => x"0c059d2c",
			2006 => x"0209ce18",
			2007 => x"08033a0c",
			2008 => x"0e078e08",
			2009 => x"0c052504",
			2010 => x"00001fc9",
			2011 => x"01621fc9",
			2012 => x"ff5f1fc9",
			2013 => x"0c056308",
			2014 => x"0209c104",
			2015 => x"fe8d1fc9",
			2016 => x"00001fc9",
			2017 => x"00001fc9",
			2018 => x"0c052808",
			2019 => x"0a02b104",
			2020 => x"00001fc9",
			2021 => x"ff811fc9",
			2022 => x"0a02f308",
			2023 => x"03087504",
			2024 => x"01b71fc9",
			2025 => x"00001fc9",
			2026 => x"ffda1fc9",
			2027 => x"0705e80c",
			2028 => x"0b061904",
			2029 => x"ff661fc9",
			2030 => x"0e082c04",
			2031 => x"001c1fc9",
			2032 => x"00001fc9",
			2033 => x"fe811fc9",
			2034 => x"09015828",
			2035 => x"0100d624",
			2036 => x"0100ca18",
			2037 => x"0209c104",
			2038 => x"fe612045",
			2039 => x"0209c908",
			2040 => x"01004104",
			2041 => x"ff682045",
			2042 => x"0b392045",
			2043 => x"0b05b408",
			2044 => x"0c054304",
			2045 => x"fe902045",
			2046 => x"187f2045",
			2047 => x"fe642045",
			2048 => x"0d06d208",
			2049 => x"0003f204",
			2050 => x"ff222045",
			2051 => x"08432045",
			2052 => x"fe552045",
			2053 => x"fc552045",
			2054 => x"0e07dc14",
			2055 => x"09018310",
			2056 => x"0e073b08",
			2057 => x"0100d804",
			2058 => x"02c72045",
			2059 => x"01e22045",
			2060 => x"0506e204",
			2061 => x"01c92045",
			2062 => x"fe332045",
			2063 => x"05822045",
			2064 => x"fe622045",
			2065 => x"0100b004",
			2066 => x"fe6c20b9",
			2067 => x"0c059b2c",
			2068 => x"0e07581c",
			2069 => x"0d06f90c",
			2070 => x"0f082b04",
			2071 => x"000020b9",
			2072 => x"0b05a704",
			2073 => x"000020b9",
			2074 => x"01dc20b9",
			2075 => x"040e6308",
			2076 => x"0003c404",
			2077 => x"000020b9",
			2078 => x"016b20b9",
			2079 => x"0f08bf04",
			2080 => x"fedc20b9",
			2081 => x"000020b9",
			2082 => x"0c056308",
			2083 => x"0a028d04",
			2084 => x"000020b9",
			2085 => x"fe3920b9",
			2086 => x"0e07dc04",
			2087 => x"015320b9",
			2088 => x"000020b9",
			2089 => x"05070d04",
			2090 => x"000020b9",
			2091 => x"0c059c04",
			2092 => x"000020b9",
			2093 => x"fe7d20b9",
			2094 => x"02096c0c",
			2095 => x"02094904",
			2096 => x"fe672135",
			2097 => x"02094d04",
			2098 => x"00002135",
			2099 => x"ff022135",
			2100 => x"0c05b42c",
			2101 => x"0e075814",
			2102 => x"09011304",
			2103 => x"fea02135",
			2104 => x"0a02e40c",
			2105 => x"0c059c08",
			2106 => x"0004c904",
			2107 => x"016e2135",
			2108 => x"02e42135",
			2109 => x"00002135",
			2110 => x"ff262135",
			2111 => x"08033908",
			2112 => x"040c3204",
			2113 => x"ff002135",
			2114 => x"01302135",
			2115 => x"0209ce04",
			2116 => x"fdba2135",
			2117 => x"0100e804",
			2118 => x"fefa2135",
			2119 => x"09019604",
			2120 => x"00dd2135",
			2121 => x"00002135",
			2122 => x"0705d004",
			2123 => x"00002135",
			2124 => x"fe622135",
			2125 => x"02096004",
			2126 => x"fe6421a9",
			2127 => x"0c059b24",
			2128 => x"0100b40c",
			2129 => x"0c054804",
			2130 => x"fe7121a9",
			2131 => x"07057304",
			2132 => x"05ee21a9",
			2133 => x"fecc21a9",
			2134 => x"0e067104",
			2135 => x"0bdf21a9",
			2136 => x"0803740c",
			2137 => x"0e07dc08",
			2138 => x"0e078e04",
			2139 => x"01b921a9",
			2140 => x"06f321a9",
			2141 => x"fe9221a9",
			2142 => x"06017c04",
			2143 => x"fce821a9",
			2144 => x"feca21a9",
			2145 => x"0705d110",
			2146 => x"0b061908",
			2147 => x"0705ce04",
			2148 => x"fe3921a9",
			2149 => x"000021a9",
			2150 => x"0307f404",
			2151 => x"019421a9",
			2152 => x"ff3b21a9",
			2153 => x"fe6121a9",
			2154 => x"02096008",
			2155 => x"02094304",
			2156 => x"fe632215",
			2157 => x"fed92215",
			2158 => x"0e07dc2c",
			2159 => x"0100ad0c",
			2160 => x"01009204",
			2161 => x"fe6c2215",
			2162 => x"01009304",
			2163 => x"07c62215",
			2164 => x"fe962215",
			2165 => x"0e065a08",
			2166 => x"0803c704",
			2167 => x"092d2215",
			2168 => x"02a62215",
			2169 => x"08037e10",
			2170 => x"0100d408",
			2171 => x"0f08cd04",
			2172 => x"041b2215",
			2173 => x"ff812215",
			2174 => x"0100dc04",
			2175 => x"00222215",
			2176 => x"01b32215",
			2177 => x"06017304",
			2178 => x"00002215",
			2179 => x"fdda2215",
			2180 => x"fe642215",
			2181 => x"02096c08",
			2182 => x"02096604",
			2183 => x"fe782289",
			2184 => x"00002289",
			2185 => x"0e055208",
			2186 => x"03061104",
			2187 => x"00002289",
			2188 => x"12f62289",
			2189 => x"06016a0c",
			2190 => x"0b062a08",
			2191 => x"0100ad04",
			2192 => x"00002289",
			2193 => x"01f62289",
			2194 => x"00002289",
			2195 => x"0e07dc1c",
			2196 => x"0100de10",
			2197 => x"0209dd08",
			2198 => x"00042904",
			2199 => x"00002289",
			2200 => x"feb62289",
			2201 => x"09015504",
			2202 => x"ff832289",
			2203 => x"00882289",
			2204 => x"0209c108",
			2205 => x"0307c404",
			2206 => x"00952289",
			2207 => x"ffa02289",
			2208 => x"01662289",
			2209 => x"fea32289",
			2210 => x"0209570c",
			2211 => x"02094304",
			2212 => x"fe65231d",
			2213 => x"02094d04",
			2214 => x"ffbf231d",
			2215 => x"fed0231d",
			2216 => x"0c059d30",
			2217 => x"09010f04",
			2218 => x"fe82231d",
			2219 => x"0e075810",
			2220 => x"0e060f04",
			2221 => x"05eb231d",
			2222 => x"08039308",
			2223 => x"0506d204",
			2224 => x"01cd231d",
			2225 => x"00f7231d",
			2226 => x"fec1231d",
			2227 => x"0803390c",
			2228 => x"0e07dc08",
			2229 => x"0c056604",
			2230 => x"00ce231d",
			2231 => x"02b1231d",
			2232 => x"feee231d",
			2233 => x"0209e808",
			2234 => x"05067e04",
			2235 => x"ffad231d",
			2236 => x"fc83231d",
			2237 => x"0f096804",
			2238 => x"00ab231d",
			2239 => x"ff1d231d",
			2240 => x"0705d10c",
			2241 => x"0b061904",
			2242 => x"febd231d",
			2243 => x"0307f404",
			2244 => x"0141231d",
			2245 => x"0000231d",
			2246 => x"fe60231d",
			2247 => x"02096004",
			2248 => x"fe6623ab",
			2249 => x"0c059d34",
			2250 => x"0100ad04",
			2251 => x"fe7723ab",
			2252 => x"0e075818",
			2253 => x"0100d40c",
			2254 => x"0803b408",
			2255 => x"0b05c704",
			2256 => x"054d23ab",
			2257 => x"032423ab",
			2258 => x"ff7023ab",
			2259 => x"0100da08",
			2260 => x"0d06f904",
			2261 => x"017823ab",
			2262 => x"fec123ab",
			2263 => x"01b423ab",
			2264 => x"0100e80c",
			2265 => x"040d8808",
			2266 => x"040c5204",
			2267 => x"fee323ab",
			2268 => x"000023ab",
			2269 => x"fa3a23ab",
			2270 => x"0e07dc08",
			2271 => x"0209ce04",
			2272 => x"00ba23ab",
			2273 => x"03b723ab",
			2274 => x"feb423ab",
			2275 => x"0705d10c",
			2276 => x"0e073b08",
			2277 => x"0506a704",
			2278 => x"ff7723ab",
			2279 => x"010c23ab",
			2280 => x"fe4c23ab",
			2281 => x"fe6523ab",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(726, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(1470, initial_addr_3'length));
	end generate gen_rom_12;

	gen_rom_13: if SELECT_ROM = 13 generate
		bank <= (
			0 => x"00000005",
			1 => x"00000009",
			2 => x"0000000d",
			3 => x"00000011",
			4 => x"00000015",
			5 => x"00000019",
			6 => x"0000001d",
			7 => x"00000021",
			8 => x"00000025",
			9 => x"00000029",
			10 => x"040c2404",
			11 => x"ffe20035",
			12 => x"00000035",
			13 => x"0100bd04",
			14 => x"00000049",
			15 => x"0100f304",
			16 => x"000a0049",
			17 => x"00000049",
			18 => x"0c054808",
			19 => x"0c04b204",
			20 => x"0000005d",
			21 => x"001e005d",
			22 => x"0000005d",
			23 => x"0900b704",
			24 => x"00000071",
			25 => x"09018704",
			26 => x"00100071",
			27 => x"00000071",
			28 => x"0307f408",
			29 => x"04100804",
			30 => x"ffc60085",
			31 => x"00000085",
			32 => x"00000085",
			33 => x"0f08dd08",
			34 => x"0f070104",
			35 => x"000000a1",
			36 => x"002700a1",
			37 => x"0f0abc04",
			38 => x"ffd900a1",
			39 => x"000000a1",
			40 => x"06016b08",
			41 => x"00040304",
			42 => x"000000bd",
			43 => x"ffdf00bd",
			44 => x"06019004",
			45 => x"000900bd",
			46 => x"000000bd",
			47 => x"02086004",
			48 => x"000000d9",
			49 => x"040e2308",
			50 => x"0f0abc04",
			51 => x"ff6a00d9",
			52 => x"000000d9",
			53 => x"000000d9",
			54 => x"0506e20c",
			55 => x"00040704",
			56 => x"000000f5",
			57 => x"0005b804",
			58 => x"ffd700f5",
			59 => x"000000f5",
			60 => x"000000f5",
			61 => x"0d07300c",
			62 => x"00040704",
			63 => x"00000111",
			64 => x"0005b804",
			65 => x"ffbf0111",
			66 => x"00000111",
			67 => x"00000111",
			68 => x"00046704",
			69 => x"0000012d",
			70 => x"01006704",
			71 => x"0000012d",
			72 => x"0100df04",
			73 => x"002f012d",
			74 => x"0000012d",
			75 => x"0306ff08",
			76 => x"06017304",
			77 => x"ffe10151",
			78 => x"00000151",
			79 => x"09018708",
			80 => x"09010604",
			81 => x"00000151",
			82 => x"00130151",
			83 => x"00000151",
			84 => x"06016b08",
			85 => x"02086004",
			86 => x"0000017d",
			87 => x"ffc0017d",
			88 => x"040dca08",
			89 => x"040ae204",
			90 => x"0000017d",
			91 => x"fff4017d",
			92 => x"0413e904",
			93 => x"0025017d",
			94 => x"0000017d",
			95 => x"0c050c0c",
			96 => x"07050104",
			97 => x"000001a9",
			98 => x"0d05f704",
			99 => x"000001a9",
			100 => x"001201a9",
			101 => x"0d075508",
			102 => x"07054904",
			103 => x"000001a9",
			104 => x"ffd801a9",
			105 => x"000001a9",
			106 => x"07058c10",
			107 => x"07050404",
			108 => x"000001cd",
			109 => x"0c052e08",
			110 => x"0c04b204",
			111 => x"000001cd",
			112 => x"003301cd",
			113 => x"000001cd",
			114 => x"fff801cd",
			115 => x"0506e210",
			116 => x"040ae204",
			117 => x"000001f1",
			118 => x"04120c08",
			119 => x"02086004",
			120 => x"000001f1",
			121 => x"ffac01f1",
			122 => x"000001f1",
			123 => x"000001f1",
			124 => x"0506e204",
			125 => x"00000215",
			126 => x"0901a10c",
			127 => x"09012d04",
			128 => x"00000215",
			129 => x"0d086d04",
			130 => x"003c0215",
			131 => x"00000215",
			132 => x"00000215",
			133 => x"00046704",
			134 => x"00000239",
			135 => x"01006704",
			136 => x"00000239",
			137 => x"0100df08",
			138 => x"0803dc04",
			139 => x"003c0239",
			140 => x"00000239",
			141 => x"00000239",
			142 => x"02086004",
			143 => x"00000265",
			144 => x"0d073008",
			145 => x"0005b804",
			146 => x"ffa80265",
			147 => x"00000265",
			148 => x"0705fd04",
			149 => x"000b0265",
			150 => x"07069b04",
			151 => x"ffe50265",
			152 => x"00000265",
			153 => x"0004670c",
			154 => x"00040304",
			155 => x"00000299",
			156 => x"040da904",
			157 => x"ffd60299",
			158 => x"00000299",
			159 => x"0803820c",
			160 => x"07050404",
			161 => x"00000299",
			162 => x"0705bb04",
			163 => x"00410299",
			164 => x"00000299",
			165 => x"00000299",
			166 => x"0004140c",
			167 => x"0a028d04",
			168 => x"000002cd",
			169 => x"0a029b04",
			170 => x"001102cd",
			171 => x"000002cd",
			172 => x"0f0a420c",
			173 => x"0a028504",
			174 => x"000002cd",
			175 => x"0005b804",
			176 => x"ffe102cd",
			177 => x"000002cd",
			178 => x"000002cd",
			179 => x"0a02920c",
			180 => x"0a028d04",
			181 => x"00000301",
			182 => x"0c050704",
			183 => x"00000301",
			184 => x"004d0301",
			185 => x"0b064b0c",
			186 => x"0c04e904",
			187 => x"00000301",
			188 => x"04120c04",
			189 => x"ffc30301",
			190 => x"00000301",
			191 => x"00000301",
			192 => x"0306ff08",
			193 => x"06017304",
			194 => x"ffdb0335",
			195 => x"00000335",
			196 => x"0601a310",
			197 => x"0100fa0c",
			198 => x"09010604",
			199 => x"00000335",
			200 => x"06016704",
			201 => x"00000335",
			202 => x"006b0335",
			203 => x"00000335",
			204 => x"00000335",
			205 => x"040c660c",
			206 => x"040ae204",
			207 => x"00000371",
			208 => x"06019604",
			209 => x"ffa20371",
			210 => x"00000371",
			211 => x"06018110",
			212 => x"01006704",
			213 => x"00000371",
			214 => x"0100de08",
			215 => x"0410bb04",
			216 => x"005b0371",
			217 => x"00000371",
			218 => x"00000371",
			219 => x"00000371",
			220 => x"0506e20c",
			221 => x"040ae204",
			222 => x"000003ad",
			223 => x"04114904",
			224 => x"ffe803ad",
			225 => x"000003ad",
			226 => x"0c05dc10",
			227 => x"0100fa0c",
			228 => x"0e071504",
			229 => x"000003ad",
			230 => x"0a028d04",
			231 => x"000003ad",
			232 => x"007103ad",
			233 => x"000003ad",
			234 => x"000003ad",
			235 => x"0705cf1c",
			236 => x"0b05f810",
			237 => x"040ae204",
			238 => x"000003f9",
			239 => x"04100808",
			240 => x"03061904",
			241 => x"000003f9",
			242 => x"ff9a03f9",
			243 => x"000003f9",
			244 => x"0d070804",
			245 => x"000003f9",
			246 => x"040d1b04",
			247 => x"000003f9",
			248 => x"005e03f9",
			249 => x"030a5c08",
			250 => x"0c057d04",
			251 => x"000003f9",
			252 => x"ff8603f9",
			253 => x"000003f9",
			254 => x"0f09b11c",
			255 => x"0d070808",
			256 => x"0e06f704",
			257 => x"fff6043d",
			258 => x"0000043d",
			259 => x"0b05f804",
			260 => x"0000043d",
			261 => x"0c059e0c",
			262 => x"0100ff08",
			263 => x"0e089604",
			264 => x"0054043d",
			265 => x"0000043d",
			266 => x"0000043d",
			267 => x"0000043d",
			268 => x"0003fb04",
			269 => x"0000043d",
			270 => x"ff89043d",
			271 => x"00040714",
			272 => x"0003f704",
			273 => x"00000489",
			274 => x"05061504",
			275 => x"00000489",
			276 => x"08033108",
			277 => x"040cbf04",
			278 => x"00610489",
			279 => x"00000489",
			280 => x"00000489",
			281 => x"0f074904",
			282 => x"00000489",
			283 => x"040e230c",
			284 => x"02088304",
			285 => x"00000489",
			286 => x"0e097704",
			287 => x"ff880489",
			288 => x"00000489",
			289 => x"00000489",
			290 => x"0d075518",
			291 => x"02088304",
			292 => x"000004bd",
			293 => x"0005b810",
			294 => x"0100eb0c",
			295 => x"0004e908",
			296 => x"0307f404",
			297 => x"ffa204bd",
			298 => x"000004bd",
			299 => x"000004bd",
			300 => x"000004bd",
			301 => x"000004bd",
			302 => x"000004bd",
			303 => x"00040718",
			304 => x"08031d04",
			305 => x"00000509",
			306 => x"0901b810",
			307 => x"0d063804",
			308 => x"00000509",
			309 => x"08033108",
			310 => x"040adc04",
			311 => x"00000509",
			312 => x"00ab0509",
			313 => x"00000509",
			314 => x"00000509",
			315 => x"09011b0c",
			316 => x"04120c08",
			317 => x"0f079d04",
			318 => x"00000509",
			319 => x"ff7a0509",
			320 => x"00000509",
			321 => x"00000509",
			322 => x"09014120",
			323 => x"02089114",
			324 => x"03060104",
			325 => x"0000055d",
			326 => x"0b05650c",
			327 => x"0b053504",
			328 => x"0000055d",
			329 => x"03067804",
			330 => x"002a055d",
			331 => x"0000055d",
			332 => x"0000055d",
			333 => x"04120c08",
			334 => x"0f073b04",
			335 => x"0000055d",
			336 => x"ff70055d",
			337 => x"0000055d",
			338 => x"0100e208",
			339 => x"09015304",
			340 => x"0000055d",
			341 => x"002e055d",
			342 => x"0000055d",
			343 => x"0c050c18",
			344 => x"0b053504",
			345 => x"000005b1",
			346 => x"08032504",
			347 => x"000005b1",
			348 => x"0208dd0c",
			349 => x"07050404",
			350 => x"000005b1",
			351 => x"0d05f704",
			352 => x"000005b1",
			353 => x"006005b1",
			354 => x"000005b1",
			355 => x"0f084f04",
			356 => x"000005b1",
			357 => x"030a5c0c",
			358 => x"0209c904",
			359 => x"000005b1",
			360 => x"07058b04",
			361 => x"000005b1",
			362 => x"ffad05b1",
			363 => x"000005b1",
			364 => x"0c05281c",
			365 => x"0c04d004",
			366 => x"000005fd",
			367 => x"00040204",
			368 => x"000005fd",
			369 => x"0e053404",
			370 => x"000005fd",
			371 => x"06014604",
			372 => x"000005fd",
			373 => x"020a8608",
			374 => x"03087504",
			375 => x"005e05fd",
			376 => x"000005fd",
			377 => x"000005fd",
			378 => x"020a6308",
			379 => x"0209c904",
			380 => x"000005fd",
			381 => x"ffc905fd",
			382 => x"000005fd",
			383 => x"0f08dd1c",
			384 => x"07050404",
			385 => x"00000641",
			386 => x"0c056514",
			387 => x"020a0610",
			388 => x"0601740c",
			389 => x"06014104",
			390 => x"00000641",
			391 => x"0f06e304",
			392 => x"00000641",
			393 => x"00680641",
			394 => x"00000641",
			395 => x"00000641",
			396 => x"00000641",
			397 => x"0c050b04",
			398 => x"00000641",
			399 => x"ffc90641",
			400 => x"09012008",
			401 => x"0005b804",
			402 => x"ffbf0685",
			403 => x"00000685",
			404 => x"0705fd18",
			405 => x"0d071604",
			406 => x"00000685",
			407 => x"09018710",
			408 => x"0100c204",
			409 => x"00000685",
			410 => x"0f08a304",
			411 => x"00000685",
			412 => x"0a028d04",
			413 => x"00000685",
			414 => x"006e0685",
			415 => x"00000685",
			416 => x"00000685",
			417 => x"09010608",
			418 => x"040fc604",
			419 => x"ff9d06d9",
			420 => x"000006d9",
			421 => x"0100d018",
			422 => x"06016b04",
			423 => x"000006d9",
			424 => x"03087510",
			425 => x"0c050a04",
			426 => x"000006d9",
			427 => x"00040304",
			428 => x"000006d9",
			429 => x"0803e604",
			430 => x"00dd06d9",
			431 => x"000006d9",
			432 => x"000006d9",
			433 => x"0f08c604",
			434 => x"000006d9",
			435 => x"06018804",
			436 => x"ffe106d9",
			437 => x"000006d9",
			438 => x"0c05281c",
			439 => x"0d05f704",
			440 => x"0000072d",
			441 => x"08032504",
			442 => x"0000072d",
			443 => x"0f08d410",
			444 => x"06017f0c",
			445 => x"00040204",
			446 => x"0000072d",
			447 => x"0c04b204",
			448 => x"0000072d",
			449 => x"0071072d",
			450 => x"0000072d",
			451 => x"0000072d",
			452 => x"0209c104",
			453 => x"0000072d",
			454 => x"00040704",
			455 => x"0000072d",
			456 => x"0005b804",
			457 => x"ffbc072d",
			458 => x"0000072d",
			459 => x"0c050c1c",
			460 => x"0c04d004",
			461 => x"00000781",
			462 => x"08032504",
			463 => x"00000781",
			464 => x"0208dd10",
			465 => x"0900b704",
			466 => x"00000781",
			467 => x"0d05f704",
			468 => x"00000781",
			469 => x"07050404",
			470 => x"00000781",
			471 => x"006c0781",
			472 => x"00000781",
			473 => x"0f084f04",
			474 => x"00000781",
			475 => x"00040304",
			476 => x"00000781",
			477 => x"07054904",
			478 => x"00000781",
			479 => x"ffb70781",
			480 => x"0900b704",
			481 => x"000007bd",
			482 => x"0100fa18",
			483 => x"0b053504",
			484 => x"000007bd",
			485 => x"08031d04",
			486 => x"000007bd",
			487 => x"0601990c",
			488 => x"0705e608",
			489 => x"0003f704",
			490 => x"000007bd",
			491 => x"005b07bd",
			492 => x"000007bd",
			493 => x"000007bd",
			494 => x"000007bd",
			495 => x"0e055204",
			496 => x"000007f9",
			497 => x"0c056518",
			498 => x"0a028d04",
			499 => x"000007f9",
			500 => x"0900b704",
			501 => x"000007f9",
			502 => x"0c04d004",
			503 => x"000007f9",
			504 => x"09018308",
			505 => x"0e087804",
			506 => x"004807f9",
			507 => x"000007f9",
			508 => x"000007f9",
			509 => x"000007f9",
			510 => x"0506b918",
			511 => x"02089110",
			512 => x"0305b004",
			513 => x"0000085d",
			514 => x"02081b04",
			515 => x"0000085d",
			516 => x"0f079d04",
			517 => x"0058085d",
			518 => x"0000085d",
			519 => x"0004e904",
			520 => x"ff2b085d",
			521 => x"0000085d",
			522 => x"0100f318",
			523 => x"0c052704",
			524 => x"0000085d",
			525 => x"020b2c10",
			526 => x"0003e104",
			527 => x"0000085d",
			528 => x"09010f04",
			529 => x"0000085d",
			530 => x"0d06f904",
			531 => x"0000085d",
			532 => x"00a4085d",
			533 => x"0000085d",
			534 => x"0000085d",
			535 => x"0100bc1c",
			536 => x"0f085c18",
			537 => x"0e055204",
			538 => x"000008b9",
			539 => x"07050404",
			540 => x"000008b9",
			541 => x"0c05460c",
			542 => x"0b053504",
			543 => x"000008b9",
			544 => x"0c04d004",
			545 => x"000008b9",
			546 => x"005d08b9",
			547 => x"000008b9",
			548 => x"ffba08b9",
			549 => x"0100de10",
			550 => x"00044e04",
			551 => x"000008b9",
			552 => x"07065608",
			553 => x"0a02b004",
			554 => x"000008b9",
			555 => x"009e08b9",
			556 => x"000008b9",
			557 => x"000008b9",
			558 => x"0209ce1c",
			559 => x"0b053504",
			560 => x"00000915",
			561 => x"0c056614",
			562 => x"00040204",
			563 => x"00000915",
			564 => x"08032504",
			565 => x"00000915",
			566 => x"0c04d004",
			567 => x"00000915",
			568 => x"07050404",
			569 => x"00000915",
			570 => x"00540915",
			571 => x"00000915",
			572 => x"00040304",
			573 => x"00000915",
			574 => x"0c052804",
			575 => x"00000915",
			576 => x"07054904",
			577 => x"00000915",
			578 => x"0005b804",
			579 => x"ffb40915",
			580 => x"00000915",
			581 => x"07058c2c",
			582 => x"01009214",
			583 => x"040cce04",
			584 => x"ff860989",
			585 => x"0e057f0c",
			586 => x"07050104",
			587 => x"00000989",
			588 => x"03055f04",
			589 => x"00000989",
			590 => x"00590989",
			591 => x"00000989",
			592 => x"06018e14",
			593 => x"06016604",
			594 => x"00000989",
			595 => x"0c050a04",
			596 => x"00000989",
			597 => x"00040304",
			598 => x"00000989",
			599 => x"0a028d04",
			600 => x"00000989",
			601 => x"00ce0989",
			602 => x"00000989",
			603 => x"0307f40c",
			604 => x"0b05e504",
			605 => x"00000989",
			606 => x"0209b104",
			607 => x"00000989",
			608 => x"ff7d0989",
			609 => x"00000989",
			610 => x"040c7f18",
			611 => x"0f077b10",
			612 => x"0e057104",
			613 => x"00000a1d",
			614 => x"0b053504",
			615 => x"00000a1d",
			616 => x"0b055204",
			617 => x"00460a1d",
			618 => x"00000a1d",
			619 => x"05084d04",
			620 => x"ff2c0a1d",
			621 => x"00000a1d",
			622 => x"08036814",
			623 => x"09018710",
			624 => x"0a028d04",
			625 => x"00000a1d",
			626 => x"00047908",
			627 => x"01006704",
			628 => x"00000a1d",
			629 => x"00d20a1d",
			630 => x"00000a1d",
			631 => x"00000a1d",
			632 => x"06018818",
			633 => x"0d06c70c",
			634 => x"04114908",
			635 => x"0305e904",
			636 => x"00000a1d",
			637 => x"ffc00a1d",
			638 => x"00000a1d",
			639 => x"040eab04",
			640 => x"00000a1d",
			641 => x"01009304",
			642 => x"00000a1d",
			643 => x"00680a1d",
			644 => x"0d07ee04",
			645 => x"ff970a1d",
			646 => x"00000a1d",
			647 => x"0d05f704",
			648 => x"ffcd0a79",
			649 => x"07058c18",
			650 => x"00040204",
			651 => x"00000a79",
			652 => x"03087510",
			653 => x"0900b704",
			654 => x"00000a79",
			655 => x"0b053504",
			656 => x"00000a79",
			657 => x"0c056304",
			658 => x"00b00a79",
			659 => x"00000a79",
			660 => x"00000a79",
			661 => x"0209c904",
			662 => x"00000a79",
			663 => x"0100c904",
			664 => x"00000a79",
			665 => x"00040704",
			666 => x"00000a79",
			667 => x"0004f704",
			668 => x"ff910a79",
			669 => x"00000a79",
			670 => x"0d061108",
			671 => x"04100804",
			672 => x"fef90af5",
			673 => x"00000af5",
			674 => x"0208dd14",
			675 => x"07051f10",
			676 => x"0c04ed04",
			677 => x"00000af5",
			678 => x"0b056908",
			679 => x"00040204",
			680 => x"00000af5",
			681 => x"01710af5",
			682 => x"00000af5",
			683 => x"00000af5",
			684 => x"0100bb10",
			685 => x"040fc608",
			686 => x"0e060004",
			687 => x"00000af5",
			688 => x"ff290af5",
			689 => x"06016a04",
			690 => x"00000af5",
			691 => x"00400af5",
			692 => x"0a028e04",
			693 => x"ffc10af5",
			694 => x"030a690c",
			695 => x"0b05e804",
			696 => x"00000af5",
			697 => x"0100fa04",
			698 => x"00d50af5",
			699 => x"00000af5",
			700 => x"00000af5",
			701 => x"0d05f704",
			702 => x"fe6a0b51",
			703 => x"0c059e1c",
			704 => x"0a036318",
			705 => x"0003f704",
			706 => x"fea30b51",
			707 => x"02086f04",
			708 => x"04830b51",
			709 => x"05060608",
			710 => x"03060104",
			711 => x"00740b51",
			712 => x"fe9a0b51",
			713 => x"06016304",
			714 => x"ffb70b51",
			715 => x"011f0b51",
			716 => x"fe8b0b51",
			717 => x"020b1c04",
			718 => x"fe650b51",
			719 => x"0f0b1c08",
			720 => x"040ce104",
			721 => x"01740b51",
			722 => x"ff780b51",
			723 => x"fe830b51",
			724 => x"040d1b24",
			725 => x"040c7f0c",
			726 => x"020b1c04",
			727 => x"fe6d0bf5",
			728 => x"020b1f04",
			729 => x"00ee0bf5",
			730 => x"fe700bf5",
			731 => x"08034114",
			732 => x"08032c0c",
			733 => x"040caf08",
			734 => x"040c9a04",
			735 => x"00000bf5",
			736 => x"01730bf5",
			737 => x"fed00bf5",
			738 => x"0a02a104",
			739 => x"04670bf5",
			740 => x"ff700bf5",
			741 => x"fe680bf5",
			742 => x"0100760c",
			743 => x"020a5008",
			744 => x"020a3a04",
			745 => x"fe6a0bf5",
			746 => x"fca20bf5",
			747 => x"00510bf5",
			748 => x"020ab518",
			749 => x"0208f904",
			750 => x"050a0bf5",
			751 => x"0e07580c",
			752 => x"0100de08",
			753 => x"0505f604",
			754 => x"fe520bf5",
			755 => x"01ae0bf5",
			756 => x"fe950bf5",
			757 => x"0100e804",
			758 => x"061c0bf5",
			759 => x"01140bf5",
			760 => x"08038108",
			761 => x"0a02cc04",
			762 => x"ff6a0bf5",
			763 => x"00b70bf5",
			764 => x"fe620bf5",
			765 => x"0f08dd34",
			766 => x"07050408",
			767 => x"0a034104",
			768 => x"ff670c69",
			769 => x"00000c69",
			770 => x"07051a14",
			771 => x"0208dd10",
			772 => x"0e050004",
			773 => x"00000c69",
			774 => x"0a028304",
			775 => x"00000c69",
			776 => x"0d05f704",
			777 => x"00000c69",
			778 => x"01020c69",
			779 => x"00000c69",
			780 => x"040d4208",
			781 => x"02088304",
			782 => x"00000c69",
			783 => x"ffa70c69",
			784 => x"0e05e004",
			785 => x"00000c69",
			786 => x"0705ce08",
			787 => x"08033a04",
			788 => x"00000c69",
			789 => x"00960c69",
			790 => x"00000c69",
			791 => x"0e086804",
			792 => x"ff360c69",
			793 => x"00000c69",
			794 => x"040d1b18",
			795 => x"040c6604",
			796 => x"fe710cdd",
			797 => x"08036610",
			798 => x"040c6c04",
			799 => x"06790cdd",
			800 => x"03087504",
			801 => x"feaa0cdd",
			802 => x"07069b04",
			803 => x"02610cdd",
			804 => x"feff0cdd",
			805 => x"fe6b0cdd",
			806 => x"01006704",
			807 => x"fe680cdd",
			808 => x"0601911c",
			809 => x"0208e204",
			810 => x"04e30cdd",
			811 => x"06016308",
			812 => x"0f07eb04",
			813 => x"016e0cdd",
			814 => x"fca70cdd",
			815 => x"0d061108",
			816 => x"0305e104",
			817 => x"00000cdd",
			818 => x"fe5d0cdd",
			819 => x"08033904",
			820 => x"ffb80cdd",
			821 => x"01b80cdd",
			822 => x"fe5d0cdd",
			823 => x"02086010",
			824 => x"0e050004",
			825 => x"00000d79",
			826 => x"040baa04",
			827 => x"00000d79",
			828 => x"0b052204",
			829 => x"00000d79",
			830 => x"00e60d79",
			831 => x"00040718",
			832 => x"0a028e04",
			833 => x"00000d79",
			834 => x"0100ff10",
			835 => x"09010604",
			836 => x"00000d79",
			837 => x"08033608",
			838 => x"040abb04",
			839 => x"00000d79",
			840 => x"009e0d79",
			841 => x"00000d79",
			842 => x"00000d79",
			843 => x"040d880c",
			844 => x"09018008",
			845 => x"02086704",
			846 => x"00000d79",
			847 => x"ff170d79",
			848 => x"00000d79",
			849 => x"06018110",
			850 => x"0e04a504",
			851 => x"00000d79",
			852 => x"0b05e908",
			853 => x"06017f04",
			854 => x"005b0d79",
			855 => x"00000d79",
			856 => x"00000d79",
			857 => x"0e08f008",
			858 => x"0307b004",
			859 => x"00000d79",
			860 => x"ff680d79",
			861 => x"00000d79",
			862 => x"040d1b1c",
			863 => x"040c4404",
			864 => x"fe700ded",
			865 => x"0b053504",
			866 => x"fe6c0ded",
			867 => x"0a02ae10",
			868 => x"0100fa0c",
			869 => x"0a028e08",
			870 => x"040caf04",
			871 => x"008e0ded",
			872 => x"ffa70ded",
			873 => x"02a90ded",
			874 => x"feeb0ded",
			875 => x"fead0ded",
			876 => x"01006704",
			877 => x"fe6a0ded",
			878 => x"06019118",
			879 => x"07060014",
			880 => x"0900ab04",
			881 => x"088f0ded",
			882 => x"0505f608",
			883 => x"0305cc04",
			884 => x"00000ded",
			885 => x"fe840ded",
			886 => x"08033904",
			887 => x"ff9b0ded",
			888 => x"01870ded",
			889 => x"fdd80ded",
			890 => x"fe600ded",
			891 => x"06019730",
			892 => x"0d05f704",
			893 => x"ff7a0e51",
			894 => x"0208dd14",
			895 => x"05063310",
			896 => x"0a028304",
			897 => x"00000e51",
			898 => x"0e050004",
			899 => x"00000e51",
			900 => x"00040304",
			901 => x"00000e51",
			902 => x"00e00e51",
			903 => x"00000e51",
			904 => x"040d4208",
			905 => x"0d07b004",
			906 => x"ff750e51",
			907 => x"00000e51",
			908 => x"01009304",
			909 => x"00000e51",
			910 => x"0b063908",
			911 => x"0b05b804",
			912 => x"00000e51",
			913 => x"00750e51",
			914 => x"00000e51",
			915 => x"ff520e51",
			916 => x"040d1b24",
			917 => x"040c4404",
			918 => x"fe670efd",
			919 => x"0004070c",
			920 => x"0100fa08",
			921 => x"0a028304",
			922 => x"feef0efd",
			923 => x"0b4b0efd",
			924 => x"fe990efd",
			925 => x"0b053504",
			926 => x"fe610efd",
			927 => x"06015b04",
			928 => x"04a60efd",
			929 => x"0a02a108",
			930 => x"0100e804",
			931 => x"07af0efd",
			932 => x"fed30efd",
			933 => x"fe760efd",
			934 => x"0900bc08",
			935 => x"01007104",
			936 => x"fe610efd",
			937 => x"ffac0efd",
			938 => x"06018820",
			939 => x"0e073b10",
			940 => x"0901580c",
			941 => x"00049604",
			942 => x"069d0efd",
			943 => x"0f08aa04",
			944 => x"02020efd",
			945 => x"04220efd",
			946 => x"fe970efd",
			947 => x"0506e208",
			948 => x"0c056104",
			949 => x"02da0efd",
			950 => x"00000efd",
			951 => x"0705b904",
			952 => x"20860efd",
			953 => x"0a130efd",
			954 => x"0a02d404",
			955 => x"00b80efd",
			956 => x"0d063704",
			957 => x"fbfb0efd",
			958 => x"fe5f0efd",
			959 => x"0900b704",
			960 => x"ff230f71",
			961 => x"0c050c18",
			962 => x"0b053504",
			963 => x"00000f71",
			964 => x"00040204",
			965 => x"00000f71",
			966 => x"0601910c",
			967 => x"0c04ce04",
			968 => x"00000f71",
			969 => x"07050104",
			970 => x"00000f71",
			971 => x"01080f71",
			972 => x"00000f71",
			973 => x"020b5b1c",
			974 => x"0b05f90c",
			975 => x"04100808",
			976 => x"0e058704",
			977 => x"00000f71",
			978 => x"ff760f71",
			979 => x"00000f71",
			980 => x"0100ed0c",
			981 => x"0100bd04",
			982 => x"00000f71",
			983 => x"040c4404",
			984 => x"00000f71",
			985 => x"00d20f71",
			986 => x"00000f71",
			987 => x"ff3d0f71",
			988 => x"0d05f704",
			989 => x"fe6d0fd5",
			990 => x"08031d04",
			991 => x"fe7f0fd5",
			992 => x"02089108",
			993 => x"0b056504",
			994 => x"02b30fd5",
			995 => x"ff470fd5",
			996 => x"06019918",
			997 => x"0b056508",
			998 => x"0305f904",
			999 => x"00d20fd5",
			1000 => x"fe950fd5",
			1001 => x"06016a08",
			1002 => x"04112a04",
			1003 => x"008b0fd5",
			1004 => x"feb50fd5",
			1005 => x"0100e204",
			1006 => x"012f0fd5",
			1007 => x"ffef0fd5",
			1008 => x"0a029b08",
			1009 => x"01011504",
			1010 => x"00c40fd5",
			1011 => x"ffb50fd5",
			1012 => x"fe810fd5",
			1013 => x"0d05f704",
			1014 => x"fe9c1059",
			1015 => x"0f07c710",
			1016 => x"0f06e304",
			1017 => x"00001059",
			1018 => x"040baa04",
			1019 => x"00001059",
			1020 => x"0c054604",
			1021 => x"01721059",
			1022 => x"00001059",
			1023 => x"09014314",
			1024 => x"04100808",
			1025 => x"0c054504",
			1026 => x"fe9a1059",
			1027 => x"00001059",
			1028 => x"0c054804",
			1029 => x"00951059",
			1030 => x"0410bb04",
			1031 => x"00001059",
			1032 => x"fecd1059",
			1033 => x"040c7f04",
			1034 => x"ff1c1059",
			1035 => x"0a02c310",
			1036 => x"0e071508",
			1037 => x"09015804",
			1038 => x"00001059",
			1039 => x"ffd91059",
			1040 => x"0705b804",
			1041 => x"01591059",
			1042 => x"00191059",
			1043 => x"0d075504",
			1044 => x"00001059",
			1045 => x"fff31059",
			1046 => x"0a028d04",
			1047 => x"ff1610cd",
			1048 => x"08033110",
			1049 => x"0100ff0c",
			1050 => x"0c050b04",
			1051 => x"000010cd",
			1052 => x"040d2e04",
			1053 => x"015c10cd",
			1054 => x"000010cd",
			1055 => x"000010cd",
			1056 => x"040c6604",
			1057 => x"ff1910cd",
			1058 => x"02089108",
			1059 => x"0305b004",
			1060 => x"000010cd",
			1061 => x"012f10cd",
			1062 => x"0100930c",
			1063 => x"08040d08",
			1064 => x"0f073b04",
			1065 => x"000010cd",
			1066 => x"ff4f10cd",
			1067 => x"000010cd",
			1068 => x"06017008",
			1069 => x"0b05b704",
			1070 => x"000010cd",
			1071 => x"009610cd",
			1072 => x"04100804",
			1073 => x"ffc410cd",
			1074 => x"000010cd",
			1075 => x"040d1b2c",
			1076 => x"0b053504",
			1077 => x"fe671171",
			1078 => x"0d064714",
			1079 => x"05061508",
			1080 => x"01007304",
			1081 => x"02c41171",
			1082 => x"fe8c1171",
			1083 => x"0208dd08",
			1084 => x"00040204",
			1085 => x"ffd11171",
			1086 => x"08b11171",
			1087 => x"ff601171",
			1088 => x"040c4404",
			1089 => x"fe6a1171",
			1090 => x"0003fb0c",
			1091 => x"0a028e04",
			1092 => x"fffa1171",
			1093 => x"01011f04",
			1094 => x"01e11171",
			1095 => x"00001171",
			1096 => x"fea31171",
			1097 => x"01006704",
			1098 => x"fe6d1171",
			1099 => x"0705ce1c",
			1100 => x"0f073904",
			1101 => x"03571171",
			1102 => x"0b056308",
			1103 => x"00059f04",
			1104 => x"fe6f1171",
			1105 => x"01381171",
			1106 => x"0c052808",
			1107 => x"00049604",
			1108 => x"04a11171",
			1109 => x"01961171",
			1110 => x"06016604",
			1111 => x"fdd31171",
			1112 => x"012b1171",
			1113 => x"0c059904",
			1114 => x"00001171",
			1115 => x"fe561171",
			1116 => x"0900c804",
			1117 => x"fe8911f5",
			1118 => x"0a02c320",
			1119 => x"0003e104",
			1120 => x"fed111f5",
			1121 => x"0c04ee04",
			1122 => x"ff1d11f5",
			1123 => x"0c050c0c",
			1124 => x"0a029304",
			1125 => x"01eb11f5",
			1126 => x"00045f04",
			1127 => x"ffc411f5",
			1128 => x"011911f5",
			1129 => x"0d06f904",
			1130 => x"ff3811f5",
			1131 => x"0901a104",
			1132 => x"00df11f5",
			1133 => x"ffe811f5",
			1134 => x"00055418",
			1135 => x"0c056210",
			1136 => x"0c05280c",
			1137 => x"07053204",
			1138 => x"ffa311f5",
			1139 => x"0f091f04",
			1140 => x"003211f5",
			1141 => x"000011f5",
			1142 => x"fe7711f5",
			1143 => x"0c059e04",
			1144 => x"007f11f5",
			1145 => x"ffbe11f5",
			1146 => x"030bd404",
			1147 => x"00e711f5",
			1148 => x"000011f5",
			1149 => x"0a028d04",
			1150 => x"ff041271",
			1151 => x"08033110",
			1152 => x"0100ff0c",
			1153 => x"0c050b04",
			1154 => x"00001271",
			1155 => x"040d2e04",
			1156 => x"017a1271",
			1157 => x"00001271",
			1158 => x"00001271",
			1159 => x"040c6604",
			1160 => x"ff0a1271",
			1161 => x"02089108",
			1162 => x"0305b004",
			1163 => x"00001271",
			1164 => x"014d1271",
			1165 => x"06017010",
			1166 => x"0e05f708",
			1167 => x"0c052e04",
			1168 => x"00001271",
			1169 => x"ffc31271",
			1170 => x"0b05b704",
			1171 => x"00001271",
			1172 => x"00a31271",
			1173 => x"04100808",
			1174 => x"040cd804",
			1175 => x"00001271",
			1176 => x"ff2b1271",
			1177 => x"0a035d04",
			1178 => x"001d1271",
			1179 => x"00001271",
			1180 => x"0b053504",
			1181 => x"fe7912e5",
			1182 => x"040baa04",
			1183 => x"fea012e5",
			1184 => x"08036814",
			1185 => x"0100fa10",
			1186 => x"02089f04",
			1187 => x"01e912e5",
			1188 => x"0506d204",
			1189 => x"ff1e12e5",
			1190 => x"0a028d04",
			1191 => x"000012e5",
			1192 => x"013312e5",
			1193 => x"ff6b12e5",
			1194 => x"0c054810",
			1195 => x"040e2304",
			1196 => x"fedf12e5",
			1197 => x"020a8608",
			1198 => x"0c052e04",
			1199 => x"015a12e5",
			1200 => x"000012e5",
			1201 => x"ff9012e5",
			1202 => x"06016b04",
			1203 => x"fe2a12e5",
			1204 => x"040eab04",
			1205 => x"ff3d12e5",
			1206 => x"0c059f04",
			1207 => x"00d912e5",
			1208 => x"ff8e12e5",
			1209 => x"0d05f704",
			1210 => x"fef71381",
			1211 => x"06014f10",
			1212 => x"0d063f0c",
			1213 => x"040baa04",
			1214 => x"00001381",
			1215 => x"0f06c104",
			1216 => x"00001381",
			1217 => x"01041381",
			1218 => x"00001381",
			1219 => x"0506b914",
			1220 => x"04100808",
			1221 => x"0f078704",
			1222 => x"00001381",
			1223 => x"fee41381",
			1224 => x"0c054808",
			1225 => x"0e04ad04",
			1226 => x"00001381",
			1227 => x"00341381",
			1228 => x"00001381",
			1229 => x"0705a210",
			1230 => x"0100c804",
			1231 => x"00001381",
			1232 => x"08033404",
			1233 => x"00001381",
			1234 => x"0308dd04",
			1235 => x"00ef1381",
			1236 => x"00001381",
			1237 => x"0100e70c",
			1238 => x"06017804",
			1239 => x"00001381",
			1240 => x"0a030404",
			1241 => x"00891381",
			1242 => x"00001381",
			1243 => x"0f0b1708",
			1244 => x"06017004",
			1245 => x"00001381",
			1246 => x"ff561381",
			1247 => x"00001381",
			1248 => x"07050408",
			1249 => x"0209ef04",
			1250 => x"feb11425",
			1251 => x"00001425",
			1252 => x"0705060c",
			1253 => x"0208e408",
			1254 => x"0d05f704",
			1255 => x"00001425",
			1256 => x"01901425",
			1257 => x"00001425",
			1258 => x"08036814",
			1259 => x"040baa04",
			1260 => x"ff111425",
			1261 => x"0100fa0c",
			1262 => x"01007e04",
			1263 => x"00001425",
			1264 => x"0d061104",
			1265 => x"00001425",
			1266 => x"00cb1425",
			1267 => x"00001425",
			1268 => x"0f084f14",
			1269 => x"0601660c",
			1270 => x"0410bb04",
			1271 => x"00001425",
			1272 => x"05061504",
			1273 => x"00001425",
			1274 => x"ff961425",
			1275 => x"02096604",
			1276 => x"00001425",
			1277 => x"00a91425",
			1278 => x"0100bb08",
			1279 => x"0306a504",
			1280 => x"00001425",
			1281 => x"fee11425",
			1282 => x"0100c908",
			1283 => x"020aaf04",
			1284 => x"006c1425",
			1285 => x"00001425",
			1286 => x"0100d404",
			1287 => x"ff3b1425",
			1288 => x"00001425",
			1289 => x"040d1b30",
			1290 => x"0b053504",
			1291 => x"fe6814e1",
			1292 => x"0d064718",
			1293 => x"0d063808",
			1294 => x"0900ba04",
			1295 => x"020114e1",
			1296 => x"fe9414e1",
			1297 => x"0c04ee04",
			1298 => x"ff3014e1",
			1299 => x"0b056908",
			1300 => x"06017004",
			1301 => x"069914e1",
			1302 => x"000014e1",
			1303 => x"000014e1",
			1304 => x"040c4404",
			1305 => x"fe6b14e1",
			1306 => x"0003fb0c",
			1307 => x"0a028e04",
			1308 => x"000014e1",
			1309 => x"0901d004",
			1310 => x"01c114e1",
			1311 => x"000014e1",
			1312 => x"feac14e1",
			1313 => x"01006704",
			1314 => x"fe6f14e1",
			1315 => x"0705ce20",
			1316 => x"06015704",
			1317 => x"035214e1",
			1318 => x"0b05630c",
			1319 => x"03061908",
			1320 => x"0d05f704",
			1321 => x"ff5814e1",
			1322 => x"015714e1",
			1323 => x"fe8214e1",
			1324 => x"0c052808",
			1325 => x"00049604",
			1326 => x"03dd14e1",
			1327 => x"018e14e1",
			1328 => x"06016604",
			1329 => x"fe1f14e1",
			1330 => x"011714e1",
			1331 => x"0a02fd08",
			1332 => x"040eab04",
			1333 => x"fef114e1",
			1334 => x"009814e1",
			1335 => x"fe4614e1",
			1336 => x"0d05f704",
			1337 => x"fe8c159d",
			1338 => x"0208dd24",
			1339 => x"07051f10",
			1340 => x"00040204",
			1341 => x"0000159d",
			1342 => x"0a02ae08",
			1343 => x"07050404",
			1344 => x"0000159d",
			1345 => x"0240159d",
			1346 => x"0000159d",
			1347 => x"040c8c04",
			1348 => x"ff7c159d",
			1349 => x"05060804",
			1350 => x"0000159d",
			1351 => x"05063308",
			1352 => x"07057304",
			1353 => x"00ae159d",
			1354 => x"0000159d",
			1355 => x"0000159d",
			1356 => x"0f08dd20",
			1357 => x"06016f0c",
			1358 => x"020a1008",
			1359 => x"0f07ce04",
			1360 => x"0000159d",
			1361 => x"ff15159d",
			1362 => x"0000159d",
			1363 => x"040d8808",
			1364 => x"040d6e04",
			1365 => x"ff90159d",
			1366 => x"0000159d",
			1367 => x"0b061908",
			1368 => x"0b054504",
			1369 => x"0000159d",
			1370 => x"0151159d",
			1371 => x"0000159d",
			1372 => x"0d079608",
			1373 => x"0f08f004",
			1374 => x"0000159d",
			1375 => x"fe86159d",
			1376 => x"0100fa0c",
			1377 => x"020b7708",
			1378 => x"08031d04",
			1379 => x"0000159d",
			1380 => x"011a159d",
			1381 => x"ffb5159d",
			1382 => x"ff26159d",
			1383 => x"0d05f704",
			1384 => x"fe6c1639",
			1385 => x"0c059e3c",
			1386 => x"0e05d81c",
			1387 => x"0f06e304",
			1388 => x"fede1639",
			1389 => x"06014e08",
			1390 => x"0b055204",
			1391 => x"03781639",
			1392 => x"00001639",
			1393 => x"040e2308",
			1394 => x"03061904",
			1395 => x"00001639",
			1396 => x"ff7f1639",
			1397 => x"07051c04",
			1398 => x"00001639",
			1399 => x"019a1639",
			1400 => x"01009204",
			1401 => x"fe811639",
			1402 => x"0506b910",
			1403 => x"09010f08",
			1404 => x"0c050704",
			1405 => x"ff4c1639",
			1406 => x"01b51639",
			1407 => x"0d06c704",
			1408 => x"fe851639",
			1409 => x"00001639",
			1410 => x"09018708",
			1411 => x"06019404",
			1412 => x"016f1639",
			1413 => x"ff451639",
			1414 => x"ff111639",
			1415 => x"06019604",
			1416 => x"fe7d1639",
			1417 => x"0f0b1c08",
			1418 => x"01010b04",
			1419 => x"013a1639",
			1420 => x"ff0e1639",
			1421 => x"fea41639",
			1422 => x"040c2404",
			1423 => x"fe8416f5",
			1424 => x"08036838",
			1425 => x"08036120",
			1426 => x"08034418",
			1427 => x"040ce10c",
			1428 => x"0e0a2a08",
			1429 => x"0a028304",
			1430 => x"000016f5",
			1431 => x"013116f5",
			1432 => x"000016f5",
			1433 => x"08033f08",
			1434 => x"0705ba04",
			1435 => x"ff5b16f5",
			1436 => x"000016f5",
			1437 => x"000016f5",
			1438 => x"040df504",
			1439 => x"ff7716f5",
			1440 => x"000016f5",
			1441 => x"0f071708",
			1442 => x"0b04c104",
			1443 => x"000016f5",
			1444 => x"04f116f5",
			1445 => x"040c6604",
			1446 => x"000016f5",
			1447 => x"0100e008",
			1448 => x"0505cc04",
			1449 => x"000016f5",
			1450 => x"017c16f5",
			1451 => x"000016f5",
			1452 => x"0601881c",
			1453 => x"040e2304",
			1454 => x"feb516f5",
			1455 => x"0c052808",
			1456 => x"0b056304",
			1457 => x"000016f5",
			1458 => x"011516f5",
			1459 => x"06017308",
			1460 => x"040fc604",
			1461 => x"000016f5",
			1462 => x"fee816f5",
			1463 => x"0100df04",
			1464 => x"009016f5",
			1465 => x"000016f5",
			1466 => x"09017404",
			1467 => x"fe6f16f5",
			1468 => x"000016f5",
			1469 => x"0d05f704",
			1470 => x"fe7317cb",
			1471 => x"0c050c1c",
			1472 => x"0e05960c",
			1473 => x"040c2404",
			1474 => x"000017cb",
			1475 => x"06017c04",
			1476 => x"01bc17cb",
			1477 => x"000017cb",
			1478 => x"0c050a08",
			1479 => x"04100804",
			1480 => x"fea417cb",
			1481 => x"002817cb",
			1482 => x"03071b04",
			1483 => x"000017cb",
			1484 => x"01e617cb",
			1485 => x"06016b1c",
			1486 => x"0c052508",
			1487 => x"0004b804",
			1488 => x"000017cb",
			1489 => x"002b17cb",
			1490 => x"0b05870c",
			1491 => x"0b058504",
			1492 => x"ff9a17cb",
			1493 => x"0d065104",
			1494 => x"000017cb",
			1495 => x"fab417cb",
			1496 => x"07055d04",
			1497 => x"000017cb",
			1498 => x"fe4317cb",
			1499 => x"0601811c",
			1500 => x"040d880c",
			1501 => x"0d075504",
			1502 => x"fef717cb",
			1503 => x"0c059e04",
			1504 => x"00d917cb",
			1505 => x"ff7817cb",
			1506 => x"00048e08",
			1507 => x"0209c904",
			1508 => x"016117cb",
			1509 => x"ff5b17cb",
			1510 => x"0305c004",
			1511 => x"000017cb",
			1512 => x"017517cb",
			1513 => x"020b0808",
			1514 => x"03079c04",
			1515 => x"000017cb",
			1516 => x"fe7717cb",
			1517 => x"030a6908",
			1518 => x"0a02d404",
			1519 => x"011f17cb",
			1520 => x"000017cb",
			1521 => x"fee817cb",
			1522 => x"000017cd",
			1523 => x"000017d1",
			1524 => x"000017d5",
			1525 => x"000017d9",
			1526 => x"000017dd",
			1527 => x"000017e1",
			1528 => x"000017e5",
			1529 => x"000017e9",
			1530 => x"000017ed",
			1531 => x"000017f1",
			1532 => x"0208dd04",
			1533 => x"000017fd",
			1534 => x"000017fd",
			1535 => x"0100bd04",
			1536 => x"ffff1811",
			1537 => x"0100f304",
			1538 => x"00081811",
			1539 => x"00001811",
			1540 => x"0c054808",
			1541 => x"0c04b204",
			1542 => x"00001825",
			1543 => x"001c1825",
			1544 => x"00001825",
			1545 => x"06019708",
			1546 => x"06014604",
			1547 => x"00001839",
			1548 => x"00181839",
			1549 => x"00001839",
			1550 => x"0e078e08",
			1551 => x"04100804",
			1552 => x"ffce184d",
			1553 => x"0000184d",
			1554 => x"0000184d",
			1555 => x"0f08dd08",
			1556 => x"0f070104",
			1557 => x"00001869",
			1558 => x"00221869",
			1559 => x"0f0abc04",
			1560 => x"ffdd1869",
			1561 => x"00001869",
			1562 => x"0f08c608",
			1563 => x"0f070104",
			1564 => x"00001885",
			1565 => x"00021885",
			1566 => x"0f0aed04",
			1567 => x"ffdd1885",
			1568 => x"00001885",
			1569 => x"02086004",
			1570 => x"000018a1",
			1571 => x"040d8808",
			1572 => x"0e097704",
			1573 => x"ff6b18a1",
			1574 => x"000018a1",
			1575 => x"000018a1",
			1576 => x"0004e90c",
			1577 => x"00041404",
			1578 => x"000018bd",
			1579 => x"0f071d04",
			1580 => x"000018bd",
			1581 => x"ffca18bd",
			1582 => x"000018bd",
			1583 => x"08034104",
			1584 => x"000018d9",
			1585 => x"0c04e904",
			1586 => x"000018d9",
			1587 => x"00043e04",
			1588 => x"000018d9",
			1589 => x"ffdc18d9",
			1590 => x"0e055a04",
			1591 => x"000018f5",
			1592 => x"0a028d04",
			1593 => x"000018f5",
			1594 => x"0e0a2a04",
			1595 => x"002518f5",
			1596 => x"000018f5",
			1597 => x"0f08c608",
			1598 => x"0f070104",
			1599 => x"00001919",
			1600 => x"00031919",
			1601 => x"0f0aed08",
			1602 => x"0f08dd04",
			1603 => x"00001919",
			1604 => x"ffd11919",
			1605 => x"00001919",
			1606 => x"0c050c0c",
			1607 => x"07050104",
			1608 => x"00001945",
			1609 => x"0d05f704",
			1610 => x"00001945",
			1611 => x"00141945",
			1612 => x"0d075508",
			1613 => x"07054904",
			1614 => x"00001945",
			1615 => x"ffd01945",
			1616 => x"00001945",
			1617 => x"040dca0c",
			1618 => x"02085b04",
			1619 => x"00001971",
			1620 => x"020b0f04",
			1621 => x"ff841971",
			1622 => x"00001971",
			1623 => x"0d06c704",
			1624 => x"00001971",
			1625 => x"0d083204",
			1626 => x"00201971",
			1627 => x"00001971",
			1628 => x"07058c10",
			1629 => x"07050404",
			1630 => x"00001995",
			1631 => x"0c052e08",
			1632 => x"0c04b204",
			1633 => x"00001995",
			1634 => x"00271995",
			1635 => x"00001995",
			1636 => x"ffff1995",
			1637 => x"0c052810",
			1638 => x"01006704",
			1639 => x"000019b9",
			1640 => x"0100d008",
			1641 => x"0c04b204",
			1642 => x"000019b9",
			1643 => x"004a19b9",
			1644 => x"000019b9",
			1645 => x"ffff19b9",
			1646 => x"0e055204",
			1647 => x"000019dd",
			1648 => x"0a028d04",
			1649 => x"000019dd",
			1650 => x"0e0a2a08",
			1651 => x"0a030804",
			1652 => x"002419dd",
			1653 => x"000019dd",
			1654 => x"000019dd",
			1655 => x"0900b704",
			1656 => x"00001a01",
			1657 => x"0901630c",
			1658 => x"0b053504",
			1659 => x"00001a01",
			1660 => x"0b073304",
			1661 => x"00211a01",
			1662 => x"00001a01",
			1663 => x"00001a01",
			1664 => x"0c052810",
			1665 => x"07050404",
			1666 => x"00001a35",
			1667 => x"07058b08",
			1668 => x"0c04b204",
			1669 => x"00001a35",
			1670 => x"002d1a35",
			1671 => x"00001a35",
			1672 => x"0a029004",
			1673 => x"00001a35",
			1674 => x"0a030404",
			1675 => x"ffe31a35",
			1676 => x"00001a35",
			1677 => x"0004140c",
			1678 => x"0a028d04",
			1679 => x"00001a69",
			1680 => x"0a029b04",
			1681 => x"00171a69",
			1682 => x"00001a69",
			1683 => x"040e230c",
			1684 => x"0f071704",
			1685 => x"00001a69",
			1686 => x"0c058004",
			1687 => x"ff991a69",
			1688 => x"00001a69",
			1689 => x"00001a69",
			1690 => x"040dca0c",
			1691 => x"02085b04",
			1692 => x"00001a9d",
			1693 => x"0f0abc04",
			1694 => x"ff7a1a9d",
			1695 => x"00001a9d",
			1696 => x"06016604",
			1697 => x"00001a9d",
			1698 => x"06019108",
			1699 => x"0d06d204",
			1700 => x"00001a9d",
			1701 => x"003e1a9d",
			1702 => x"00001a9d",
			1703 => x"040e2310",
			1704 => x"0a029004",
			1705 => x"00001ad9",
			1706 => x"0f071704",
			1707 => x"00001ad9",
			1708 => x"0003fb04",
			1709 => x"00001ad9",
			1710 => x"ff961ad9",
			1711 => x"0100c90c",
			1712 => x"01007304",
			1713 => x"00001ad9",
			1714 => x"0f09a304",
			1715 => x"00311ad9",
			1716 => x"00001ad9",
			1717 => x"00001ad9",
			1718 => x"0e073b08",
			1719 => x"05070d04",
			1720 => x"fff31b0d",
			1721 => x"00001b0d",
			1722 => x"0100fa10",
			1723 => x"0100c204",
			1724 => x"00001b0d",
			1725 => x"0506d504",
			1726 => x"00001b0d",
			1727 => x"05086a04",
			1728 => x"00561b0d",
			1729 => x"00001b0d",
			1730 => x"00001b0d",
			1731 => x"06016608",
			1732 => x"040c2404",
			1733 => x"ffd71b49",
			1734 => x"00001b49",
			1735 => x"06017410",
			1736 => x"01009b04",
			1737 => x"00001b49",
			1738 => x"0100f308",
			1739 => x"040adc04",
			1740 => x"00001b49",
			1741 => x"005e1b49",
			1742 => x"00001b49",
			1743 => x"040fc604",
			1744 => x"ffec1b49",
			1745 => x"00001b49",
			1746 => x"09014110",
			1747 => x"0f07d504",
			1748 => x"00001b8d",
			1749 => x"04120c08",
			1750 => x"05070d04",
			1751 => x"ffb71b8d",
			1752 => x"00001b8d",
			1753 => x"00001b8d",
			1754 => x"0100f510",
			1755 => x"0901870c",
			1756 => x"0100f308",
			1757 => x"0100c204",
			1758 => x"00001b8d",
			1759 => x"00091b8d",
			1760 => x"00001b8d",
			1761 => x"00001b8d",
			1762 => x"00001b8d",
			1763 => x"03071b08",
			1764 => x"0306ff04",
			1765 => x"ffef1bc9",
			1766 => x"00001bc9",
			1767 => x"0100fa14",
			1768 => x"0100bb04",
			1769 => x"00001bc9",
			1770 => x"0e071504",
			1771 => x"00001bc9",
			1772 => x"03078c04",
			1773 => x"00001bc9",
			1774 => x"030a8104",
			1775 => x"00521bc9",
			1776 => x"00001bc9",
			1777 => x"00001bc9",
			1778 => x"040cce0c",
			1779 => x"06019608",
			1780 => x"0a02ac04",
			1781 => x"ff8b1c0d",
			1782 => x"00001c0d",
			1783 => x"00001c0d",
			1784 => x"06019114",
			1785 => x"0705fd10",
			1786 => x"06016604",
			1787 => x"00001c0d",
			1788 => x"0900e704",
			1789 => x"00001c0d",
			1790 => x"0a028d04",
			1791 => x"00001c0d",
			1792 => x"00511c0d",
			1793 => x"00001c0d",
			1794 => x"00001c0d",
			1795 => x"00040714",
			1796 => x"0003f704",
			1797 => x"00001c61",
			1798 => x"05061504",
			1799 => x"00001c61",
			1800 => x"0100fa08",
			1801 => x"08033404",
			1802 => x"006d1c61",
			1803 => x"00001c61",
			1804 => x"00001c61",
			1805 => x"0f074908",
			1806 => x"0e050004",
			1807 => x"00001c61",
			1808 => x"00061c61",
			1809 => x"040e230c",
			1810 => x"02088304",
			1811 => x"00001c61",
			1812 => x"0e097704",
			1813 => x"ff7f1c61",
			1814 => x"00001c61",
			1815 => x"00001c61",
			1816 => x"0e055a04",
			1817 => x"00001c95",
			1818 => x"0a028d04",
			1819 => x"00001c95",
			1820 => x"07064610",
			1821 => x"0900b704",
			1822 => x"00001c95",
			1823 => x"0100fa08",
			1824 => x"07050404",
			1825 => x"00001c95",
			1826 => x"003a1c95",
			1827 => x"00001c95",
			1828 => x"00001c95",
			1829 => x"0c052818",
			1830 => x"0d05f704",
			1831 => x"00001ce1",
			1832 => x"08032504",
			1833 => x"00001ce1",
			1834 => x"020a9b0c",
			1835 => x"00040204",
			1836 => x"00001ce1",
			1837 => x"07050104",
			1838 => x"00001ce1",
			1839 => x"00701ce1",
			1840 => x"00001ce1",
			1841 => x"0209c104",
			1842 => x"00001ce1",
			1843 => x"00040704",
			1844 => x"00001ce1",
			1845 => x"0005b804",
			1846 => x"ffb31ce1",
			1847 => x"00001ce1",
			1848 => x"00040714",
			1849 => x"0003f704",
			1850 => x"00001d3d",
			1851 => x"05061504",
			1852 => x"00001d3d",
			1853 => x"08033108",
			1854 => x"040cbf04",
			1855 => x"00721d3d",
			1856 => x"00001d3d",
			1857 => x"00001d3d",
			1858 => x"0f07490c",
			1859 => x"0e050004",
			1860 => x"00001d3d",
			1861 => x"0305b004",
			1862 => x"00001d3d",
			1863 => x"00121d3d",
			1864 => x"0005b80c",
			1865 => x"0e08f008",
			1866 => x"02088304",
			1867 => x"00001d3d",
			1868 => x"ffa71d3d",
			1869 => x"00001d3d",
			1870 => x"00001d3d",
			1871 => x"09010608",
			1872 => x"040fc604",
			1873 => x"ffa41d89",
			1874 => x"00001d89",
			1875 => x"0100d018",
			1876 => x"06016b04",
			1877 => x"00001d89",
			1878 => x"03087510",
			1879 => x"00040304",
			1880 => x"00001d89",
			1881 => x"0b056504",
			1882 => x"00001d89",
			1883 => x"06019104",
			1884 => x"00c71d89",
			1885 => x"00001d89",
			1886 => x"00001d89",
			1887 => x"0f08c604",
			1888 => x"00001d89",
			1889 => x"fffa1d89",
			1890 => x"040cce0c",
			1891 => x"06019608",
			1892 => x"0a02ac04",
			1893 => x"ff801dd5",
			1894 => x"00001dd5",
			1895 => x"00001dd5",
			1896 => x"06019118",
			1897 => x"0705fd14",
			1898 => x"06016604",
			1899 => x"00001dd5",
			1900 => x"01008604",
			1901 => x"00001dd5",
			1902 => x"0a028d04",
			1903 => x"00001dd5",
			1904 => x"07051c04",
			1905 => x"00001dd5",
			1906 => x"005c1dd5",
			1907 => x"00001dd5",
			1908 => x"00001dd5",
			1909 => x"0f08dd1c",
			1910 => x"0c04b204",
			1911 => x"00001e19",
			1912 => x"0a027f04",
			1913 => x"00001e19",
			1914 => x"0f06e304",
			1915 => x"00001e19",
			1916 => x"020a060c",
			1917 => x"0a02fd08",
			1918 => x"0c056504",
			1919 => x"00631e19",
			1920 => x"00001e19",
			1921 => x"00001e19",
			1922 => x"00001e19",
			1923 => x"0c050b04",
			1924 => x"00001e19",
			1925 => x"ffcf1e19",
			1926 => x"040c7f18",
			1927 => x"02086010",
			1928 => x"0b053504",
			1929 => x"00001e8d",
			1930 => x"0b054508",
			1931 => x"06014104",
			1932 => x"00001e8d",
			1933 => x"003c1e8d",
			1934 => x"00001e8d",
			1935 => x"07069b04",
			1936 => x"ff241e8d",
			1937 => x"00001e8d",
			1938 => x"0a02d410",
			1939 => x"0100fa0c",
			1940 => x"0a028d04",
			1941 => x"00001e8d",
			1942 => x"0d05f704",
			1943 => x"00001e8d",
			1944 => x"00ab1e8d",
			1945 => x"00001e8d",
			1946 => x"0f080504",
			1947 => x"00001e8d",
			1948 => x"020a0604",
			1949 => x"00001e8d",
			1950 => x"03068304",
			1951 => x"00001e8d",
			1952 => x"0d073004",
			1953 => x"ff5e1e8d",
			1954 => x"00001e8d",
			1955 => x"06016b10",
			1956 => x"0901760c",
			1957 => x"0f074904",
			1958 => x"00001ee1",
			1959 => x"0a030804",
			1960 => x"ff931ee1",
			1961 => x"00001ee1",
			1962 => x"00001ee1",
			1963 => x"09016318",
			1964 => x"09010604",
			1965 => x"00001ee1",
			1966 => x"03087510",
			1967 => x"0c050a04",
			1968 => x"00001ee1",
			1969 => x"040adc04",
			1970 => x"00001ee1",
			1971 => x"0a031004",
			1972 => x"00bf1ee1",
			1973 => x"00001ee1",
			1974 => x"00001ee1",
			1975 => x"00001ee1",
			1976 => x"0f09b124",
			1977 => x"03071b0c",
			1978 => x"04100808",
			1979 => x"0f074904",
			1980 => x"00001f35",
			1981 => x"ffc71f35",
			1982 => x"00001f35",
			1983 => x"01009b04",
			1984 => x"00001f35",
			1985 => x"0c059e10",
			1986 => x"06016704",
			1987 => x"00001f35",
			1988 => x"0c050a04",
			1989 => x"00001f35",
			1990 => x"040adc04",
			1991 => x"00001f35",
			1992 => x"00591f35",
			1993 => x"00001f35",
			1994 => x"0003fb04",
			1995 => x"00001f35",
			1996 => x"ff791f35",
			1997 => x"0d05f704",
			1998 => x"ffd61f71",
			1999 => x"07058c18",
			2000 => x"00040204",
			2001 => x"00001f71",
			2002 => x"03087510",
			2003 => x"08036f0c",
			2004 => x"0c056308",
			2005 => x"07050404",
			2006 => x"00001f71",
			2007 => x"00a81f71",
			2008 => x"00001f71",
			2009 => x"00001f71",
			2010 => x"00001f71",
			2011 => x"00001f71",
			2012 => x"01008e04",
			2013 => x"00001fad",
			2014 => x"0100fa18",
			2015 => x"0a027f04",
			2016 => x"00001fad",
			2017 => x"07050504",
			2018 => x"00001fad",
			2019 => x"0d063804",
			2020 => x"00001fad",
			2021 => x"0601a608",
			2022 => x"0c04ed04",
			2023 => x"00001fad",
			2024 => x"00501fad",
			2025 => x"00001fad",
			2026 => x"00001fad",
			2027 => x"0e055a04",
			2028 => x"00001fe9",
			2029 => x"07058c18",
			2030 => x"08032504",
			2031 => x"00001fe9",
			2032 => x"0900b704",
			2033 => x"00001fe9",
			2034 => x"07050404",
			2035 => x"00001fe9",
			2036 => x"06018e08",
			2037 => x"040adc04",
			2038 => x"00001fe9",
			2039 => x"005e1fe9",
			2040 => x"00001fe9",
			2041 => x"00001fe9",
			2042 => x"01008e14",
			2043 => x"0f07490c",
			2044 => x"0e050004",
			2045 => x"0000205d",
			2046 => x"040c2404",
			2047 => x"0000205d",
			2048 => x"0065205d",
			2049 => x"08040d04",
			2050 => x"ff70205d",
			2051 => x"0000205d",
			2052 => x"0100c918",
			2053 => x"00040204",
			2054 => x"0000205d",
			2055 => x"07050504",
			2056 => x"0000205d",
			2057 => x"0308750c",
			2058 => x"05061504",
			2059 => x"0000205d",
			2060 => x"0c04ee04",
			2061 => x"0000205d",
			2062 => x"00d0205d",
			2063 => x"0000205d",
			2064 => x"0209c904",
			2065 => x"0000205d",
			2066 => x"07057504",
			2067 => x"0000205d",
			2068 => x"07069b04",
			2069 => x"ffc1205d",
			2070 => x"0000205d",
			2071 => x"0209ce1c",
			2072 => x"0900b704",
			2073 => x"000020b9",
			2074 => x"00040204",
			2075 => x"000020b9",
			2076 => x"0b053504",
			2077 => x"000020b9",
			2078 => x"0601710c",
			2079 => x"08032504",
			2080 => x"000020b9",
			2081 => x"07050404",
			2082 => x"000020b9",
			2083 => x"006a20b9",
			2084 => x"000020b9",
			2085 => x"0c052804",
			2086 => x"000020b9",
			2087 => x"0e09770c",
			2088 => x"00040304",
			2089 => x"000020b9",
			2090 => x"0005b804",
			2091 => x"ff6b20b9",
			2092 => x"000020b9",
			2093 => x"000020b9",
			2094 => x"07058c24",
			2095 => x"0d05f704",
			2096 => x"ffa72115",
			2097 => x"06018e1c",
			2098 => x"040c8c10",
			2099 => x"0803370c",
			2100 => x"07051a08",
			2101 => x"08032804",
			2102 => x"00002115",
			2103 => x"00602115",
			2104 => x"00002115",
			2105 => x"ffff2115",
			2106 => x"01006704",
			2107 => x"00002115",
			2108 => x"08033a04",
			2109 => x"00002115",
			2110 => x"00a42115",
			2111 => x"00002115",
			2112 => x"0d075508",
			2113 => x"0209b104",
			2114 => x"00002115",
			2115 => x"ff792115",
			2116 => x"00002115",
			2117 => x"0d05f704",
			2118 => x"fecd2179",
			2119 => x"07058c24",
			2120 => x"08036e10",
			2121 => x"00040204",
			2122 => x"00002179",
			2123 => x"07050404",
			2124 => x"00002179",
			2125 => x"06019004",
			2126 => x"01702179",
			2127 => x"00002179",
			2128 => x"04100808",
			2129 => x"0b058504",
			2130 => x"ff5b2179",
			2131 => x"00002179",
			2132 => x"06016604",
			2133 => x"00002179",
			2134 => x"00076604",
			2135 => x"00ad2179",
			2136 => x"00002179",
			2137 => x"0209e808",
			2138 => x"0a028e04",
			2139 => x"fffc2179",
			2140 => x"00002179",
			2141 => x"ff252179",
			2142 => x"07050408",
			2143 => x"0209e804",
			2144 => x"fe6b21dd",
			2145 => x"000021dd",
			2146 => x"0c059e1c",
			2147 => x"0a036318",
			2148 => x"0003f704",
			2149 => x"feba21dd",
			2150 => x"02086004",
			2151 => x"035521dd",
			2152 => x"0b055608",
			2153 => x"040e6304",
			2154 => x"fea121dd",
			2155 => x"001621dd",
			2156 => x"06019004",
			2157 => x"00f721dd",
			2158 => x"febc21dd",
			2159 => x"fea021dd",
			2160 => x"020b1c04",
			2161 => x"fe6c21dd",
			2162 => x"030a6908",
			2163 => x"030a2804",
			2164 => x"ffd421dd",
			2165 => x"016c21dd",
			2166 => x"fe8e21dd",
			2167 => x"00040718",
			2168 => x"08031d04",
			2169 => x"ffde2261",
			2170 => x"0c04ee04",
			2171 => x"00002261",
			2172 => x"0100fa0c",
			2173 => x"08033608",
			2174 => x"040adc04",
			2175 => x"00002261",
			2176 => x"012f2261",
			2177 => x"00002261",
			2178 => x"00002261",
			2179 => x"06014e10",
			2180 => x"0305f904",
			2181 => x"ff9f2261",
			2182 => x"01006f04",
			2183 => x"00002261",
			2184 => x"040b9704",
			2185 => x"00002261",
			2186 => x"00d92261",
			2187 => x"040d4204",
			2188 => x"ff1f2261",
			2189 => x"06018110",
			2190 => x"0e07580c",
			2191 => x"0100ca08",
			2192 => x"0900e704",
			2193 => x"00002261",
			2194 => x"00242261",
			2195 => x"ffc22261",
			2196 => x"006a2261",
			2197 => x"04117604",
			2198 => x"ff512261",
			2199 => x"00002261",
			2200 => x"0f08dd34",
			2201 => x"07050408",
			2202 => x"0a034f04",
			2203 => x"ff7722dd",
			2204 => x"000022dd",
			2205 => x"07051f14",
			2206 => x"0208dd10",
			2207 => x"0e050004",
			2208 => x"000022dd",
			2209 => x"00040204",
			2210 => x"000022dd",
			2211 => x"08036804",
			2212 => x"010c22dd",
			2213 => x"000022dd",
			2214 => x"000022dd",
			2215 => x"0803960c",
			2216 => x"0f08a308",
			2217 => x"0305e104",
			2218 => x"000022dd",
			2219 => x"ff7f22dd",
			2220 => x"000022dd",
			2221 => x"06015f04",
			2222 => x"000022dd",
			2223 => x"0006ce04",
			2224 => x"005a22dd",
			2225 => x"000022dd",
			2226 => x"0b064b04",
			2227 => x"ff2922dd",
			2228 => x"0c059e04",
			2229 => x"000322dd",
			2230 => x"000022dd",
			2231 => x"040c2404",
			2232 => x"ff342341",
			2233 => x"08036618",
			2234 => x"0100fa14",
			2235 => x"01006704",
			2236 => x"00002341",
			2237 => x"0a02b30c",
			2238 => x"0a028e04",
			2239 => x"00002341",
			2240 => x"0d05f704",
			2241 => x"00002341",
			2242 => x"007d2341",
			2243 => x"00002341",
			2244 => x"00002341",
			2245 => x"06018814",
			2246 => x"040eab08",
			2247 => x"0100da04",
			2248 => x"fff72341",
			2249 => x"00002341",
			2250 => x"06016a04",
			2251 => x"00002341",
			2252 => x"01007304",
			2253 => x"00002341",
			2254 => x"00762341",
			2255 => x"ff8a2341",
			2256 => x"040d1b24",
			2257 => x"040c7f0c",
			2258 => x"020b1c04",
			2259 => x"fe7123c5",
			2260 => x"020b1f04",
			2261 => x"00da23c5",
			2262 => x"fe7523c5",
			2263 => x"08034114",
			2264 => x"0a028e0c",
			2265 => x"040caf08",
			2266 => x"06015f04",
			2267 => x"000023c5",
			2268 => x"013423c5",
			2269 => x"fef123c5",
			2270 => x"0c066f04",
			2271 => x"030e23c5",
			2272 => x"ff9d23c5",
			2273 => x"fe6b23c5",
			2274 => x"03055f04",
			2275 => x"fe6823c5",
			2276 => x"06019118",
			2277 => x"0c05a014",
			2278 => x"0505f604",
			2279 => x"fea523c5",
			2280 => x"0209c108",
			2281 => x"0a028e04",
			2282 => x"ff0323c5",
			2283 => x"02d523c5",
			2284 => x"040dca04",
			2285 => x"fe7f23c5",
			2286 => x"01a323c5",
			2287 => x"fd9923c5",
			2288 => x"fe5c23c5",
			2289 => x"040e2338",
			2290 => x"040cce1c",
			2291 => x"040c2404",
			2292 => x"bf9b2471",
			2293 => x"0803370c",
			2294 => x"030a7808",
			2295 => x"0a028304",
			2296 => x"bfcb2471",
			2297 => x"e14a2471",
			2298 => x"bfae2471",
			2299 => x"0b053504",
			2300 => x"bf992471",
			2301 => x"0d060304",
			2302 => x"c33a2471",
			2303 => x"bfa72471",
			2304 => x"0506e20c",
			2305 => x"05060604",
			2306 => x"bf9b2471",
			2307 => x"03073b04",
			2308 => x"cc652471",
			2309 => x"bfa52471",
			2310 => x"0a029304",
			2311 => x"df212471",
			2312 => x"08034208",
			2313 => x"0100eb04",
			2314 => x"d2f52471",
			2315 => x"c0722471",
			2316 => x"bfbc2471",
			2317 => x"01007104",
			2318 => x"bf982471",
			2319 => x"0f08b80c",
			2320 => x"040f7008",
			2321 => x"0d06e204",
			2322 => x"c03a2471",
			2323 => x"fb1b2471",
			2324 => x"10012471",
			2325 => x"0c059b0c",
			2326 => x"040eab08",
			2327 => x"0b060904",
			2328 => x"c0322471",
			2329 => x"cc652471",
			2330 => x"f3062471",
			2331 => x"bf992471",
			2332 => x"0d05f704",
			2333 => x"ff9b24e5",
			2334 => x"0208910c",
			2335 => x"00040204",
			2336 => x"000024e5",
			2337 => x"0c050c04",
			2338 => x"00d524e5",
			2339 => x"000024e5",
			2340 => x"0100bb0c",
			2341 => x"0e058704",
			2342 => x"000024e5",
			2343 => x"0005b804",
			2344 => x"ff6224e5",
			2345 => x"000024e5",
			2346 => x"0100c90c",
			2347 => x"0a02bb04",
			2348 => x"000024e5",
			2349 => x"0f09e104",
			2350 => x"009024e5",
			2351 => x"000024e5",
			2352 => x"0209c90c",
			2353 => x"0506d204",
			2354 => x"000024e5",
			2355 => x"0e07dc04",
			2356 => x"004f24e5",
			2357 => x"000024e5",
			2358 => x"020b0804",
			2359 => x"ff9424e5",
			2360 => x"000024e5",
			2361 => x"040c4404",
			2362 => x"fea52571",
			2363 => x"08036628",
			2364 => x"00046818",
			2365 => x"0209c10c",
			2366 => x"0a028e04",
			2367 => x"00002571",
			2368 => x"0c050704",
			2369 => x"00002571",
			2370 => x"006f2571",
			2371 => x"0e09c104",
			2372 => x"ffc62571",
			2373 => x"020b5b04",
			2374 => x"00012571",
			2375 => x"00002571",
			2376 => x"08035e04",
			2377 => x"00002571",
			2378 => x"00047908",
			2379 => x"0305b004",
			2380 => x"00002571",
			2381 => x"01f22571",
			2382 => x"00002571",
			2383 => x"0f08f014",
			2384 => x"0900e408",
			2385 => x"020a0604",
			2386 => x"ff002571",
			2387 => x"00002571",
			2388 => x"09015a08",
			2389 => x"0b05b804",
			2390 => x"00002571",
			2391 => x"01152571",
			2392 => x"00002571",
			2393 => x"0100c504",
			2394 => x"febe2571",
			2395 => x"00002571",
			2396 => x"040c4404",
			2397 => x"feb125f5",
			2398 => x"08036624",
			2399 => x"00046814",
			2400 => x"06016f08",
			2401 => x"06015e04",
			2402 => x"000025f5",
			2403 => x"ffda25f5",
			2404 => x"0c056204",
			2405 => x"000025f5",
			2406 => x"0c063404",
			2407 => x"005825f5",
			2408 => x"000025f5",
			2409 => x"08035e04",
			2410 => x"000025f5",
			2411 => x"00047908",
			2412 => x"0305b004",
			2413 => x"000025f5",
			2414 => x"01b925f5",
			2415 => x"000025f5",
			2416 => x"06018818",
			2417 => x"05063508",
			2418 => x"00056a04",
			2419 => x"ff1625f5",
			2420 => x"000025f5",
			2421 => x"06016b04",
			2422 => x"000025f5",
			2423 => x"09015a08",
			2424 => x"040e6304",
			2425 => x"000025f5",
			2426 => x"011525f5",
			2427 => x"000025f5",
			2428 => x"fecb25f5",
			2429 => x"040c7f0c",
			2430 => x"020b1c04",
			2431 => x"fe7a2689",
			2432 => x"0f0b1c04",
			2433 => x"01292689",
			2434 => x"fea02689",
			2435 => x"01007c18",
			2436 => x"08036108",
			2437 => x"08035b04",
			2438 => x"ff512689",
			2439 => x"06d62689",
			2440 => x"020a500c",
			2441 => x"01007604",
			2442 => x"fe712689",
			2443 => x"01007804",
			2444 => x"00382689",
			2445 => x"fec12689",
			2446 => x"00002689",
			2447 => x"020b5b24",
			2448 => x"03067808",
			2449 => x"05060604",
			2450 => x"00002689",
			2451 => x"01c02689",
			2452 => x"06016b0c",
			2453 => x"0c052a04",
			2454 => x"00002689",
			2455 => x"0209ab04",
			2456 => x"00002689",
			2457 => x"fdb62689",
			2458 => x"040df508",
			2459 => x"0b061904",
			2460 => x"fe9f2689",
			2461 => x"014a2689",
			2462 => x"0100df04",
			2463 => x"01842689",
			2464 => x"feeb2689",
			2465 => x"fe732689",
			2466 => x"040d1b1c",
			2467 => x"040c6604",
			2468 => x"fe732705",
			2469 => x"00046b14",
			2470 => x"02086204",
			2471 => x"057d2705",
			2472 => x"0a02a10c",
			2473 => x"0209dd04",
			2474 => x"feea2705",
			2475 => x"0508de04",
			2476 => x"02352705",
			2477 => x"00002705",
			2478 => x"fec92705",
			2479 => x"fe6d2705",
			2480 => x"01006704",
			2481 => x"fe692705",
			2482 => x"0601911c",
			2483 => x"0c04b304",
			2484 => x"0a862705",
			2485 => x"01007c08",
			2486 => x"0e053404",
			2487 => x"015a2705",
			2488 => x"fdde2705",
			2489 => x"0209c108",
			2490 => x"06017404",
			2491 => x"029f2705",
			2492 => x"00002705",
			2493 => x"0100de04",
			2494 => x"01782705",
			2495 => x"fe802705",
			2496 => x"fe5f2705",
			2497 => x"0900b704",
			2498 => x"ff382779",
			2499 => x"0c050c18",
			2500 => x"0d061104",
			2501 => x"00002779",
			2502 => x"0c04ed04",
			2503 => x"00002779",
			2504 => x"08032504",
			2505 => x"00002779",
			2506 => x"06019108",
			2507 => x"07050404",
			2508 => x"00002779",
			2509 => x"00fe2779",
			2510 => x"00002779",
			2511 => x"020b5b1c",
			2512 => x"0b05f90c",
			2513 => x"04100808",
			2514 => x"0e058704",
			2515 => x"00002779",
			2516 => x"ff862779",
			2517 => x"00002779",
			2518 => x"0a028d04",
			2519 => x"00002779",
			2520 => x"0100bf04",
			2521 => x"00002779",
			2522 => x"0100fa04",
			2523 => x"00ab2779",
			2524 => x"00002779",
			2525 => x"ff4e2779",
			2526 => x"01007c18",
			2527 => x"0d05f704",
			2528 => x"fe6827fd",
			2529 => x"0505ce04",
			2530 => x"08b527fd",
			2531 => x"0705450c",
			2532 => x"0d060304",
			2533 => x"ff2827fd",
			2534 => x"0d061104",
			2535 => x"005927fd",
			2536 => x"ffff27fd",
			2537 => x"fe5b27fd",
			2538 => x"0a028e04",
			2539 => x"fe6b27fd",
			2540 => x"0601a324",
			2541 => x"05060608",
			2542 => x"0e053404",
			2543 => x"000027fd",
			2544 => x"fe9827fd",
			2545 => x"0208dd0c",
			2546 => x"0e065a08",
			2547 => x"00043e04",
			2548 => x"ffb227fd",
			2549 => x"022227fd",
			2550 => x"064827fd",
			2551 => x"06016b08",
			2552 => x"0100b404",
			2553 => x"010927fd",
			2554 => x"fd8127fd",
			2555 => x"02099d04",
			2556 => x"ff0027fd",
			2557 => x"014c27fd",
			2558 => x"fe6d27fd",
			2559 => x"07050408",
			2560 => x"0a034f04",
			2561 => x"fee12891",
			2562 => x"00002891",
			2563 => x"02086710",
			2564 => x"02083004",
			2565 => x"00002891",
			2566 => x"040baa04",
			2567 => x"00002891",
			2568 => x"07055f04",
			2569 => x"01252891",
			2570 => x"00002891",
			2571 => x"040d420c",
			2572 => x"020b0f04",
			2573 => x"fef62891",
			2574 => x"030a6904",
			2575 => x"00732891",
			2576 => x"00002891",
			2577 => x"0004bc10",
			2578 => x"0308750c",
			2579 => x"0705b808",
			2580 => x"0c057204",
			2581 => x"01032891",
			2582 => x"00002891",
			2583 => x"00002891",
			2584 => x"00002891",
			2585 => x"04100808",
			2586 => x"09014504",
			2587 => x"ff0e2891",
			2588 => x"00002891",
			2589 => x"0e05e908",
			2590 => x"0c054304",
			2591 => x"00002891",
			2592 => x"ff912891",
			2593 => x"03092204",
			2594 => x"00672891",
			2595 => x"00002891",
			2596 => x"040c4404",
			2597 => x"feab291d",
			2598 => x"08036628",
			2599 => x"00046818",
			2600 => x"06016f08",
			2601 => x"0b058304",
			2602 => x"0000291d",
			2603 => x"ffaf291d",
			2604 => x"0b060904",
			2605 => x"0000291d",
			2606 => x"0a02ab08",
			2607 => x"0e0a2a04",
			2608 => x"007b291d",
			2609 => x"0000291d",
			2610 => x"0000291d",
			2611 => x"08035e04",
			2612 => x"0000291d",
			2613 => x"00047908",
			2614 => x"0305b004",
			2615 => x"0000291d",
			2616 => x"01cd291d",
			2617 => x"0000291d",
			2618 => x"06018818",
			2619 => x"05063508",
			2620 => x"00056a04",
			2621 => x"ff08291d",
			2622 => x"0000291d",
			2623 => x"06016b04",
			2624 => x"0000291d",
			2625 => x"0a02be04",
			2626 => x"0000291d",
			2627 => x"040e2304",
			2628 => x"0000291d",
			2629 => x"011d291d",
			2630 => x"fec1291d",
			2631 => x"040c7f1c",
			2632 => x"06016b04",
			2633 => x"fe6929d9",
			2634 => x"06016c0c",
			2635 => x"09010604",
			2636 => x"ff7a29d9",
			2637 => x"0d077004",
			2638 => x"057129d9",
			2639 => x"000029d9",
			2640 => x"09015f08",
			2641 => x"0100d004",
			2642 => x"feae29d9",
			2643 => x"012d29d9",
			2644 => x"fe7429d9",
			2645 => x"01007c1c",
			2646 => x"00047908",
			2647 => x"00047804",
			2648 => x"ff4029d9",
			2649 => x"050029d9",
			2650 => x"0900b104",
			2651 => x"fe6429d9",
			2652 => x"0100780c",
			2653 => x"01007308",
			2654 => x"0900b304",
			2655 => x"000029d9",
			2656 => x"ff6a29d9",
			2657 => x"006729d9",
			2658 => x"febd29d9",
			2659 => x"0601a324",
			2660 => x"03067808",
			2661 => x"05060604",
			2662 => x"000029d9",
			2663 => x"01bf29d9",
			2664 => x"06016b0c",
			2665 => x"0c052a04",
			2666 => x"000029d9",
			2667 => x"0c056304",
			2668 => x"fdf329d9",
			2669 => x"000029d9",
			2670 => x"01009f08",
			2671 => x"04110304",
			2672 => x"fecc29d9",
			2673 => x"00ac29d9",
			2674 => x"0100de04",
			2675 => x"016d29d9",
			2676 => x"005629d9",
			2677 => x"fe7829d9",
			2678 => x"0b053504",
			2679 => x"fe882a65",
			2680 => x"0f07490c",
			2681 => x"0f070104",
			2682 => x"00002a65",
			2683 => x"040c2404",
			2684 => x"00002a65",
			2685 => x"029f2a65",
			2686 => x"09014318",
			2687 => x"04120c10",
			2688 => x"0f078704",
			2689 => x"00002a65",
			2690 => x"09011304",
			2691 => x"feb12a65",
			2692 => x"09014004",
			2693 => x"00002a65",
			2694 => x"ff0f2a65",
			2695 => x"0506e204",
			2696 => x"00ad2a65",
			2697 => x"00002a65",
			2698 => x"0100e210",
			2699 => x"06016b04",
			2700 => x"ffec2a65",
			2701 => x"00049c08",
			2702 => x"0506d204",
			2703 => x"00002a65",
			2704 => x"012d2a65",
			2705 => x"00002a65",
			2706 => x"0100fa0c",
			2707 => x"0d075504",
			2708 => x"ff192a65",
			2709 => x"040c7f04",
			2710 => x"00002a65",
			2711 => x"00cc2a65",
			2712 => x"ff002a65",
			2713 => x"01007e04",
			2714 => x"fe832b01",
			2715 => x"0c052820",
			2716 => x"0c04ee08",
			2717 => x"04100804",
			2718 => x"fee62b01",
			2719 => x"00002b01",
			2720 => x"0c050c10",
			2721 => x"00040204",
			2722 => x"00002b01",
			2723 => x"0a029304",
			2724 => x"02152b01",
			2725 => x"0a02be04",
			2726 => x"00002b01",
			2727 => x"010e2b01",
			2728 => x"040e6304",
			2729 => x"ff482b01",
			2730 => x"01062b01",
			2731 => x"0506b910",
			2732 => x"0803e60c",
			2733 => x"0c054c08",
			2734 => x"0209d404",
			2735 => x"00002b01",
			2736 => x"fe122b01",
			2737 => x"00002b01",
			2738 => x"00062b01",
			2739 => x"040c4404",
			2740 => x"fed52b01",
			2741 => x"0a02b30c",
			2742 => x"0100fa08",
			2743 => x"0b060904",
			2744 => x"00002b01",
			2745 => x"01342b01",
			2746 => x"00002b01",
			2747 => x"00048e04",
			2748 => x"ff312b01",
			2749 => x"0c059e04",
			2750 => x"00e82b01",
			2751 => x"ff7f2b01",
			2752 => x"0d05f704",
			2753 => x"fe712ba5",
			2754 => x"0c050c1c",
			2755 => x"0e05960c",
			2756 => x"040c2404",
			2757 => x"00002ba5",
			2758 => x"03063204",
			2759 => x"01cd2ba5",
			2760 => x"00002ba5",
			2761 => x"0c050a08",
			2762 => x"04100804",
			2763 => x"fe9d2ba5",
			2764 => x"003e2ba5",
			2765 => x"09010604",
			2766 => x"00002ba5",
			2767 => x"02142ba5",
			2768 => x"0b058710",
			2769 => x"0b058508",
			2770 => x"00051504",
			2771 => x"ff402ba5",
			2772 => x"00002ba5",
			2773 => x"01009204",
			2774 => x"00002ba5",
			2775 => x"f0e22ba5",
			2776 => x"0c05dc20",
			2777 => x"0100bc10",
			2778 => x"0803d008",
			2779 => x"020a0604",
			2780 => x"00002ba5",
			2781 => x"fe1b2ba5",
			2782 => x"01008204",
			2783 => x"ff1b2ba5",
			2784 => x"01242ba5",
			2785 => x"0a028e08",
			2786 => x"0209dd04",
			2787 => x"ff162ba5",
			2788 => x"00002ba5",
			2789 => x"0209c904",
			2790 => x"01422ba5",
			2791 => x"003f2ba5",
			2792 => x"feb12ba5",
			2793 => x"040c2404",
			2794 => x"fe812c51",
			2795 => x"08036838",
			2796 => x"08036120",
			2797 => x"08034418",
			2798 => x"040ce10c",
			2799 => x"0e0a2a08",
			2800 => x"0a028304",
			2801 => x"00002c51",
			2802 => x"01402c51",
			2803 => x"00002c51",
			2804 => x"0209c108",
			2805 => x"0f08a304",
			2806 => x"00002c51",
			2807 => x"006f2c51",
			2808 => x"ff652c51",
			2809 => x"040df504",
			2810 => x"ff6a2c51",
			2811 => x"00002c51",
			2812 => x"0f071708",
			2813 => x"040c8504",
			2814 => x"00002c51",
			2815 => x"06852c51",
			2816 => x"0100e00c",
			2817 => x"040c6604",
			2818 => x"00002c51",
			2819 => x"0505cc04",
			2820 => x"00002c51",
			2821 => x"018e2c51",
			2822 => x"00002c51",
			2823 => x"04120c10",
			2824 => x"09014104",
			2825 => x"fef02c51",
			2826 => x"0100df08",
			2827 => x"0f0ad104",
			2828 => x"00652c51",
			2829 => x"00002c51",
			2830 => x"fffc2c51",
			2831 => x"0900b104",
			2832 => x"ff6a2c51",
			2833 => x"020ac304",
			2834 => x"00ce2c51",
			2835 => x"00002c51",
			2836 => x"0d05f704",
			2837 => x"fe902cfd",
			2838 => x"0f08dd3c",
			2839 => x"07051f18",
			2840 => x"06016c10",
			2841 => x"00040204",
			2842 => x"00002cfd",
			2843 => x"0a02ae08",
			2844 => x"07050404",
			2845 => x"00002cfd",
			2846 => x"02052cfd",
			2847 => x"00002cfd",
			2848 => x"00059f04",
			2849 => x"ffea2cfd",
			2850 => x"00002cfd",
			2851 => x"06016f14",
			2852 => x"0c052e0c",
			2853 => x"00043e04",
			2854 => x"ffa12cfd",
			2855 => x"05060804",
			2856 => x"00002cfd",
			2857 => x"00ba2cfd",
			2858 => x"06016804",
			2859 => x"fee32cfd",
			2860 => x"00002cfd",
			2861 => x"040d8804",
			2862 => x"00002cfd",
			2863 => x"0b061908",
			2864 => x"08034804",
			2865 => x"00002cfd",
			2866 => x"014d2cfd",
			2867 => x"00002cfd",
			2868 => x"05070d08",
			2869 => x"0f08e604",
			2870 => x"00002cfd",
			2871 => x"fe9d2cfd",
			2872 => x"0c05dc0c",
			2873 => x"040c7f04",
			2874 => x"00002cfd",
			2875 => x"0d079604",
			2876 => x"00002cfd",
			2877 => x"00f42cfd",
			2878 => x"ff672cfd",
			2879 => x"07050408",
			2880 => x"08044304",
			2881 => x"ff062d99",
			2882 => x"00002d99",
			2883 => x"07051a14",
			2884 => x"0208dd10",
			2885 => x"0e050004",
			2886 => x"00002d99",
			2887 => x"08032804",
			2888 => x"00002d99",
			2889 => x"0d05f704",
			2890 => x"00002d99",
			2891 => x"017f2d99",
			2892 => x"00002d99",
			2893 => x"040c4404",
			2894 => x"ff402d99",
			2895 => x"00041410",
			2896 => x"0c056204",
			2897 => x"00002d99",
			2898 => x"0100fa08",
			2899 => x"0506e204",
			2900 => x"00002d99",
			2901 => x"00b42d99",
			2902 => x"00002d99",
			2903 => x"06017010",
			2904 => x"0c054808",
			2905 => x"040e2304",
			2906 => x"00002d99",
			2907 => x"00c32d99",
			2908 => x"06016b04",
			2909 => x"ff9b2d99",
			2910 => x"00002d99",
			2911 => x"04100808",
			2912 => x"03099604",
			2913 => x"ff452d99",
			2914 => x"00002d99",
			2915 => x"08046104",
			2916 => x"000a2d99",
			2917 => x"00002d99",
			2918 => x"0d05f704",
			2919 => x"fe6e2e45",
			2920 => x"0c05282c",
			2921 => x"0c050714",
			2922 => x"0e05960c",
			2923 => x"040d2e04",
			2924 => x"fff92e45",
			2925 => x"06017804",
			2926 => x"01d32e45",
			2927 => x"00002e45",
			2928 => x"04100804",
			2929 => x"fe8f2e45",
			2930 => x"00002e45",
			2931 => x"00040304",
			2932 => x"fff42e45",
			2933 => x"0a029304",
			2934 => x"02f22e45",
			2935 => x"00047808",
			2936 => x"00045f04",
			2937 => x"ffcd2e45",
			2938 => x"00002e45",
			2939 => x"01007e04",
			2940 => x"00002e45",
			2941 => x"018d2e45",
			2942 => x"06016608",
			2943 => x"0c052e04",
			2944 => x"00002e45",
			2945 => x"fe3f2e45",
			2946 => x"0100fa1c",
			2947 => x"00043e0c",
			2948 => x"0506d504",
			2949 => x"ff7b2e45",
			2950 => x"0a028d04",
			2951 => x"00002e45",
			2952 => x"015c2e45",
			2953 => x"0f094508",
			2954 => x"0004dd04",
			2955 => x"ff712e45",
			2956 => x"01372e45",
			2957 => x"0100dc04",
			2958 => x"fe822e45",
			2959 => x"00002e45",
			2960 => x"fe8b2e45",
			2961 => x"0d05f704",
			2962 => x"fe702ed1",
			2963 => x"08031d04",
			2964 => x"fe8d2ed1",
			2965 => x"0a029318",
			2966 => x"0c050704",
			2967 => x"ffa52ed1",
			2968 => x"0209be08",
			2969 => x"08032804",
			2970 => x"00002ed1",
			2971 => x"02182ed1",
			2972 => x"0307f404",
			2973 => x"00002ed1",
			2974 => x"030a6904",
			2975 => x"01062ed1",
			2976 => x"00002ed1",
			2977 => x"0e05c314",
			2978 => x"0c05450c",
			2979 => x"040d2e04",
			2980 => x"ffa52ed1",
			2981 => x"01006704",
			2982 => x"00002ed1",
			2983 => x"018c2ed1",
			2984 => x"01008404",
			2985 => x"fedf2ed1",
			2986 => x"00002ed1",
			2987 => x"0d069408",
			2988 => x"0410e104",
			2989 => x"fe5a2ed1",
			2990 => x"00002ed1",
			2991 => x"0c05dc08",
			2992 => x"0c058004",
			2993 => x"fffd2ed1",
			2994 => x"00fa2ed1",
			2995 => x"fe9c2ed1",
			2996 => x"0d05f704",
			2997 => x"feac2f7d",
			2998 => x"08036830",
			2999 => x"0003f708",
			3000 => x"040c4404",
			3001 => x"ff342f7d",
			3002 => x"00002f7d",
			3003 => x"00040710",
			3004 => x"0a029b0c",
			3005 => x"05061504",
			3006 => x"00002f7d",
			3007 => x"0100fa04",
			3008 => x"01a72f7d",
			3009 => x"00002f7d",
			3010 => x"00002f7d",
			3011 => x"00046710",
			3012 => x"0a029008",
			3013 => x"0c056204",
			3014 => x"00002f7d",
			3015 => x"00cb2f7d",
			3016 => x"0c058004",
			3017 => x"ff3d2f7d",
			3018 => x"00002f7d",
			3019 => x"09016304",
			3020 => x"016b2f7d",
			3021 => x"00002f7d",
			3022 => x"06018820",
			3023 => x"0100ca18",
			3024 => x"0900e70c",
			3025 => x"0305e904",
			3026 => x"00002f7d",
			3027 => x"0005b004",
			3028 => x"ff432f7d",
			3029 => x"00002f7d",
			3030 => x"040eab04",
			3031 => x"00002f7d",
			3032 => x"06016b04",
			3033 => x"00002f7d",
			3034 => x"01062f7d",
			3035 => x"06017804",
			3036 => x"ff3f2f7d",
			3037 => x"00002f7d",
			3038 => x"fedc2f7d",
			3039 => x"0b053504",
			3040 => x"fe76300b",
			3041 => x"040baa04",
			3042 => x"fe94300b",
			3043 => x"08036818",
			3044 => x"0100fa14",
			3045 => x"02089f04",
			3046 => x"022f300b",
			3047 => x"0d071608",
			3048 => x"00046804",
			3049 => x"fef7300b",
			3050 => x"0000300b",
			3051 => x"0e073b04",
			3052 => x"0000300b",
			3053 => x"017a300b",
			3054 => x"ff4b300b",
			3055 => x"0c054810",
			3056 => x"040e2304",
			3057 => x"fecd300b",
			3058 => x"020a8608",
			3059 => x"0c052e04",
			3060 => x"0176300b",
			3061 => x"0000300b",
			3062 => x"ff80300b",
			3063 => x"0d06af0c",
			3064 => x"05067e08",
			3065 => x"0b05b704",
			3066 => x"fdb8300b",
			3067 => x"0000300b",
			3068 => x"0000300b",
			3069 => x"0c059e08",
			3070 => x"00049604",
			3071 => x"ffa1300b",
			3072 => x"011f300b",
			3073 => x"ff11300b",
			3074 => x"0000300d",
			3075 => x"00003011",
			3076 => x"00003015",
			3077 => x"00003019",
			3078 => x"0000301d",
			3079 => x"00003021",
			3080 => x"00003025",
			3081 => x"00003029",
			3082 => x"0000302d",
			3083 => x"040c2404",
			3084 => x"ffdd3039",
			3085 => x"00003039",
			3086 => x"06016b04",
			3087 => x"ffe6304d",
			3088 => x"06019004",
			3089 => x"0008304d",
			3090 => x"0000304d",
			3091 => x"0100bd04",
			3092 => x"ffff3061",
			3093 => x"0100f304",
			3094 => x"00063061",
			3095 => x"00003061",
			3096 => x"03071b08",
			3097 => x"06017304",
			3098 => x"ffdd3075",
			3099 => x"00003075",
			3100 => x"00003075",
			3101 => x"0e078e08",
			3102 => x"04100804",
			3103 => x"ffc43089",
			3104 => x"00003089",
			3105 => x"00003089",
			3106 => x"0e055a04",
			3107 => x"0000309d",
			3108 => x"0e0a2a04",
			3109 => x"0010309d",
			3110 => x"0000309d",
			3111 => x"0f08dd08",
			3112 => x"0f070104",
			3113 => x"000030b9",
			3114 => x"001e30b9",
			3115 => x"0f0abc04",
			3116 => x"ffe030b9",
			3117 => x"000030b9",
			3118 => x"02086004",
			3119 => x"000030d5",
			3120 => x"0e097708",
			3121 => x"00048604",
			3122 => x"ff6830d5",
			3123 => x"000030d5",
			3124 => x"000030d5",
			3125 => x"02086004",
			3126 => x"000030f1",
			3127 => x"040d5508",
			3128 => x"0f0abc04",
			3129 => x"ff7530f1",
			3130 => x"000030f1",
			3131 => x"000030f1",
			3132 => x"0100dc0c",
			3133 => x"01006704",
			3134 => x"0000310d",
			3135 => x"0100c904",
			3136 => x"0028310d",
			3137 => x"0000310d",
			3138 => x"ffff310d",
			3139 => x"0306ff04",
			3140 => x"ffee3129",
			3141 => x"09018708",
			3142 => x"09010604",
			3143 => x"00003129",
			3144 => x"00153129",
			3145 => x"00003129",
			3146 => x"0c052808",
			3147 => x"0d064504",
			3148 => x"0000314d",
			3149 => x"000d314d",
			3150 => x"0f0abc08",
			3151 => x"07054904",
			3152 => x"0000314d",
			3153 => x"ffde314d",
			3154 => x"0000314d",
			3155 => x"0f08c608",
			3156 => x"0f070104",
			3157 => x"00003171",
			3158 => x"00023171",
			3159 => x"0f0aed08",
			3160 => x"0f08dd04",
			3161 => x"00003171",
			3162 => x"ffd53171",
			3163 => x"00003171",
			3164 => x"0c050c0c",
			3165 => x"07050104",
			3166 => x"0000319d",
			3167 => x"0b052404",
			3168 => x"0000319d",
			3169 => x"0013319d",
			3170 => x"030a5c08",
			3171 => x"07054904",
			3172 => x"0000319d",
			3173 => x"ffdd319d",
			3174 => x"0000319d",
			3175 => x"040dca0c",
			3176 => x"02085b04",
			3177 => x"000031c9",
			3178 => x"020b0f04",
			3179 => x"ff8c31c9",
			3180 => x"000031c9",
			3181 => x"0d06c704",
			3182 => x"000031c9",
			3183 => x"0d083204",
			3184 => x"001d31c9",
			3185 => x"000031c9",
			3186 => x"02086004",
			3187 => x"000031ed",
			3188 => x"040e630c",
			3189 => x"0f0abc08",
			3190 => x"0f071f04",
			3191 => x"000031ed",
			3192 => x"ff5d31ed",
			3193 => x"000031ed",
			3194 => x"000031ed",
			3195 => x"0c052810",
			3196 => x"01006704",
			3197 => x"00003211",
			3198 => x"0100d008",
			3199 => x"0c04b204",
			3200 => x"00003211",
			3201 => x"00463211",
			3202 => x"00003211",
			3203 => x"fffe3211",
			3204 => x"0506e210",
			3205 => x"04120c0c",
			3206 => x"02088304",
			3207 => x"00003235",
			3208 => x"0f071d04",
			3209 => x"00003235",
			3210 => x"ffa93235",
			3211 => x"00003235",
			3212 => x"00003235",
			3213 => x"00046708",
			3214 => x"00040304",
			3215 => x"00003261",
			3216 => x"ffd33261",
			3217 => x"0803820c",
			3218 => x"07050404",
			3219 => x"00003261",
			3220 => x"0705bb04",
			3221 => x"00523261",
			3222 => x"00003261",
			3223 => x"00003261",
			3224 => x"0004670c",
			3225 => x"00040304",
			3226 => x"00003295",
			3227 => x"040da904",
			3228 => x"ffd13295",
			3229 => x"00003295",
			3230 => x"0803820c",
			3231 => x"07050404",
			3232 => x"00003295",
			3233 => x"0705bb04",
			3234 => x"00493295",
			3235 => x"00003295",
			3236 => x"00003295",
			3237 => x"0004140c",
			3238 => x"0a028d04",
			3239 => x"000032c9",
			3240 => x"0a029b04",
			3241 => x"001232c9",
			3242 => x"000032c9",
			3243 => x"0a028504",
			3244 => x"000032c9",
			3245 => x"0005b808",
			3246 => x"0c058004",
			3247 => x"ffdf32c9",
			3248 => x"000032c9",
			3249 => x"000032c9",
			3250 => x"0506e210",
			3251 => x"04120c0c",
			3252 => x"02088304",
			3253 => x"000032fd",
			3254 => x"0f071d04",
			3255 => x"000032fd",
			3256 => x"ffb332fd",
			3257 => x"000032fd",
			3258 => x"0c05dc08",
			3259 => x"0c056204",
			3260 => x"000032fd",
			3261 => x"001032fd",
			3262 => x"000032fd",
			3263 => x"040e2310",
			3264 => x"0a029004",
			3265 => x"00003339",
			3266 => x"0f071704",
			3267 => x"00003339",
			3268 => x"0003fb04",
			3269 => x"00003339",
			3270 => x"ff9d3339",
			3271 => x"0100c90c",
			3272 => x"01007304",
			3273 => x"00003339",
			3274 => x"0f09a304",
			3275 => x"002c3339",
			3276 => x"00003339",
			3277 => x"00003339",
			3278 => x"0100dc14",
			3279 => x"01006704",
			3280 => x"00003365",
			3281 => x"00040204",
			3282 => x"00003365",
			3283 => x"0a02fd08",
			3284 => x"0a027f04",
			3285 => x"00003365",
			3286 => x"00423365",
			3287 => x"00003365",
			3288 => x"00003365",
			3289 => x"06016608",
			3290 => x"040c2404",
			3291 => x"ffdf33a1",
			3292 => x"000033a1",
			3293 => x"06017410",
			3294 => x"01009b04",
			3295 => x"000033a1",
			3296 => x"0100f308",
			3297 => x"040adc04",
			3298 => x"000033a1",
			3299 => x"005333a1",
			3300 => x"000033a1",
			3301 => x"040fc604",
			3302 => x"fff133a1",
			3303 => x"000033a1",
			3304 => x"0901411c",
			3305 => x"0208910c",
			3306 => x"03060104",
			3307 => x"000033ed",
			3308 => x"0e060004",
			3309 => x"001d33ed",
			3310 => x"000033ed",
			3311 => x"04120c0c",
			3312 => x"0f073b04",
			3313 => x"000033ed",
			3314 => x"05070d04",
			3315 => x"ff7b33ed",
			3316 => x"000033ed",
			3317 => x"000033ed",
			3318 => x"0100e208",
			3319 => x"09015304",
			3320 => x"000033ed",
			3321 => x"002933ed",
			3322 => x"000033ed",
			3323 => x"0c052818",
			3324 => x"0c04d004",
			3325 => x"00003431",
			3326 => x"040adc04",
			3327 => x"00003431",
			3328 => x"0305f004",
			3329 => x"00003431",
			3330 => x"020a8608",
			3331 => x"03087504",
			3332 => x"004c3431",
			3333 => x"00003431",
			3334 => x"00003431",
			3335 => x"020a6308",
			3336 => x"0209c904",
			3337 => x"00003431",
			3338 => x"ffd23431",
			3339 => x"00003431",
			3340 => x"0901060c",
			3341 => x"0f074904",
			3342 => x"0000347d",
			3343 => x"0803fa04",
			3344 => x"ffa9347d",
			3345 => x"0000347d",
			3346 => x"06019714",
			3347 => x"0a028d04",
			3348 => x"0000347d",
			3349 => x"06016b04",
			3350 => x"0000347d",
			3351 => x"09016108",
			3352 => x"0c050a04",
			3353 => x"0000347d",
			3354 => x"00d2347d",
			3355 => x"0000347d",
			3356 => x"0a029b04",
			3357 => x"0000347d",
			3358 => x"fffc347d",
			3359 => x"0900b704",
			3360 => x"000034b1",
			3361 => x"040c2404",
			3362 => x"000034b1",
			3363 => x"0901a110",
			3364 => x"0410bb0c",
			3365 => x"030a7808",
			3366 => x"0b053504",
			3367 => x"000034b1",
			3368 => x"004634b1",
			3369 => x"000034b1",
			3370 => x"000034b1",
			3371 => x"000034b1",
			3372 => x"00040718",
			3373 => x"08031d04",
			3374 => x"000034fd",
			3375 => x"0100fa10",
			3376 => x"0d063804",
			3377 => x"000034fd",
			3378 => x"08033108",
			3379 => x"040adc04",
			3380 => x"000034fd",
			3381 => x"00ba34fd",
			3382 => x"000034fd",
			3383 => x"000034fd",
			3384 => x"0100bc0c",
			3385 => x"04120c08",
			3386 => x"0f079d04",
			3387 => x"000034fd",
			3388 => x"ff8434fd",
			3389 => x"000034fd",
			3390 => x"000034fd",
			3391 => x"040cce0c",
			3392 => x"02083d04",
			3393 => x"00003551",
			3394 => x"07069b04",
			3395 => x"ff563551",
			3396 => x"00003551",
			3397 => x"08038814",
			3398 => x"0100f310",
			3399 => x"0004a70c",
			3400 => x"01006704",
			3401 => x"00003551",
			3402 => x"08032804",
			3403 => x"00003551",
			3404 => x"00733551",
			3405 => x"00003551",
			3406 => x"00003551",
			3407 => x"04100804",
			3408 => x"ffbd3551",
			3409 => x"04143604",
			3410 => x"00053551",
			3411 => x"00003551",
			3412 => x"040cce0c",
			3413 => x"02083d04",
			3414 => x"000035a5",
			3415 => x"06019604",
			3416 => x"ff4335a5",
			3417 => x"000035a5",
			3418 => x"0601891c",
			3419 => x"0d06d410",
			3420 => x"0f082208",
			3421 => x"03055f04",
			3422 => x"000035a5",
			3423 => x"000e35a5",
			3424 => x"0e05c304",
			3425 => x"000035a5",
			3426 => x"fff035a5",
			3427 => x"0c059e08",
			3428 => x"08032804",
			3429 => x"000035a5",
			3430 => x"009a35a5",
			3431 => x"000035a5",
			3432 => x"000035a5",
			3433 => x"0803661c",
			3434 => x"0b053504",
			3435 => x"000035f1",
			3436 => x"08031d04",
			3437 => x"000035f1",
			3438 => x"0100fa10",
			3439 => x"0a02b30c",
			3440 => x"0c04d004",
			3441 => x"000035f1",
			3442 => x"040adc04",
			3443 => x"000035f1",
			3444 => x"006635f1",
			3445 => x"000035f1",
			3446 => x"000035f1",
			3447 => x"04120c08",
			3448 => x"0b066c04",
			3449 => x"ffb735f1",
			3450 => x"000035f1",
			3451 => x"000035f1",
			3452 => x"07058c1c",
			3453 => x"0b053504",
			3454 => x"0000363d",
			3455 => x"0100cb14",
			3456 => x"00040204",
			3457 => x"0000363d",
			3458 => x"01006f04",
			3459 => x"0000363d",
			3460 => x"020a8608",
			3461 => x"0c04d004",
			3462 => x"0000363d",
			3463 => x"0054363d",
			3464 => x"0000363d",
			3465 => x"0000363d",
			3466 => x"00040304",
			3467 => x"0000363d",
			3468 => x"0209e804",
			3469 => x"0000363d",
			3470 => x"ff8e363d",
			3471 => x"0f08dd1c",
			3472 => x"07050404",
			3473 => x"00003681",
			3474 => x"08032504",
			3475 => x"00003681",
			3476 => x"0c052810",
			3477 => x"0705750c",
			3478 => x"08046108",
			3479 => x"0c04b204",
			3480 => x"00003681",
			3481 => x"00543681",
			3482 => x"00003681",
			3483 => x"00003681",
			3484 => x"00003681",
			3485 => x"0c050b04",
			3486 => x"00003681",
			3487 => x"ffd13681",
			3488 => x"07058c1c",
			3489 => x"0d05f704",
			3490 => x"ffa036d5",
			3491 => x"06018e14",
			3492 => x"00040304",
			3493 => x"000036d5",
			3494 => x"01006704",
			3495 => x"000036d5",
			3496 => x"08032804",
			3497 => x"000036d5",
			3498 => x"07050104",
			3499 => x"000036d5",
			3500 => x"009736d5",
			3501 => x"000036d5",
			3502 => x"0d07550c",
			3503 => x"0b05e504",
			3504 => x"000036d5",
			3505 => x"0209b104",
			3506 => x"000036d5",
			3507 => x"ff5a36d5",
			3508 => x"000036d5",
			3509 => x"09015324",
			3510 => x"02089118",
			3511 => x"03060104",
			3512 => x"00003729",
			3513 => x"0e060010",
			3514 => x"0b053504",
			3515 => x"00003729",
			3516 => x"0b056508",
			3517 => x"0c050904",
			3518 => x"00333729",
			3519 => x"00003729",
			3520 => x"00003729",
			3521 => x"00003729",
			3522 => x"04120c08",
			3523 => x"0e04f704",
			3524 => x"00003729",
			3525 => x"ff793729",
			3526 => x"00003729",
			3527 => x"0100e204",
			3528 => x"00313729",
			3529 => x"00003729",
			3530 => x"0209ce1c",
			3531 => x"0900b704",
			3532 => x"0000377d",
			3533 => x"00040204",
			3534 => x"0000377d",
			3535 => x"0b053504",
			3536 => x"0000377d",
			3537 => x"0601710c",
			3538 => x"07050404",
			3539 => x"0000377d",
			3540 => x"0d05f704",
			3541 => x"0000377d",
			3542 => x"0073377d",
			3543 => x"0000377d",
			3544 => x"0f0abc0c",
			3545 => x"04120c08",
			3546 => x"00040304",
			3547 => x"0000377d",
			3548 => x"ff78377d",
			3549 => x"0000377d",
			3550 => x"0000377d",
			3551 => x"0705a91c",
			3552 => x"0d05f704",
			3553 => x"000037b9",
			3554 => x"0a02c314",
			3555 => x"00040204",
			3556 => x"000037b9",
			3557 => x"07050404",
			3558 => x"000037b9",
			3559 => x"0f09b108",
			3560 => x"08032504",
			3561 => x"000037b9",
			3562 => x"007537b9",
			3563 => x"000037b9",
			3564 => x"000037b9",
			3565 => x"ffd137b9",
			3566 => x"01008e04",
			3567 => x"000037f5",
			3568 => x"0100fa18",
			3569 => x"0a027f04",
			3570 => x"000037f5",
			3571 => x"07050504",
			3572 => x"000037f5",
			3573 => x"0d063804",
			3574 => x"000037f5",
			3575 => x"0b073308",
			3576 => x"05061504",
			3577 => x"000037f5",
			3578 => x"004537f5",
			3579 => x"000037f5",
			3580 => x"000037f5",
			3581 => x"0e055a04",
			3582 => x"00003831",
			3583 => x"0f09b118",
			3584 => x"0100dc14",
			3585 => x"0a027f04",
			3586 => x"00003831",
			3587 => x"0900b704",
			3588 => x"00003831",
			3589 => x"09016308",
			3590 => x"06018e04",
			3591 => x"005a3831",
			3592 => x"00003831",
			3593 => x"00003831",
			3594 => x"00003831",
			3595 => x"00003831",
			3596 => x"040c2404",
			3597 => x"ff3e388d",
			3598 => x"08036610",
			3599 => x"07050404",
			3600 => x"0000388d",
			3601 => x"020b5b08",
			3602 => x"08031d04",
			3603 => x"0000388d",
			3604 => x"004c388d",
			3605 => x"0000388d",
			3606 => x"06018814",
			3607 => x"040eab08",
			3608 => x"020a2004",
			3609 => x"fffe388d",
			3610 => x"0000388d",
			3611 => x"06016a04",
			3612 => x"0000388d",
			3613 => x"00064804",
			3614 => x"006e388d",
			3615 => x"0000388d",
			3616 => x"0d07ee04",
			3617 => x"ff88388d",
			3618 => x"0000388d",
			3619 => x"0209ce1c",
			3620 => x"0900b704",
			3621 => x"000038e9",
			3622 => x"00040204",
			3623 => x"000038e9",
			3624 => x"0b053504",
			3625 => x"000038e9",
			3626 => x"0601710c",
			3627 => x"08032504",
			3628 => x"000038e9",
			3629 => x"07050404",
			3630 => x"000038e9",
			3631 => x"006138e9",
			3632 => x"000038e9",
			3633 => x"0c052804",
			3634 => x"000038e9",
			3635 => x"0f0abc0c",
			3636 => x"00040304",
			3637 => x"000038e9",
			3638 => x"0005b804",
			3639 => x"ff7a38e9",
			3640 => x"000038e9",
			3641 => x"000038e9",
			3642 => x"00040718",
			3643 => x"08031d04",
			3644 => x"ffd2395d",
			3645 => x"0c04ee04",
			3646 => x"0000395d",
			3647 => x"0100fa0c",
			3648 => x"08033608",
			3649 => x"040adc04",
			3650 => x"0000395d",
			3651 => x"014d395d",
			3652 => x"0000395d",
			3653 => x"0000395d",
			3654 => x"02086008",
			3655 => x"0305e104",
			3656 => x"ffe5395d",
			3657 => x"00e7395d",
			3658 => x"040d4204",
			3659 => x"fef8395d",
			3660 => x"0209ce0c",
			3661 => x"05062304",
			3662 => x"0000395d",
			3663 => x"0e052004",
			3664 => x"0000395d",
			3665 => x"006f395d",
			3666 => x"0005b808",
			3667 => x"0506e204",
			3668 => x"ff44395d",
			3669 => x"0000395d",
			3670 => x"0000395d",
			3671 => x"00040718",
			3672 => x"08031d04",
			3673 => x"ffd939d1",
			3674 => x"0c04ee04",
			3675 => x"000039d1",
			3676 => x"0100fa0c",
			3677 => x"08033608",
			3678 => x"040adc04",
			3679 => x"000039d1",
			3680 => x"013b39d1",
			3681 => x"000039d1",
			3682 => x"000039d1",
			3683 => x"02086008",
			3684 => x"0305e104",
			3685 => x"ffea39d1",
			3686 => x"00dc39d1",
			3687 => x"040d4204",
			3688 => x"ff0439d1",
			3689 => x"0209ce08",
			3690 => x"01008a04",
			3691 => x"000039d1",
			3692 => x"007039d1",
			3693 => x"0005b80c",
			3694 => x"0506e208",
			3695 => x"0f07d504",
			3696 => x"000039d1",
			3697 => x"ff5539d1",
			3698 => x"000039d1",
			3699 => x"000039d1",
			3700 => x"02086010",
			3701 => x"07050404",
			3702 => x"00003a55",
			3703 => x"0e050004",
			3704 => x"00003a55",
			3705 => x"08032504",
			3706 => x"00003a55",
			3707 => x"00f93a55",
			3708 => x"00040718",
			3709 => x"0a028e04",
			3710 => x"00003a55",
			3711 => x"0100ff10",
			3712 => x"03071b04",
			3713 => x"00003a55",
			3714 => x"08033608",
			3715 => x"040ad504",
			3716 => x"00003a55",
			3717 => x"00ad3a55",
			3718 => x"00003a55",
			3719 => x"00003a55",
			3720 => x"0410080c",
			3721 => x"0b05fa08",
			3722 => x"02086704",
			3723 => x"00003a55",
			3724 => x"ff323a55",
			3725 => x"00003a55",
			3726 => x"0a03630c",
			3727 => x"0b063908",
			3728 => x"06015604",
			3729 => x"00003a55",
			3730 => x"00793a55",
			3731 => x"00003a55",
			3732 => x"fffe3a55",
			3733 => x"040c2404",
			3734 => x"ff2b3ab9",
			3735 => x"08036618",
			3736 => x"0100fa14",
			3737 => x"01006704",
			3738 => x"00003ab9",
			3739 => x"0a02b30c",
			3740 => x"0a028e04",
			3741 => x"00003ab9",
			3742 => x"0d05f704",
			3743 => x"00003ab9",
			3744 => x"008c3ab9",
			3745 => x"00003ab9",
			3746 => x"00003ab9",
			3747 => x"06018810",
			3748 => x"06016a04",
			3749 => x"00003ab9",
			3750 => x"040eab04",
			3751 => x"00003ab9",
			3752 => x"01007304",
			3753 => x"00003ab9",
			3754 => x"007e3ab9",
			3755 => x"0d07ee04",
			3756 => x"ff7b3ab9",
			3757 => x"00003ab9",
			3758 => x"0f08dd34",
			3759 => x"07050408",
			3760 => x"0a034104",
			3761 => x"ff5e3b3d",
			3762 => x"00003b3d",
			3763 => x"07051a14",
			3764 => x"0208dd10",
			3765 => x"0a028304",
			3766 => x"00003b3d",
			3767 => x"0d05f704",
			3768 => x"00003b3d",
			3769 => x"06016c04",
			3770 => x"00fd3b3d",
			3771 => x"00003b3d",
			3772 => x"00003b3d",
			3773 => x"040d4208",
			3774 => x"02088304",
			3775 => x"00003b3d",
			3776 => x"ff9f3b3d",
			3777 => x"01007c04",
			3778 => x"00003b3d",
			3779 => x"06016604",
			3780 => x"00003b3d",
			3781 => x"0705ce04",
			3782 => x"00933b3d",
			3783 => x"00003b3d",
			3784 => x"09015a08",
			3785 => x"0f08f004",
			3786 => x"00003b3d",
			3787 => x"ff153b3d",
			3788 => x"0100e704",
			3789 => x"00563b3d",
			3790 => x"ff9c3b3d",
			3791 => x"0100bc1c",
			3792 => x"0f085c18",
			3793 => x"0d05f704",
			3794 => x"00003ba9",
			3795 => x"0c054610",
			3796 => x"0a028304",
			3797 => x"00003ba9",
			3798 => x"06018008",
			3799 => x"03055f04",
			3800 => x"00003ba9",
			3801 => x"007f3ba9",
			3802 => x"00003ba9",
			3803 => x"00003ba9",
			3804 => x"ffb23ba9",
			3805 => x"0a028d04",
			3806 => x"00003ba9",
			3807 => x"0100fa14",
			3808 => x"0d06e204",
			3809 => x"00003ba9",
			3810 => x"020b690c",
			3811 => x"0601a608",
			3812 => x"040c4404",
			3813 => x"00003ba9",
			3814 => x"009e3ba9",
			3815 => x"00003ba9",
			3816 => x"00003ba9",
			3817 => x"00003ba9",
			3818 => x"0505f908",
			3819 => x"04100804",
			3820 => x"feef3c1d",
			3821 => x"00003c1d",
			3822 => x"0c050c10",
			3823 => x"0c04ed04",
			3824 => x"00003c1d",
			3825 => x"0f09b108",
			3826 => x"08032504",
			3827 => x"00003c1d",
			3828 => x"013c3c1d",
			3829 => x"00003c1d",
			3830 => x"0a028e04",
			3831 => x"ff973c1d",
			3832 => x"07057310",
			3833 => x"0a030d0c",
			3834 => x"06016304",
			3835 => x"00003c1d",
			3836 => x"09012d04",
			3837 => x"ff9c3c1d",
			3838 => x"00003c1d",
			3839 => x"00003c1d",
			3840 => x"030a690c",
			3841 => x"06016304",
			3842 => x"00003c1d",
			3843 => x"09010a04",
			3844 => x"00003c1d",
			3845 => x"008f3c1d",
			3846 => x"00003c1d",
			3847 => x"0d05f704",
			3848 => x"fe6c3c81",
			3849 => x"0c059e20",
			3850 => x"0601911c",
			3851 => x"0003f704",
			3852 => x"fec03c81",
			3853 => x"02089108",
			3854 => x"0b056504",
			3855 => x"03553c81",
			3856 => x"ff273c81",
			3857 => x"0b056308",
			3858 => x"03060904",
			3859 => x"00ba3c81",
			3860 => x"fe913c81",
			3861 => x"0c052804",
			3862 => x"019b3c81",
			3863 => x"007a3c81",
			3864 => x"fe6f3c81",
			3865 => x"020b1c04",
			3866 => x"fe783c81",
			3867 => x"0f0b1c08",
			3868 => x"00040b04",
			3869 => x"01453c81",
			3870 => x"fff13c81",
			3871 => x"fe9a3c81",
			3872 => x"0d05f704",
			3873 => x"fed53cfd",
			3874 => x"07058c2c",
			3875 => x"08036e14",
			3876 => x"00040204",
			3877 => x"00003cfd",
			3878 => x"07050404",
			3879 => x"00003cfd",
			3880 => x"0c056308",
			3881 => x"0e088604",
			3882 => x"01593cfd",
			3883 => x"00003cfd",
			3884 => x"00003cfd",
			3885 => x"0410080c",
			3886 => x"0c051108",
			3887 => x"06016404",
			3888 => x"00003cfd",
			3889 => x"ff4b3cfd",
			3890 => x"00003cfd",
			3891 => x"06016604",
			3892 => x"00003cfd",
			3893 => x"00076604",
			3894 => x"00a23cfd",
			3895 => x"00003cfd",
			3896 => x"0209e808",
			3897 => x"0c056404",
			3898 => x"00003cfd",
			3899 => x"fff73cfd",
			3900 => x"0e05e004",
			3901 => x"00003cfd",
			3902 => x"ff363cfd",
			3903 => x"0505f908",
			3904 => x"04100804",
			3905 => x"fedf3d89",
			3906 => x"00003d89",
			3907 => x"0208dd10",
			3908 => x"0b05690c",
			3909 => x"0c050c08",
			3910 => x"00040204",
			3911 => x"00003d89",
			3912 => x"01863d89",
			3913 => x"00003d89",
			3914 => x"00003d89",
			3915 => x"07057310",
			3916 => x"0005540c",
			3917 => x"0f07c704",
			3918 => x"00003d89",
			3919 => x"09012d04",
			3920 => x"ff443d89",
			3921 => x"00003d89",
			3922 => x"00003d89",
			3923 => x"040dca10",
			3924 => x"020b0f08",
			3925 => x"0209c104",
			3926 => x"00003d89",
			3927 => x"ff6d3d89",
			3928 => x"030a6904",
			3929 => x"00883d89",
			3930 => x"00003d89",
			3931 => x"0705d10c",
			3932 => x"06016304",
			3933 => x"00003d89",
			3934 => x"08034f04",
			3935 => x"00003d89",
			3936 => x"00fc3d89",
			3937 => x"00003d89",
			3938 => x"0601661c",
			3939 => x"0900c408",
			3940 => x"0f084f04",
			3941 => x"fe663e3d",
			3942 => x"fccf3e3d",
			3943 => x"0f079d0c",
			3944 => x"08032504",
			3945 => x"fe7d3e3d",
			3946 => x"05060604",
			3947 => x"febe3e3d",
			3948 => x"05453e3d",
			3949 => x"0305e904",
			3950 => x"00d13e3d",
			3951 => x"fe553e3d",
			3952 => x"0c059e30",
			3953 => x"0209ab14",
			3954 => x"0b056504",
			3955 => x"fe733e3d",
			3956 => x"07050804",
			3957 => x"080b3e3d",
			3958 => x"00052904",
			3959 => x"fe953e3d",
			3960 => x"0e034304",
			3961 => x"ff153e3d",
			3962 => x"015a3e3d",
			3963 => x"06019018",
			3964 => x"0f097d10",
			3965 => x"0f08dd08",
			3966 => x"0e071504",
			3967 => x"01ae3e3d",
			3968 => x"03a13e3d",
			3969 => x"09018304",
			3970 => x"00223e3d",
			3971 => x"fe8d3e3d",
			3972 => x"00040204",
			3973 => x"00003e3d",
			3974 => x"04033e3d",
			3975 => x"fe2b3e3d",
			3976 => x"0e0a2a0c",
			3977 => x"030a5c04",
			3978 => x"fe6d3e3d",
			3979 => x"030a6904",
			3980 => x"02963e3d",
			3981 => x"feeb3e3d",
			3982 => x"fe663e3d",
			3983 => x"0d05f704",
			3984 => x"fede3ec1",
			3985 => x"07058c30",
			3986 => x"08036e18",
			3987 => x"00040204",
			3988 => x"00003ec1",
			3989 => x"07050404",
			3990 => x"00003ec1",
			3991 => x"07051f08",
			3992 => x"06016c04",
			3993 => x"01a13ec1",
			3994 => x"00003ec1",
			3995 => x"03079c04",
			3996 => x"fffa3ec1",
			3997 => x"00ea3ec1",
			3998 => x"0100930c",
			3999 => x"0f07d504",
			4000 => x"00003ec1",
			4001 => x"00055404",
			4002 => x"ff293ec1",
			4003 => x"00003ec1",
			4004 => x"0004c904",
			4005 => x"00003ec1",
			4006 => x"0a034404",
			4007 => x"007f3ec1",
			4008 => x"00003ec1",
			4009 => x"0209e808",
			4010 => x"0c056404",
			4011 => x"00003ec1",
			4012 => x"fffe3ec1",
			4013 => x"0b05e704",
			4014 => x"00003ec1",
			4015 => x"ff3b3ec1",
			4016 => x"0900b704",
			4017 => x"ff2e3f3d",
			4018 => x"0208dd18",
			4019 => x"0b053504",
			4020 => x"00003f3d",
			4021 => x"0c052510",
			4022 => x"08032504",
			4023 => x"00003f3d",
			4024 => x"07050404",
			4025 => x"00003f3d",
			4026 => x"06016c04",
			4027 => x"011f3f3d",
			4028 => x"00003f3d",
			4029 => x"00003f3d",
			4030 => x"0100bb08",
			4031 => x"0e068d04",
			4032 => x"00003f3d",
			4033 => x"ff183f3d",
			4034 => x"0d06e208",
			4035 => x"06018104",
			4036 => x"ffec3f3d",
			4037 => x"00003f3d",
			4038 => x"0c059e0c",
			4039 => x"08033a04",
			4040 => x"00003f3d",
			4041 => x"0100ed04",
			4042 => x"00d93f3d",
			4043 => x"00003f3d",
			4044 => x"06019604",
			4045 => x"ffed3f3d",
			4046 => x"00003f3d",
			4047 => x"040d1b24",
			4048 => x"040c2404",
			4049 => x"fe633ff1",
			4050 => x"08034114",
			4051 => x"0004240c",
			4052 => x"0100fa08",
			4053 => x"0705ba04",
			4054 => x"fedc3ff1",
			4055 => x"02563ff1",
			4056 => x"fe803ff1",
			4057 => x"0e04a004",
			4058 => x"ff763ff1",
			4059 => x"06863ff1",
			4060 => x"0b053504",
			4061 => x"fe653ff1",
			4062 => x"0505df04",
			4063 => x"025b3ff1",
			4064 => x"fe7c3ff1",
			4065 => x"0900c410",
			4066 => x"0f08160c",
			4067 => x"0900b104",
			4068 => x"fe653ff1",
			4069 => x"0e054404",
			4070 => x"01323ff1",
			4071 => x"ff353ff1",
			4072 => x"fd253ff1",
			4073 => x"07060024",
			4074 => x"0004bc14",
			4075 => x"08033f08",
			4076 => x"0705ba04",
			4077 => x"fe763ff1",
			4078 => x"03193ff1",
			4079 => x"08039008",
			4080 => x"0209c104",
			4081 => x"05d83ff1",
			4082 => x"02903ff1",
			4083 => x"00003ff1",
			4084 => x"0004dd04",
			4085 => x"ff653ff1",
			4086 => x"040f7004",
			4087 => x"feda3ff1",
			4088 => x"0a02f304",
			4089 => x"00fa3ff1",
			4090 => x"01d13ff1",
			4091 => x"fe673ff1",
			4092 => x"0d05f704",
			4093 => x"fe984075",
			4094 => x"0f079d10",
			4095 => x"0f06e304",
			4096 => x"00004075",
			4097 => x"040baa04",
			4098 => x"00004075",
			4099 => x"0c054604",
			4100 => x"01a24075",
			4101 => x"00004075",
			4102 => x"0100bb0c",
			4103 => x"04120c04",
			4104 => x"fef84075",
			4105 => x"0506e204",
			4106 => x"00674075",
			4107 => x"00004075",
			4108 => x"07058c0c",
			4109 => x"0b05d904",
			4110 => x"00004075",
			4111 => x"08033a04",
			4112 => x"00004075",
			4113 => x"017e4075",
			4114 => x"0506d20c",
			4115 => x"020a1808",
			4116 => x"0c056404",
			4117 => x"fece4075",
			4118 => x"00004075",
			4119 => x"00004075",
			4120 => x"0c05dc08",
			4121 => x"0a029904",
			4122 => x"00004075",
			4123 => x"00b84075",
			4124 => x"ff114075",
			4125 => x"07050408",
			4126 => x"0a034f04",
			4127 => x"fee94109",
			4128 => x"00004109",
			4129 => x"02086710",
			4130 => x"02083004",
			4131 => x"00004109",
			4132 => x"040baa04",
			4133 => x"00004109",
			4134 => x"07055f04",
			4135 => x"01194109",
			4136 => x"00004109",
			4137 => x"040d420c",
			4138 => x"020b0f04",
			4139 => x"ff044109",
			4140 => x"030a6904",
			4141 => x"00664109",
			4142 => x"00004109",
			4143 => x"0004bc10",
			4144 => x"0308750c",
			4145 => x"0705b808",
			4146 => x"0c057204",
			4147 => x"00f84109",
			4148 => x"00004109",
			4149 => x"00004109",
			4150 => x"00004109",
			4151 => x"04100808",
			4152 => x"09014504",
			4153 => x"ff214109",
			4154 => x"00004109",
			4155 => x"0e05e908",
			4156 => x"0c054304",
			4157 => x"00004109",
			4158 => x"ffa24109",
			4159 => x"03092204",
			4160 => x"00624109",
			4161 => x"00004109",
			4162 => x"040d1b20",
			4163 => x"040c2404",
			4164 => x"fe6241bd",
			4165 => x"08034110",
			4166 => x"030a780c",
			4167 => x"08033608",
			4168 => x"0c058204",
			4169 => x"feaa41bd",
			4170 => x"023541bd",
			4171 => x"07e341bd",
			4172 => x"fe9341bd",
			4173 => x"0d05f704",
			4174 => x"fe6341bd",
			4175 => x"03062104",
			4176 => x"03dc41bd",
			4177 => x"fe7741bd",
			4178 => x"0900c410",
			4179 => x"0f08160c",
			4180 => x"0900b104",
			4181 => x"fe6341bd",
			4182 => x"0e054404",
			4183 => x"016241bd",
			4184 => x"ff1e41bd",
			4185 => x"fcb541bd",
			4186 => x"06019128",
			4187 => x"040f0214",
			4188 => x"03066904",
			4189 => x"0e9a41bd",
			4190 => x"0307c408",
			4191 => x"0100da04",
			4192 => x"03e941bd",
			4193 => x"fe8c41bd",
			4194 => x"0506e204",
			4195 => x"238241bd",
			4196 => x"054341bd",
			4197 => x"06016608",
			4198 => x"0209c104",
			4199 => x"01bd41bd",
			4200 => x"fee341bd",
			4201 => x"0f08aa08",
			4202 => x"0a02f304",
			4203 => x"016241bd",
			4204 => x"01ed41bd",
			4205 => x"02fc41bd",
			4206 => x"fe6341bd",
			4207 => x"040d1b30",
			4208 => x"0b053504",
			4209 => x"fe674259",
			4210 => x"0d064718",
			4211 => x"0d063808",
			4212 => x"0900ba04",
			4213 => x"02c04259",
			4214 => x"fe8b4259",
			4215 => x"00040204",
			4216 => x"ff654259",
			4217 => x"00042004",
			4218 => x"18e94259",
			4219 => x"07051f04",
			4220 => x"00004259",
			4221 => x"040e4259",
			4222 => x"040c4404",
			4223 => x"fe694259",
			4224 => x"0003fb0c",
			4225 => x"01011108",
			4226 => x"08031204",
			4227 => x"00004259",
			4228 => x"02024259",
			4229 => x"fffc4259",
			4230 => x"fe9b4259",
			4231 => x"01006704",
			4232 => x"fe6c4259",
			4233 => x"0705eb18",
			4234 => x"06019114",
			4235 => x"07050408",
			4236 => x"0c04d004",
			4237 => x"feac4259",
			4238 => x"00004259",
			4239 => x"0208f704",
			4240 => x"03a34259",
			4241 => x"06016604",
			4242 => x"00004259",
			4243 => x"01804259",
			4244 => x"fe5d4259",
			4245 => x"fe584259",
			4246 => x"040d1b1c",
			4247 => x"040c2404",
			4248 => x"fe624305",
			4249 => x"0b053504",
			4250 => x"fe644305",
			4251 => x"0208bb04",
			4252 => x"073f4305",
			4253 => x"0a02a10c",
			4254 => x"0209dd04",
			4255 => x"feb04305",
			4256 => x"030a8a04",
			4257 => x"034e4305",
			4258 => x"fed94305",
			4259 => x"fe744305",
			4260 => x"0900c410",
			4261 => x"0f08160c",
			4262 => x"0900b104",
			4263 => x"fe644305",
			4264 => x"02094304",
			4265 => x"ff2d4305",
			4266 => x"01484305",
			4267 => x"fcf34305",
			4268 => x"06019128",
			4269 => x"0004bc18",
			4270 => x"00042e08",
			4271 => x"0f08d404",
			4272 => x"feb74305",
			4273 => x"01cc4305",
			4274 => x"0307b008",
			4275 => x"0e062e04",
			4276 => x"078c4305",
			4277 => x"02624305",
			4278 => x"0506f104",
			4279 => x"10274305",
			4280 => x"02fb4305",
			4281 => x"06016604",
			4282 => x"00204305",
			4283 => x"04100804",
			4284 => x"006d4305",
			4285 => x"0f08aa04",
			4286 => x"01d24305",
			4287 => x"02ad4305",
			4288 => x"fe654305",
			4289 => x"07050408",
			4290 => x"0209ef04",
			4291 => x"fea643a1",
			4292 => x"000043a1",
			4293 => x"0705060c",
			4294 => x"0208e408",
			4295 => x"0d05f704",
			4296 => x"000043a1",
			4297 => x"01cc43a1",
			4298 => x"000043a1",
			4299 => x"08036814",
			4300 => x"040baa04",
			4301 => x"fefe43a1",
			4302 => x"0100fa0c",
			4303 => x"01007e04",
			4304 => x"000043a1",
			4305 => x"0c04ee04",
			4306 => x"000043a1",
			4307 => x"00e143a1",
			4308 => x"000043a1",
			4309 => x"0f084f18",
			4310 => x"0e05520c",
			4311 => x"0209dd08",
			4312 => x"0c04f104",
			4313 => x"000043a1",
			4314 => x"ff9943a1",
			4315 => x"000043a1",
			4316 => x"040e2304",
			4317 => x"000043a1",
			4318 => x"0c04ed04",
			4319 => x"000043a1",
			4320 => x"009a43a1",
			4321 => x"0209f704",
			4322 => x"000043a1",
			4323 => x"0d073004",
			4324 => x"fec543a1",
			4325 => x"03087504",
			4326 => x"000043a1",
			4327 => x"ffec43a1",
			4328 => x"0d05f704",
			4329 => x"fe6a443d",
			4330 => x"0c05631c",
			4331 => x"00040204",
			4332 => x"feb2443d",
			4333 => x"00040708",
			4334 => x"08033404",
			4335 => x"052d443d",
			4336 => x"0000443d",
			4337 => x"040c6604",
			4338 => x"fea8443d",
			4339 => x"0505ce04",
			4340 => x"0391443d",
			4341 => x"040d4204",
			4342 => x"ff71443d",
			4343 => x"0115443d",
			4344 => x"0c059e1c",
			4345 => x"0d079614",
			4346 => x"0d07300c",
			4347 => x"07058e08",
			4348 => x"07058c04",
			4349 => x"ff6b443d",
			4350 => x"0000443d",
			4351 => x"fe96443d",
			4352 => x"0100e804",
			4353 => x"00ea443d",
			4354 => x"feca443d",
			4355 => x"040bd804",
			4356 => x"0000443d",
			4357 => x"01b5443d",
			4358 => x"020b1c04",
			4359 => x"fe68443d",
			4360 => x"0c05dc04",
			4361 => x"0136443d",
			4362 => x"020b1f08",
			4363 => x"0c063404",
			4364 => x"006e443d",
			4365 => x"0000443d",
			4366 => x"fe87443d",
			4367 => x"0d05f704",
			4368 => x"fe9444e1",
			4369 => x"0208dd18",
			4370 => x"05062310",
			4371 => x"0803660c",
			4372 => x"00040204",
			4373 => x"000044e1",
			4374 => x"0c050c04",
			4375 => x"01e144e1",
			4376 => x"000044e1",
			4377 => x"000044e1",
			4378 => x"0a02cb04",
			4379 => x"ffc544e1",
			4380 => x"000044e1",
			4381 => x"0100b418",
			4382 => x"0e06ac14",
			4383 => x"05063508",
			4384 => x"0e054b04",
			4385 => x"000044e1",
			4386 => x"ff0344e1",
			4387 => x"06016304",
			4388 => x"000044e1",
			4389 => x"00072404",
			4390 => x"00c344e1",
			4391 => x"000044e1",
			4392 => x"fe9344e1",
			4393 => x"0100e710",
			4394 => x"020b2c0c",
			4395 => x"06016f04",
			4396 => x"000044e1",
			4397 => x"0100bb04",
			4398 => x"000044e1",
			4399 => x"00e944e1",
			4400 => x"ffd344e1",
			4401 => x"020b5304",
			4402 => x"ff3644e1",
			4403 => x"0a029b08",
			4404 => x"0901bc04",
			4405 => x"005d44e1",
			4406 => x"000044e1",
			4407 => x"000044e1",
			4408 => x"02099528",
			4409 => x"01006f04",
			4410 => x"fe6145b5",
			4411 => x"0a02dd1c",
			4412 => x"0f077b18",
			4413 => x"0a02a810",
			4414 => x"0f077908",
			4415 => x"0a028304",
			4416 => x"fe6a45b5",
			4417 => x"ff3745b5",
			4418 => x"0a027804",
			4419 => x"ff8c45b5",
			4420 => x"05e245b5",
			4421 => x"0305e904",
			4422 => x"fea645b5",
			4423 => x"0cc845b5",
			4424 => x"fe6d45b5",
			4425 => x"0b055604",
			4426 => x"fee345b5",
			4427 => x"01d245b5",
			4428 => x"0c059e34",
			4429 => x"06018928",
			4430 => x"0d070814",
			4431 => x"0900bc08",
			4432 => x"02099d04",
			4433 => x"002645b5",
			4434 => x"fe5345b5",
			4435 => x"0a02b004",
			4436 => x"fea445b5",
			4437 => x"06016604",
			4438 => x"ffb845b5",
			4439 => x"020045b5",
			4440 => x"09019010",
			4441 => x"0e073b08",
			4442 => x"09015c04",
			4443 => x"032f45b5",
			4444 => x"ff2545b5",
			4445 => x"08033904",
			4446 => x"03ef45b5",
			4447 => x"077a45b5",
			4448 => x"fe9f45b5",
			4449 => x"05079008",
			4450 => x"0803dc04",
			4451 => x"fe6445b5",
			4452 => x"fc9345b5",
			4453 => x"01b445b5",
			4454 => x"0e0a2a0c",
			4455 => x"020b1c04",
			4456 => x"fe6645b5",
			4457 => x"08037f04",
			4458 => x"054345b5",
			4459 => x"ff0745b5",
			4460 => x"fe6245b5",
			4461 => x"0d05f704",
			4462 => x"fe744669",
			4463 => x"0c050c1c",
			4464 => x"0e05960c",
			4465 => x"040c2404",
			4466 => x"00004669",
			4467 => x"06017c04",
			4468 => x"01a64669",
			4469 => x"00004669",
			4470 => x"0c050a08",
			4471 => x"04100804",
			4472 => x"feaa4669",
			4473 => x"00144669",
			4474 => x"09010604",
			4475 => x"00004669",
			4476 => x"01c74669",
			4477 => x"06016b0c",
			4478 => x"0c052508",
			4479 => x"0e05b304",
			4480 => x"000b4669",
			4481 => x"00004669",
			4482 => x"fdf44669",
			4483 => x"0601811c",
			4484 => x"040d880c",
			4485 => x"0d075504",
			4486 => x"ff0a4669",
			4487 => x"0100f504",
			4488 => x"00f14669",
			4489 => x"ff6b4669",
			4490 => x"0100de08",
			4491 => x"0900cb04",
			4492 => x"00004669",
			4493 => x"01584669",
			4494 => x"0209d404",
			4495 => x"005d4669",
			4496 => x"ff624669",
			4497 => x"020b0808",
			4498 => x"03079c04",
			4499 => x"00004669",
			4500 => x"fe804669",
			4501 => x"030a6908",
			4502 => x"0a02d404",
			4503 => x"01164669",
			4504 => x"00004669",
			4505 => x"fef94669",
			4506 => x"0d05f704",
			4507 => x"fe6f4715",
			4508 => x"0c05282c",
			4509 => x"0c050718",
			4510 => x"0e059610",
			4511 => x"040d2e04",
			4512 => x"fffa4715",
			4513 => x"06017808",
			4514 => x"0d066b04",
			4515 => x"01ce4715",
			4516 => x"00004715",
			4517 => x"00004715",
			4518 => x"04100804",
			4519 => x"fe964715",
			4520 => x"00004715",
			4521 => x"0f08d410",
			4522 => x"08032804",
			4523 => x"00004715",
			4524 => x"01007c04",
			4525 => x"00004715",
			4526 => x"0a029304",
			4527 => x"02914715",
			4528 => x"01404715",
			4529 => x"00004715",
			4530 => x"06016308",
			4531 => x"0c052e04",
			4532 => x"00004715",
			4533 => x"fe434715",
			4534 => x"0100fa1c",
			4535 => x"0a02a10c",
			4536 => x"0d071604",
			4537 => x"ff6b4715",
			4538 => x"0a028d04",
			4539 => x"ffed4715",
			4540 => x"01444715",
			4541 => x"0f094508",
			4542 => x"0a02d704",
			4543 => x"ff884715",
			4544 => x"01024715",
			4545 => x"09017404",
			4546 => x"fe884715",
			4547 => x"00004715",
			4548 => x"fe904715",
			4549 => x"0d05f704",
			4550 => x"fea247a1",
			4551 => x"02083d0c",
			4552 => x"0b054508",
			4553 => x"0409db04",
			4554 => x"000047a1",
			4555 => x"019f47a1",
			4556 => x"000047a1",
			4557 => x"040c7f04",
			4558 => x"febf47a1",
			4559 => x"0a02c31c",
			4560 => x"0c05630c",
			4561 => x"0c04ef04",
			4562 => x"000047a1",
			4563 => x"0a028d04",
			4564 => x"000047a1",
			4565 => x"012247a1",
			4566 => x"0f093d08",
			4567 => x"0f08aa04",
			4568 => x"000047a1",
			4569 => x"ff8c47a1",
			4570 => x"0100fc04",
			4571 => x"00e447a1",
			4572 => x"000047a1",
			4573 => x"06018810",
			4574 => x"06017308",
			4575 => x"0c052804",
			4576 => x"003b47a1",
			4577 => x"ff5947a1",
			4578 => x"040eab04",
			4579 => x"000047a1",
			4580 => x"00ba47a1",
			4581 => x"0100dc04",
			4582 => x"feac47a1",
			4583 => x"000047a1",
			4584 => x"0b053504",
			4585 => x"fe77482d",
			4586 => x"040baa04",
			4587 => x"fe9a482d",
			4588 => x"08036818",
			4589 => x"0100fa14",
			4590 => x"0c050b04",
			4591 => x"01dd482d",
			4592 => x"0c056208",
			4593 => x"0d071604",
			4594 => x"ff5d482d",
			4595 => x"0000482d",
			4596 => x"0d071604",
			4597 => x"0000482d",
			4598 => x"013c482d",
			4599 => x"ff5a482d",
			4600 => x"06016a14",
			4601 => x"0c052e0c",
			4602 => x"040e2304",
			4603 => x"ff7a482d",
			4604 => x"01007304",
			4605 => x"0000482d",
			4606 => x"0100482d",
			4607 => x"0e05f704",
			4608 => x"fdf2482d",
			4609 => x"0000482d",
			4610 => x"0601810c",
			4611 => x"040e6304",
			4612 => x"ff34482d",
			4613 => x"0100d204",
			4614 => x"016d482d",
			4615 => x"0000482d",
			4616 => x"0f08b104",
			4617 => x"0000482d",
			4618 => x"fede482d",
			4619 => x"01007e04",
			4620 => x"fe7e48db",
			4621 => x"0a02c324",
			4622 => x"0003e104",
			4623 => x"fec048db",
			4624 => x"0c04ee04",
			4625 => x"ff2148db",
			4626 => x"0a02920c",
			4627 => x"0100f308",
			4628 => x"0a027f04",
			4629 => x"000048db",
			4630 => x"01ba48db",
			4631 => x"000048db",
			4632 => x"040dca08",
			4633 => x"0c057f04",
			4634 => x"ff2848db",
			4635 => x"000048db",
			4636 => x"0e071504",
			4637 => x"000048db",
			4638 => x"019248db",
			4639 => x"00055428",
			4640 => x"0c05601c",
			4641 => x"0c052810",
			4642 => x"05063208",
			4643 => x"06016b04",
			4644 => x"000048db",
			4645 => x"ffbb48db",
			4646 => x"06018d04",
			4647 => x"005048db",
			4648 => x"000048db",
			4649 => x"0209d404",
			4650 => x"000048db",
			4651 => x"020a6304",
			4652 => x"fdf648db",
			4653 => x"000048db",
			4654 => x"0c059e08",
			4655 => x"09012004",
			4656 => x"000048db",
			4657 => x"00c648db",
			4658 => x"ffa948db",
			4659 => x"020b2c04",
			4660 => x"010248db",
			4661 => x"000048db",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1522, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(3074, initial_addr_3'length));
	end generate gen_rom_13;

	gen_rom_14: if SELECT_ROM = 14 generate
		bank <= (
			0 => x"07057358",
			1 => x"040f7054",
			2 => x"06010714",
			3 => x"03043508",
			4 => x"0f061a04",
			5 => x"025f00d5",
			6 => x"ff5500d5",
			7 => x"03047f08",
			8 => x"0e039704",
			9 => x"feaf00d5",
			10 => x"007400d5",
			11 => x"fe6200d5",
			12 => x"0704be20",
			13 => x"03051b10",
			14 => x"07047808",
			15 => x"0208c004",
			16 => x"01fb00d5",
			17 => x"fe6100d5",
			18 => x"0a024704",
			19 => x"029200d5",
			20 => x"006400d5",
			21 => x"02082a08",
			22 => x"040bb204",
			23 => x"018400d5",
			24 => x"031d00d5",
			25 => x"0a028504",
			26 => x"003600d5",
			27 => x"012b00d5",
			28 => x"0e057110",
			29 => x"0208bb08",
			30 => x"06012b04",
			31 => x"fef700d5",
			32 => x"007700d5",
			33 => x"0704ef04",
			34 => x"ff1a00d5",
			35 => x"013f00d5",
			36 => x"0704ee08",
			37 => x"0e06ac04",
			38 => x"013700d5",
			39 => x"fe8500d5",
			40 => x"06017d04",
			41 => x"008400d5",
			42 => x"fefc00d5",
			43 => x"fe5e00d5",
			44 => x"0a024510",
			45 => x"0f0a420c",
			46 => x"07058d08",
			47 => x"0801e404",
			48 => x"febd00d5",
			49 => x"015a00d5",
			50 => x"fe5f00d5",
			51 => x"039700d5",
			52 => x"fe5e00d5",
			53 => x"0004b888",
			54 => x"0504e71c",
			55 => x"00047d0c",
			56 => x"09005d08",
			57 => x"0504c804",
			58 => x"00000259",
			59 => x"ffb80259",
			60 => x"020b0259",
			61 => x"040c9304",
			62 => x"feb70259",
			63 => x"0b045c04",
			64 => x"00000259",
			65 => x"0a029304",
			66 => x"00000259",
			67 => x"01c20259",
			68 => x"01004b30",
			69 => x"09007d20",
			70 => x"02082f10",
			71 => x"06013508",
			72 => x"0f06e504",
			73 => x"ffb70259",
			74 => x"030f0259",
			75 => x"01004904",
			76 => x"00340259",
			77 => x"022e0259",
			78 => x"02084b08",
			79 => x"00043f04",
			80 => x"01f30259",
			81 => x"fe6b0259",
			82 => x"01004704",
			83 => x"00840259",
			84 => x"ff520259",
			85 => x"05051408",
			86 => x"0e047104",
			87 => x"fe520259",
			88 => x"00e20259",
			89 => x"0a02b004",
			90 => x"fdcd0259",
			91 => x"ffb20259",
			92 => x"0d054d1c",
			93 => x"0305330c",
			94 => x"0b04c308",
			95 => x"0b04b104",
			96 => x"fffb0259",
			97 => x"00d30259",
			98 => x"fd760259",
			99 => x"0208ab08",
			100 => x"00043e04",
			101 => x"007d0259",
			102 => x"01a60259",
			103 => x"09009104",
			104 => x"00d00259",
			105 => x"fe220259",
			106 => x"01005c10",
			107 => x"0b04d208",
			108 => x"0d057504",
			109 => x"ffae0259",
			110 => x"fe200259",
			111 => x"01005804",
			112 => x"01df0259",
			113 => x"ffdb0259",
			114 => x"09009c08",
			115 => x"03057704",
			116 => x"003e0259",
			117 => x"01770259",
			118 => x"01006204",
			119 => x"ff840259",
			120 => x"00020259",
			121 => x"0208c224",
			122 => x"0e04b420",
			123 => x"0304d614",
			124 => x"0f06f310",
			125 => x"0a02d108",
			126 => x"0e041604",
			127 => x"fe750259",
			128 => x"00630259",
			129 => x"0004e904",
			130 => x"00990259",
			131 => x"ff6c0259",
			132 => x"02c80259",
			133 => x"0a02e404",
			134 => x"fe850259",
			135 => x"0f06e504",
			136 => x"00f10259",
			137 => x"ff620259",
			138 => x"01310259",
			139 => x"01007110",
			140 => x"0803be04",
			141 => x"fe510259",
			142 => x"01005608",
			143 => x"0f071704",
			144 => x"ffe20259",
			145 => x"01840259",
			146 => x"febc0259",
			147 => x"0b052404",
			148 => x"011d0259",
			149 => x"feeb0259",
			150 => x"09007b50",
			151 => x"0c04912c",
			152 => x"0c048f28",
			153 => x"0208c220",
			154 => x"040d6e10",
			155 => x"0e03e708",
			156 => x"0b049104",
			157 => x"ffe703bd",
			158 => x"fe6803bd",
			159 => x"0c045704",
			160 => x"ff9103bd",
			161 => x"007603bd",
			162 => x"0a02ed08",
			163 => x"0d04f304",
			164 => x"034703bd",
			165 => x"00fb03bd",
			166 => x"0b047d04",
			167 => x"ff5603bd",
			168 => x"012c03bd",
			169 => x"040c7204",
			170 => x"006003bd",
			171 => x"fdf103bd",
			172 => x"fe5703bd",
			173 => x"0100430c",
			174 => x"0e044408",
			175 => x"01003904",
			176 => x"000003bd",
			177 => x"fe5f03bd",
			178 => x"004d03bd",
			179 => x"0c04b014",
			180 => x"0e046810",
			181 => x"0d052608",
			182 => x"09007504",
			183 => x"01dc03bd",
			184 => x"005c03bd",
			185 => x"0b04a004",
			186 => x"ff0d03bd",
			187 => x"00c303bd",
			188 => x"02b703bd",
			189 => x"fe6b03bd",
			190 => x"01005130",
			191 => x"0c045504",
			192 => x"019203bd",
			193 => x"02087614",
			194 => x"040cf510",
			195 => x"0e048808",
			196 => x"07047804",
			197 => x"016103bd",
			198 => x"ff8503bd",
			199 => x"01004f04",
			200 => x"ffd603bd",
			201 => x"014703bd",
			202 => x"01bf03bd",
			203 => x"0900800c",
			204 => x"09007f08",
			205 => x"0f072b04",
			206 => x"fe0603bd",
			207 => x"ffe803bd",
			208 => x"009103bd",
			209 => x"06014604",
			210 => x"fe0803bd",
			211 => x"0004a304",
			212 => x"000f03bd",
			213 => x"fe3203bd",
			214 => x"07047a04",
			215 => x"017303bd",
			216 => x"0c045b14",
			217 => x"0d05410c",
			218 => x"01005508",
			219 => x"0e048804",
			220 => x"fe7103bd",
			221 => x"002f03bd",
			222 => x"016e03bd",
			223 => x"040c1e04",
			224 => x"fe3003bd",
			225 => x"ffc003bd",
			226 => x"0c04720c",
			227 => x"02081d04",
			228 => x"ff6c03bd",
			229 => x"07049504",
			230 => x"02ae03bd",
			231 => x"009603bd",
			232 => x"0d052608",
			233 => x"040c3204",
			234 => x"fe1203bd",
			235 => x"004503bd",
			236 => x"0c04ec04",
			237 => x"001103bd",
			238 => x"ffbb03bd",
			239 => x"0c04d194",
			240 => x"07050464",
			241 => x"0704f13c",
			242 => x"0c04ca20",
			243 => x"02086210",
			244 => x"02086008",
			245 => x"01007504",
			246 => x"000a0571",
			247 => x"00d80571",
			248 => x"0a02a804",
			249 => x"016b0571",
			250 => x"ff8b0571",
			251 => x"0a02b108",
			252 => x"0e052004",
			253 => x"ff970571",
			254 => x"fff80571",
			255 => x"0c049104",
			256 => x"ff8e0571",
			257 => x"006e0571",
			258 => x"0a02bb10",
			259 => x"0b04d008",
			260 => x"02083104",
			261 => x"ffeb0571",
			262 => x"01890571",
			263 => x"0f07c004",
			264 => x"fef80571",
			265 => x"fffa0571",
			266 => x"0a02be04",
			267 => x"01f40571",
			268 => x"06016304",
			269 => x"ff0c0571",
			270 => x"012d0571",
			271 => x"00047520",
			272 => x"08034210",
			273 => x"0f07eb08",
			274 => x"0c04b404",
			275 => x"ff900571",
			276 => x"01410571",
			277 => x"0a029504",
			278 => x"fe360571",
			279 => x"01150571",
			280 => x"0a02b008",
			281 => x"0d05dc04",
			282 => x"02490571",
			283 => x"014e0571",
			284 => x"03065904",
			285 => x"ff8e0571",
			286 => x"01c20571",
			287 => x"0d05cf04",
			288 => x"fdeb0571",
			289 => x"008c0571",
			290 => x"0209131c",
			291 => x"01008c10",
			292 => x"02084b04",
			293 => x"00fd0571",
			294 => x"07051804",
			295 => x"fde60571",
			296 => x"0e05e904",
			297 => x"ffef0571",
			298 => x"fdf10571",
			299 => x"0d062a04",
			300 => x"01810571",
			301 => x"07051a04",
			302 => x"fe2c0571",
			303 => x"00620571",
			304 => x"00043a08",
			305 => x"0b056904",
			306 => x"fdfe0571",
			307 => x"00140571",
			308 => x"06016b04",
			309 => x"01ed0571",
			310 => x"07051804",
			311 => x"fe6c0571",
			312 => x"00d40571",
			313 => x"0c04d218",
			314 => x"02089308",
			315 => x"02082404",
			316 => x"00000571",
			317 => x"02290571",
			318 => x"0208b204",
			319 => x"ff490571",
			320 => x"0d05b504",
			321 => x"ffc40571",
			322 => x"01008604",
			323 => x"02010571",
			324 => x"00000571",
			325 => x"00049628",
			326 => x"08038a20",
			327 => x"0c04ea10",
			328 => x"0c04e908",
			329 => x"0e05d804",
			330 => x"ffb70571",
			331 => x"01610571",
			332 => x"06015204",
			333 => x"ffda0571",
			334 => x"fe210571",
			335 => x"01006b08",
			336 => x"06015204",
			337 => x"00000571",
			338 => x"fdf30571",
			339 => x"06015404",
			340 => x"00ea0571",
			341 => x"00050571",
			342 => x"02098e04",
			343 => x"032e0571",
			344 => x"00000571",
			345 => x"0b050204",
			346 => x"000d0571",
			347 => x"fe600571",
			348 => x"07053278",
			349 => x"01002d08",
			350 => x"06014604",
			351 => x"fe5606d5",
			352 => x"00ed06d5",
			353 => x"040c263c",
			354 => x"06013a20",
			355 => x"02084d10",
			356 => x"00044b08",
			357 => x"06013504",
			358 => x"00b606d5",
			359 => x"019f06d5",
			360 => x"040bf104",
			361 => x"fe8506d5",
			362 => x"007f06d5",
			363 => x"0003ed08",
			364 => x"040abb04",
			365 => x"000006d5",
			366 => x"fe0706d5",
			367 => x"03057904",
			368 => x"ffb506d5",
			369 => x"013806d5",
			370 => x"0c04cb0c",
			371 => x"01009508",
			372 => x"040b9704",
			373 => x"020106d5",
			374 => x"016706d5",
			375 => x"fe1a06d5",
			376 => x"0c04cc08",
			377 => x"040ba404",
			378 => x"fd3e06d5",
			379 => x"fe7506d5",
			380 => x"06017904",
			381 => x"00e906d5",
			382 => x"fe8406d5",
			383 => x"0c049314",
			384 => x"0a028304",
			385 => x"fe5b06d5",
			386 => x"09007b08",
			387 => x"0304b704",
			388 => x"00e206d5",
			389 => x"030506d5",
			390 => x"03050004",
			391 => x"ffd406d5",
			392 => x"012406d5",
			393 => x"06014a10",
			394 => x"02086f08",
			395 => x"07049104",
			396 => x"fe9306d5",
			397 => x"006906d5",
			398 => x"0900a004",
			399 => x"ff5d06d5",
			400 => x"fded06d5",
			401 => x"040cbf08",
			402 => x"09009804",
			403 => x"01be06d5",
			404 => x"007906d5",
			405 => x"0c049704",
			406 => x"00a306d5",
			407 => x"ff2a06d5",
			408 => x"0c054524",
			409 => x"0d069f10",
			410 => x"0e062e04",
			411 => x"fe5206d5",
			412 => x"0e06ac08",
			413 => x"0003d104",
			414 => x"fea106d5",
			415 => x"01da06d5",
			416 => x"fe3f06d5",
			417 => x"040c0c10",
			418 => x"00032c04",
			419 => x"fe7306d5",
			420 => x"06017c04",
			421 => x"039006d5",
			422 => x"0a02b804",
			423 => x"fe7406d5",
			424 => x"005206d5",
			425 => x"fe6206d5",
			426 => x"0c05b814",
			427 => x"07063d10",
			428 => x"0705730c",
			429 => x"07056104",
			430 => x"fe8206d5",
			431 => x"0c054c04",
			432 => x"00cc06d5",
			433 => x"ff0406d5",
			434 => x"fe5e06d5",
			435 => x"049f06d5",
			436 => x"fe5506d5",
			437 => x"0e061e90",
			438 => x"0900cd5c",
			439 => x"01007930",
			440 => x"0900c220",
			441 => x"06014f10",
			442 => x"0208bb08",
			443 => x"0c04b404",
			444 => x"fff908a9",
			445 => x"006a08a9",
			446 => x"0900b304",
			447 => x"ffb008a9",
			448 => x"fe6308a9",
			449 => x"0c04d008",
			450 => x"03053704",
			451 => x"ffad08a9",
			452 => x"007408a9",
			453 => x"0305f204",
			454 => x"ff1d08a9",
			455 => x"00f808a9",
			456 => x"040c850c",
			457 => x"0505cc08",
			458 => x"00046704",
			459 => x"ffcf08a9",
			460 => x"fdf808a9",
			461 => x"fd8c08a9",
			462 => x"013408a9",
			463 => x"040b5d14",
			464 => x"06012d08",
			465 => x"0900c404",
			466 => x"000008a9",
			467 => x"048208a9",
			468 => x"0305e908",
			469 => x"0704ec04",
			470 => x"01ad08a9",
			471 => x"000008a9",
			472 => x"01d308a9",
			473 => x"0306190c",
			474 => x"0900c204",
			475 => x"01be08a9",
			476 => x"00044a04",
			477 => x"ffae08a9",
			478 => x"fe2008a9",
			479 => x"040c5e08",
			480 => x"01007c04",
			481 => x"02b208a9",
			482 => x"00da08a9",
			483 => x"ffc208a9",
			484 => x"00044f1c",
			485 => x"01007d04",
			486 => x"fe5a08a9",
			487 => x"040b910c",
			488 => x"01008e08",
			489 => x"03062104",
			490 => x"ff1308a9",
			491 => x"008308a9",
			492 => x"fdcf08a9",
			493 => x"040baa04",
			494 => x"01ff08a9",
			495 => x"0208d604",
			496 => x"fec908a9",
			497 => x"011e08a9",
			498 => x"0900ec10",
			499 => x"06017404",
			500 => x"fe4e08a9",
			501 => x"0505f604",
			502 => x"fef708a9",
			503 => x"01008604",
			504 => x"016608a9",
			505 => x"000008a9",
			506 => x"0b058504",
			507 => x"015c08a9",
			508 => x"000008a9",
			509 => x"06017944",
			510 => x"0c04e924",
			511 => x"0c04af08",
			512 => x"040b6904",
			513 => x"01b308a9",
			514 => x"fd9308a9",
			515 => x"08035010",
			516 => x"08032808",
			517 => x"02086e04",
			518 => x"000008a9",
			519 => x"018408a9",
			520 => x"08033704",
			521 => x"fef908a9",
			522 => x"008a08a9",
			523 => x"0c04d008",
			524 => x"0c04b904",
			525 => x"010508a9",
			526 => x"028a08a9",
			527 => x"00c408a9",
			528 => x"0c04ea04",
			529 => x"fdc208a9",
			530 => x"0306830c",
			531 => x"07052f04",
			532 => x"fe9d08a9",
			533 => x"05065f04",
			534 => x"015608a9",
			535 => x"000008a9",
			536 => x"0306a508",
			537 => x"0c050b04",
			538 => x"01e008a9",
			539 => x"ff0f08a9",
			540 => x"0d065f04",
			541 => x"ff9708a9",
			542 => x"00b408a9",
			543 => x"0d061f08",
			544 => x"0e067104",
			545 => x"ff7308a9",
			546 => x"013308a9",
			547 => x"06018c04",
			548 => x"fe5e08a9",
			549 => x"02096c08",
			550 => x"05064204",
			551 => x"000008a9",
			552 => x"018908a9",
			553 => x"feb408a9",
			554 => x"0c054388",
			555 => x"0100320c",
			556 => x"06014604",
			557 => x"fe5a09e5",
			558 => x"07048004",
			559 => x"01a409e5",
			560 => x"fee609e5",
			561 => x"09008240",
			562 => x"0304d820",
			563 => x"09007e10",
			564 => x"03049708",
			565 => x"0c045504",
			566 => x"01aa09e5",
			567 => x"ffe809e5",
			568 => x"0f064a04",
			569 => x"04a209e5",
			570 => x"00a409e5",
			571 => x"01004f08",
			572 => x"0c047304",
			573 => x"ff8909e5",
			574 => x"fe2009e5",
			575 => x"0f069604",
			576 => x"01da09e5",
			577 => x"fefe09e5",
			578 => x"0f06d010",
			579 => x"0e045308",
			580 => x"0a029204",
			581 => x"ff4b09e5",
			582 => x"02fb09e5",
			583 => x"0003e604",
			584 => x"ff3d09e5",
			585 => x"038d09e5",
			586 => x"08032908",
			587 => x"0e049604",
			588 => x"fe2309e5",
			589 => x"007e09e5",
			590 => x"0304fe04",
			591 => x"002809e5",
			592 => x"019c09e5",
			593 => x"0e04e21c",
			594 => x"03055f10",
			595 => x"03055308",
			596 => x"03054f04",
			597 => x"002109e5",
			598 => x"fe3109e5",
			599 => x"02086f04",
			600 => x"01cc09e5",
			601 => x"ffb209e5",
			602 => x"08039908",
			603 => x"0f06d604",
			604 => x"009209e5",
			605 => x"fee009e5",
			606 => x"04e909e5",
			607 => x"0900af10",
			608 => x"0208d008",
			609 => x"0704c404",
			610 => x"00ad09e5",
			611 => x"015809e5",
			612 => x"06014f04",
			613 => x"ff1809e5",
			614 => x"008b09e5",
			615 => x"0e057808",
			616 => x"0d057404",
			617 => x"021c09e5",
			618 => x"ffbe09e5",
			619 => x"0900cf04",
			620 => x"00be09e5",
			621 => x"fff909e5",
			622 => x"0c05b814",
			623 => x"0d083010",
			624 => x"0705730c",
			625 => x"07056104",
			626 => x"feb409e5",
			627 => x"0c054c04",
			628 => x"006109e5",
			629 => x"000009e5",
			630 => x"fe6b09e5",
			631 => x"030709e5",
			632 => x"fe6509e5",
			633 => x"0705326c",
			634 => x"01002a04",
			635 => x"fe5a0b41",
			636 => x"040c2638",
			637 => x"07050420",
			638 => x"06013e10",
			639 => x"02086c08",
			640 => x"0e04e204",
			641 => x"009a0b41",
			642 => x"015f0b41",
			643 => x"00040b04",
			644 => x"feb30b41",
			645 => x"00400b41",
			646 => x"0704be08",
			647 => x"0f072d04",
			648 => x"02620b41",
			649 => x"018b0b41",
			650 => x"0e054b04",
			651 => x"00a70b41",
			652 => x"01820b41",
			653 => x"0803610c",
			654 => x"06017308",
			655 => x"0f074f04",
			656 => x"feb90b41",
			657 => x"01130b41",
			658 => x"fe5a0b41",
			659 => x"040c0c08",
			660 => x"02095104",
			661 => x"fdf20b41",
			662 => x"00000b41",
			663 => x"fff70b41",
			664 => x"09008f14",
			665 => x"06012304",
			666 => x"fe5f0b41",
			667 => x"0e049d08",
			668 => x"07047d04",
			669 => x"018a0b41",
			670 => x"006e0b41",
			671 => x"0208a604",
			672 => x"02ba0b41",
			673 => x"01080b41",
			674 => x"0305370c",
			675 => x"0d054104",
			676 => x"01f60b41",
			677 => x"02081d04",
			678 => x"001d0b41",
			679 => x"feab0b41",
			680 => x"06014a08",
			681 => x"0e050004",
			682 => x"00030b41",
			683 => x"fe5b0b41",
			684 => x"040c9304",
			685 => x"00d40b41",
			686 => x"ffe60b41",
			687 => x"07058b24",
			688 => x"0e062e04",
			689 => x"fe570b41",
			690 => x"02098e1c",
			691 => x"0d069f0c",
			692 => x"0e06ac08",
			693 => x"0003d104",
			694 => x"fe9c0b41",
			695 => x"01380b41",
			696 => x"fe480b41",
			697 => x"06014508",
			698 => x"0b05d804",
			699 => x"fe660b41",
			700 => x"00000b41",
			701 => x"0b05bf04",
			702 => x"03fd0b41",
			703 => x"00dd0b41",
			704 => x"fe670b41",
			705 => x"0802cc1c",
			706 => x"040abb10",
			707 => x"0705a40c",
			708 => x"0705a208",
			709 => x"07058d04",
			710 => x"00000b41",
			711 => x"ffca0b41",
			712 => x"00dc0b41",
			713 => x"fe5a0b41",
			714 => x"00036804",
			715 => x"04dc0b41",
			716 => x"040af704",
			717 => x"fe830b41",
			718 => x"01d10b41",
			719 => x"fe580b41",
			720 => x"09007b68",
			721 => x"0c049138",
			722 => x"0c048f34",
			723 => x"040d6e1c",
			724 => x"0e03e70c",
			725 => x"0b049108",
			726 => x"02079b04",
			727 => x"00c90cdd",
			728 => x"ff810cdd",
			729 => x"fe5d0cdd",
			730 => x"0f06b208",
			731 => x"08036504",
			732 => x"00570cdd",
			733 => x"01780cdd",
			734 => x"0c047a04",
			735 => x"ffe40cdd",
			736 => x"02400cdd",
			737 => x"0a02ed0c",
			738 => x"0207c504",
			739 => x"05db0cdd",
			740 => x"040dca04",
			741 => x"01e00cdd",
			742 => x"ffff0cdd",
			743 => x"0a02f704",
			744 => x"fe600cdd",
			745 => x"040fc604",
			746 => x"00f40cdd",
			747 => x"ff710cdd",
			748 => x"fe480cdd",
			749 => x"01004308",
			750 => x"0e044404",
			751 => x"fe6b0cdd",
			752 => x"00720cdd",
			753 => x"02080714",
			754 => x"0207d70c",
			755 => x"07049708",
			756 => x"06012804",
			757 => x"010c0cdd",
			758 => x"fe870cdd",
			759 => x"02740cdd",
			760 => x"040c2c04",
			761 => x"fe320cdd",
			762 => x"00660cdd",
			763 => x"0c04950c",
			764 => x"0d051a04",
			765 => x"031d0cdd",
			766 => x"0e043604",
			767 => x"ffa60cdd",
			768 => x"02b60cdd",
			769 => x"0a02b804",
			770 => x"01840cdd",
			771 => x"ff2e0cdd",
			772 => x"01005128",
			773 => x"0c045504",
			774 => x"01b30cdd",
			775 => x"02087614",
			776 => x"040cf510",
			777 => x"0e048808",
			778 => x"0b049104",
			779 => x"000b0cdd",
			780 => x"ff430cdd",
			781 => x"06013104",
			782 => x"01810cdd",
			783 => x"ffeb0cdd",
			784 => x"01ef0cdd",
			785 => x"0900860c",
			786 => x"0a029604",
			787 => x"fdda0cdd",
			788 => x"00049604",
			789 => x"00340cdd",
			790 => x"feaf0cdd",
			791 => x"fdec0cdd",
			792 => x"07047a04",
			793 => x"01990cdd",
			794 => x"0c04ec20",
			795 => x"0a027a10",
			796 => x"0a027708",
			797 => x"0e04e204",
			798 => x"ffb30cdd",
			799 => x"00360cdd",
			800 => x"040af504",
			801 => x"fd8d0cdd",
			802 => x"ff820cdd",
			803 => x"08032e08",
			804 => x"0f079604",
			805 => x"01180cdd",
			806 => x"ffd90cdd",
			807 => x"0a028504",
			808 => x"ffb90cdd",
			809 => x"001e0cdd",
			810 => x"040c3210",
			811 => x"040b6308",
			812 => x"08032e04",
			813 => x"ffd00cdd",
			814 => x"fdd70cdd",
			815 => x"00047104",
			816 => x"00880cdd",
			817 => x"fe920cdd",
			818 => x"08037a04",
			819 => x"fe190cdd",
			820 => x"00048604",
			821 => x"00d40cdd",
			822 => x"fea40cdd",
			823 => x"0207a164",
			824 => x"02076728",
			825 => x"0003c418",
			826 => x"0305170c",
			827 => x"01004504",
			828 => x"ff8d0ed9",
			829 => x"0e043604",
			830 => x"00b10ed9",
			831 => x"022c0ed9",
			832 => x"0f067404",
			833 => x"fe830ed9",
			834 => x"04089204",
			835 => x"00000ed9",
			836 => x"00850ed9",
			837 => x"0c045c0c",
			838 => x"07047908",
			839 => x"07046604",
			840 => x"ffe10ed9",
			841 => x"013a0ed9",
			842 => x"fef40ed9",
			843 => x"fe4b0ed9",
			844 => x"0a026718",
			845 => x"040b0f10",
			846 => x"0304df04",
			847 => x"fea30ed9",
			848 => x"0003cc08",
			849 => x"02079204",
			850 => x"ffcf0ed9",
			851 => x"01a70ed9",
			852 => x"01de0ed9",
			853 => x"01004e04",
			854 => x"004a0ed9",
			855 => x"03a20ed9",
			856 => x"0a027508",
			857 => x"040b7004",
			858 => x"fdd90ed9",
			859 => x"00000ed9",
			860 => x"06012d0c",
			861 => x"0c045b08",
			862 => x"0c045a04",
			863 => x"fffd0ed9",
			864 => x"019e0ed9",
			865 => x"fe640ed9",
			866 => x"0c045a08",
			867 => x"01002d04",
			868 => x"00070ed9",
			869 => x"fe7c0ed9",
			870 => x"07047a04",
			871 => x"03410ed9",
			872 => x"01070ed9",
			873 => x"0e03e758",
			874 => x"0f064a24",
			875 => x"03047718",
			876 => x"01003f10",
			877 => x"03041608",
			878 => x"0d04d904",
			879 => x"00000ed9",
			880 => x"fe990ed9",
			881 => x"0a02d104",
			882 => x"ffcb0ed9",
			883 => x"02a00ed9",
			884 => x"040c0a04",
			885 => x"00000ed9",
			886 => x"fe6c0ed9",
			887 => x"03047f04",
			888 => x"021d0ed9",
			889 => x"06014d04",
			890 => x"001d0ed9",
			891 => x"00000ed9",
			892 => x"0e03bd20",
			893 => x"0f066d10",
			894 => x"06012d08",
			895 => x"0a02a004",
			896 => x"00000ed9",
			897 => x"011e0ed9",
			898 => x"0e037004",
			899 => x"006b0ed9",
			900 => x"fe590ed9",
			901 => x"0004a308",
			902 => x"00046804",
			903 => x"00000ed9",
			904 => x"025c0ed9",
			905 => x"0704a604",
			906 => x"ff690ed9",
			907 => x"00f70ed9",
			908 => x"01004b0c",
			909 => x"09006208",
			910 => x"0f068704",
			911 => x"01070ed9",
			912 => x"fe680ed9",
			913 => x"fe230ed9",
			914 => x"040c9a04",
			915 => x"00760ed9",
			916 => x"ff6a0ed9",
			917 => x"0f064a04",
			918 => x"01cf0ed9",
			919 => x"0a027020",
			920 => x"0a026a10",
			921 => x"06014908",
			922 => x"00040804",
			923 => x"ffbc0ed9",
			924 => x"00a50ed9",
			925 => x"0c04ec04",
			926 => x"01de0ed9",
			927 => x"00000ed9",
			928 => x"06013808",
			929 => x"08031704",
			930 => x"01480ed9",
			931 => x"ff480ed9",
			932 => x"0d059b04",
			933 => x"fe190ed9",
			934 => x"ffc50ed9",
			935 => x"0c049010",
			936 => x"01005e08",
			937 => x"0704a704",
			938 => x"002a0ed9",
			939 => x"ffa70ed9",
			940 => x"08034404",
			941 => x"001d0ed9",
			942 => x"011b0ed9",
			943 => x"0c049208",
			944 => x"01005a04",
			945 => x"ffee0ed9",
			946 => x"ff0d0ed9",
			947 => x"0c049304",
			948 => x"00c80ed9",
			949 => x"fffa0ed9",
			950 => x"07057380",
			951 => x"040fc67c",
			952 => x"0704913c",
			953 => x"0304af20",
			954 => x"09006210",
			955 => x"03043708",
			956 => x"0207d104",
			957 => x"ff560ffd",
			958 => x"01da0ffd",
			959 => x"06011c04",
			960 => x"fe970ffd",
			961 => x"02e30ffd",
			962 => x"02078b08",
			963 => x"03046704",
			964 => x"000b0ffd",
			965 => x"02c80ffd",
			966 => x"0a02d404",
			967 => x"ff150ffd",
			968 => x"015e0ffd",
			969 => x"0a027010",
			970 => x"0207f308",
			971 => x"0b049f04",
			972 => x"ff4f0ffd",
			973 => x"02140ffd",
			974 => x"0a026a04",
			975 => x"000d0ffd",
			976 => x"fd4d0ffd",
			977 => x"0207da04",
			978 => x"04fc0ffd",
			979 => x"09007704",
			980 => x"021f0ffd",
			981 => x"00f40ffd",
			982 => x"06014220",
			983 => x"02087b10",
			984 => x"0704d708",
			985 => x"0e053b04",
			986 => x"00420ffd",
			987 => x"015a0ffd",
			988 => x"040b8e04",
			989 => x"ffb90ffd",
			990 => x"fdc50ffd",
			991 => x"09007b08",
			992 => x"08035b04",
			993 => x"ffd80ffd",
			994 => x"03920ffd",
			995 => x"0b04e404",
			996 => x"ff0a0ffd",
			997 => x"fdeb0ffd",
			998 => x"09009710",
			999 => x"0d056808",
			1000 => x"02083004",
			1001 => x"019a0ffd",
			1002 => x"00470ffd",
			1003 => x"0a02d404",
			1004 => x"028a0ffd",
			1005 => x"fe7f0ffd",
			1006 => x"03055308",
			1007 => x"0a028b04",
			1008 => x"fcc10ffd",
			1009 => x"ff620ffd",
			1010 => x"09009e04",
			1011 => x"018f0ffd",
			1012 => x"005e0ffd",
			1013 => x"fe660ffd",
			1014 => x"0a024510",
			1015 => x"0f0a420c",
			1016 => x"0705a408",
			1017 => x"06010c04",
			1018 => x"feba0ffd",
			1019 => x"01cd0ffd",
			1020 => x"fe650ffd",
			1021 => x"03730ffd",
			1022 => x"fe630ffd",
			1023 => x"0e0526a8",
			1024 => x"0d05a974",
			1025 => x"0f071f40",
			1026 => x"0e04db20",
			1027 => x"0f06d610",
			1028 => x"0304c008",
			1029 => x"0b049104",
			1030 => x"00301209",
			1031 => x"ff9f1209",
			1032 => x"09007904",
			1033 => x"018f1209",
			1034 => x"00361209",
			1035 => x"01006a08",
			1036 => x"0e048804",
			1037 => x"ff9c1209",
			1038 => x"00201209",
			1039 => x"0e04bb04",
			1040 => x"ff5f1209",
			1041 => x"fd5a1209",
			1042 => x"040b3610",
			1043 => x"0f070508",
			1044 => x"06012504",
			1045 => x"fedc1209",
			1046 => x"01311209",
			1047 => x"0704bc04",
			1048 => x"00411209",
			1049 => x"fddb1209",
			1050 => x"0c04b108",
			1051 => x"0704d604",
			1052 => x"01041209",
			1053 => x"feed1209",
			1054 => x"0b04f004",
			1055 => x"02dd1209",
			1056 => x"009e1209",
			1057 => x"0c04b420",
			1058 => x"0c047210",
			1059 => x"0c045b08",
			1060 => x"0f078104",
			1061 => x"ff401209",
			1062 => x"01aa1209",
			1063 => x"06014904",
			1064 => x"02461209",
			1065 => x"00aa1209",
			1066 => x"08033c08",
			1067 => x"0d055a04",
			1068 => x"fdef1209",
			1069 => x"ffa71209",
			1070 => x"00042904",
			1071 => x"025c1209",
			1072 => x"ffc01209",
			1073 => x"0c04b504",
			1074 => x"04101209",
			1075 => x"0c04cc08",
			1076 => x"0f073b04",
			1077 => x"ff401209",
			1078 => x"fdf81209",
			1079 => x"0e04f704",
			1080 => x"ff571209",
			1081 => x"01081209",
			1082 => x"0c04ef24",
			1083 => x"0f07791c",
			1084 => x"0305a010",
			1085 => x"0e04c308",
			1086 => x"0e04b404",
			1087 => x"ff501209",
			1088 => x"002c1209",
			1089 => x"0c04cd04",
			1090 => x"fd641209",
			1091 => x"fe8a1209",
			1092 => x"0704d804",
			1093 => x"01031209",
			1094 => x"0e051004",
			1095 => x"ff951209",
			1096 => x"fdcd1209",
			1097 => x"0900be04",
			1098 => x"00501209",
			1099 => x"02c91209",
			1100 => x"0f073908",
			1101 => x"0207b504",
			1102 => x"01931209",
			1103 => x"fedd1209",
			1104 => x"0e050d04",
			1105 => x"05de1209",
			1106 => x"ffcb1209",
			1107 => x"0d058020",
			1108 => x"0208e414",
			1109 => x"01005304",
			1110 => x"fd461209",
			1111 => x"07049404",
			1112 => x"ffb41209",
			1113 => x"0b04e308",
			1114 => x"0b04d304",
			1115 => x"015e1209",
			1116 => x"ffb91209",
			1117 => x"02901209",
			1118 => x"0f07eb08",
			1119 => x"0704bc04",
			1120 => x"017e1209",
			1121 => x"fe9a1209",
			1122 => x"fe081209",
			1123 => x"0305890c",
			1124 => x"0b04d304",
			1125 => x"009a1209",
			1126 => x"01007104",
			1127 => x"fc951209",
			1128 => x"00631209",
			1129 => x"08039318",
			1130 => x"040cbf10",
			1131 => x"0003ea08",
			1132 => x"040aef04",
			1133 => x"fffa1209",
			1134 => x"feb71209",
			1135 => x"08031d04",
			1136 => x"01601209",
			1137 => x"00231209",
			1138 => x"0d059c04",
			1139 => x"00001209",
			1140 => x"fe401209",
			1141 => x"0c04cf0c",
			1142 => x"0f079604",
			1143 => x"06fb1209",
			1144 => x"0f07e304",
			1145 => x"ff0a1209",
			1146 => x"02a31209",
			1147 => x"0e064308",
			1148 => x"0704ee04",
			1149 => x"00781209",
			1150 => x"fe951209",
			1151 => x"06018d04",
			1152 => x"02481209",
			1153 => x"ff231209",
			1154 => x"0c0543ac",
			1155 => x"09007e58",
			1156 => x"0304df3c",
			1157 => x"08034520",
			1158 => x"040bb710",
			1159 => x"0c047408",
			1160 => x"08033004",
			1161 => x"01b61375",
			1162 => x"ff7f1375",
			1163 => x"0e042604",
			1164 => x"fe711375",
			1165 => x"002d1375",
			1166 => x"05050308",
			1167 => x"0207df04",
			1168 => x"00f11375",
			1169 => x"feed1375",
			1170 => x"05051404",
			1171 => x"04701375",
			1172 => x"00781375",
			1173 => x"05052e10",
			1174 => x"09007108",
			1175 => x"03045e04",
			1176 => x"ffb11375",
			1177 => x"00dd1375",
			1178 => x"08035304",
			1179 => x"fe5f1375",
			1180 => x"ffa61375",
			1181 => x"08038504",
			1182 => x"050f1375",
			1183 => x"0d055904",
			1184 => x"ff801375",
			1185 => x"02bb1375",
			1186 => x"0b04bf18",
			1187 => x"0208380c",
			1188 => x"0003f704",
			1189 => x"fef11375",
			1190 => x"08034704",
			1191 => x"03cc1375",
			1192 => x"01ac1375",
			1193 => x"00044604",
			1194 => x"fe1a1375",
			1195 => x"05052b04",
			1196 => x"009a1375",
			1197 => x"02211375",
			1198 => x"fdf61375",
			1199 => x"01004d18",
			1200 => x"05051104",
			1201 => x"00a61375",
			1202 => x"01004b08",
			1203 => x"0e048504",
			1204 => x"fe711375",
			1205 => x"fcd21375",
			1206 => x"0e048f08",
			1207 => x"00048a04",
			1208 => x"fdfa1375",
			1209 => x"ffc01375",
			1210 => x"00911375",
			1211 => x"0c047920",
			1212 => x"09008010",
			1213 => x"05051d08",
			1214 => x"0c047504",
			1215 => x"00a81375",
			1216 => x"fe3b1375",
			1217 => x"08035604",
			1218 => x"02c41375",
			1219 => x"01ab1375",
			1220 => x"0208a408",
			1221 => x"02085904",
			1222 => x"ffdd1375",
			1223 => x"ff0f1375",
			1224 => x"05051e04",
			1225 => x"02991375",
			1226 => x"ffe71375",
			1227 => x"0c049010",
			1228 => x"05056808",
			1229 => x"09009304",
			1230 => x"00841375",
			1231 => x"02121375",
			1232 => x"0b04e204",
			1233 => x"fe661375",
			1234 => x"01951375",
			1235 => x"05051004",
			1236 => x"02721375",
			1237 => x"0b049d04",
			1238 => x"fedf1375",
			1239 => x"00131375",
			1240 => x"0a024c08",
			1241 => x"020a3a04",
			1242 => x"fe8f1375",
			1243 => x"01751375",
			1244 => x"fe721375",
			1245 => x"0803298c",
			1246 => x"08031d40",
			1247 => x"0d053324",
			1248 => x"07049214",
			1249 => x"06012910",
			1250 => x"0e046808",
			1251 => x"0b048f04",
			1252 => x"00da15a1",
			1253 => x"fed615a1",
			1254 => x"040ac204",
			1255 => x"ff6715a1",
			1256 => x"021615a1",
			1257 => x"fee915a1",
			1258 => x"0207c50c",
			1259 => x"03049704",
			1260 => x"000915a1",
			1261 => x"0207a104",
			1262 => x"02e815a1",
			1263 => x"016a15a1",
			1264 => x"ff8b15a1",
			1265 => x"0e044b04",
			1266 => x"fe4f15a1",
			1267 => x"07049008",
			1268 => x"01005104",
			1269 => x"ffd915a1",
			1270 => x"028015a1",
			1271 => x"0b04b008",
			1272 => x"040b5604",
			1273 => x"fe7b15a1",
			1274 => x"007815a1",
			1275 => x"05055504",
			1276 => x"00ab15a1",
			1277 => x"fff115a1",
			1278 => x"02083828",
			1279 => x"0a026f10",
			1280 => x"0a026904",
			1281 => x"003f15a1",
			1282 => x"06013108",
			1283 => x"0b04bf04",
			1284 => x"fe9615a1",
			1285 => x"007215a1",
			1286 => x"fda015a1",
			1287 => x"01004e08",
			1288 => x"09007b04",
			1289 => x"ffb015a1",
			1290 => x"fe3515a1",
			1291 => x"05057508",
			1292 => x"0c04ae04",
			1293 => x"008a15a1",
			1294 => x"028215a1",
			1295 => x"05058504",
			1296 => x"fe6f15a1",
			1297 => x"007515a1",
			1298 => x"0b049008",
			1299 => x"0c044304",
			1300 => x"000015a1",
			1301 => x"028d15a1",
			1302 => x"0100620c",
			1303 => x"0704a804",
			1304 => x"fd3415a1",
			1305 => x"0e04e204",
			1306 => x"fdff15a1",
			1307 => x"ffb415a1",
			1308 => x"0d058308",
			1309 => x"01006604",
			1310 => x"005415a1",
			1311 => x"022a15a1",
			1312 => x"01007904",
			1313 => x"fe7215a1",
			1314 => x"000615a1",
			1315 => x"08032e34",
			1316 => x"06015628",
			1317 => x"040b8a14",
			1318 => x"0d05670c",
			1319 => x"0b04ae04",
			1320 => x"014f15a1",
			1321 => x"040b5004",
			1322 => x"011a15a1",
			1323 => x"fecf15a1",
			1324 => x"02087e04",
			1325 => x"021215a1",
			1326 => x"011815a1",
			1327 => x"02084d0c",
			1328 => x"040ba404",
			1329 => x"003015a1",
			1330 => x"06012904",
			1331 => x"009815a1",
			1332 => x"02ac15a1",
			1333 => x"07049504",
			1334 => x"01a515a1",
			1335 => x"fe1d15a1",
			1336 => x"02096c04",
			1337 => x"fda815a1",
			1338 => x"0307c404",
			1339 => x"021f15a1",
			1340 => x"000015a1",
			1341 => x"0505f640",
			1342 => x"0900b920",
			1343 => x"01006c10",
			1344 => x"0208d008",
			1345 => x"03057904",
			1346 => x"000e15a1",
			1347 => x"007c15a1",
			1348 => x"0704da04",
			1349 => x"ff5e15a1",
			1350 => x"00a915a1",
			1351 => x"0b04d208",
			1352 => x"0900b104",
			1353 => x"fd6a15a1",
			1354 => x"004815a1",
			1355 => x"0900a904",
			1356 => x"025d15a1",
			1357 => x"009515a1",
			1358 => x"0e05bb10",
			1359 => x"0c04ef08",
			1360 => x"08033304",
			1361 => x"fd1915a1",
			1362 => x"ff5115a1",
			1363 => x"040c2c04",
			1364 => x"01b215a1",
			1365 => x"feb215a1",
			1366 => x"0900d308",
			1367 => x"06015b04",
			1368 => x"fff115a1",
			1369 => x"014515a1",
			1370 => x"0a029204",
			1371 => x"00ed15a1",
			1372 => x"ff0815a1",
			1373 => x"040cbf14",
			1374 => x"0e05c304",
			1375 => x"035f15a1",
			1376 => x"040b8508",
			1377 => x"07050304",
			1378 => x"01c015a1",
			1379 => x"ff1015a1",
			1380 => x"0c04cf04",
			1381 => x"ff5b15a1",
			1382 => x"015c15a1",
			1383 => x"fe7f15a1",
			1384 => x"050606b0",
			1385 => x"040c7f60",
			1386 => x"0e048f30",
			1387 => x"0e046114",
			1388 => x"04098704",
			1389 => x"06611775",
			1390 => x"06013e08",
			1391 => x"0b048e04",
			1392 => x"01331775",
			1393 => x"ffbf1775",
			1394 => x"00048a04",
			1395 => x"03021775",
			1396 => x"fee81775",
			1397 => x"08030a0c",
			1398 => x"06012b08",
			1399 => x"05053c04",
			1400 => x"00911775",
			1401 => x"fe721775",
			1402 => x"03401775",
			1403 => x"0207da08",
			1404 => x"00040c04",
			1405 => x"028b1775",
			1406 => x"07151775",
			1407 => x"09008004",
			1408 => x"04571775",
			1409 => x"01651775",
			1410 => x"06011f10",
			1411 => x"0802e80c",
			1412 => x"03051b04",
			1413 => x"fff31775",
			1414 => x"0c047504",
			1415 => x"feef1775",
			1416 => x"fe441775",
			1417 => x"02ad1775",
			1418 => x"040bd810",
			1419 => x"06017408",
			1420 => x"06013504",
			1421 => x"02f11775",
			1422 => x"04b81775",
			1423 => x"0a02b804",
			1424 => x"fe311775",
			1425 => x"01541775",
			1426 => x"0c04d208",
			1427 => x"0e052604",
			1428 => x"024d1775",
			1429 => x"03ee1775",
			1430 => x"02091b04",
			1431 => x"ffd41775",
			1432 => x"02c51775",
			1433 => x"06013414",
			1434 => x"040ca704",
			1435 => x"02551775",
			1436 => x"01003904",
			1437 => x"fe3a1775",
			1438 => x"09006c08",
			1439 => x"040ce104",
			1440 => x"fe781775",
			1441 => x"00771775",
			1442 => x"fe631775",
			1443 => x"0b04b920",
			1444 => x"00049a10",
			1445 => x"0c047608",
			1446 => x"040cb604",
			1447 => x"03e31775",
			1448 => x"07a41775",
			1449 => x"05053a04",
			1450 => x"02991775",
			1451 => x"ff3f1775",
			1452 => x"040d6e08",
			1453 => x"09006804",
			1454 => x"03011775",
			1455 => x"00281775",
			1456 => x"0a031504",
			1457 => x"04a41775",
			1458 => x"fe421775",
			1459 => x"0f07eb10",
			1460 => x"02087608",
			1461 => x"03053704",
			1462 => x"ff9b1775",
			1463 => x"03e21775",
			1464 => x"0c047504",
			1465 => x"01881775",
			1466 => x"fee61775",
			1467 => x"00048a04",
			1468 => x"fe361775",
			1469 => x"040ce104",
			1470 => x"03af1775",
			1471 => x"ff5d1775",
			1472 => x"0c054324",
			1473 => x"05070d20",
			1474 => x"03066904",
			1475 => x"fe4f1775",
			1476 => x"0601640c",
			1477 => x"06013104",
			1478 => x"fe581775",
			1479 => x"0208b404",
			1480 => x"05ca1775",
			1481 => x"01e01775",
			1482 => x"06017908",
			1483 => x"02092004",
			1484 => x"fee41775",
			1485 => x"00c51775",
			1486 => x"0c04b904",
			1487 => x"ff6a1775",
			1488 => x"fe4b1775",
			1489 => x"05c61775",
			1490 => x"0c054814",
			1491 => x"08035210",
			1492 => x"0803410c",
			1493 => x"0802c704",
			1494 => x"fe631775",
			1495 => x"08030804",
			1496 => x"00981775",
			1497 => x"fe8d1775",
			1498 => x"01ee1775",
			1499 => x"fe4e1775",
			1500 => x"fe3a1775",
			1501 => x"0208bb8c",
			1502 => x"040d5560",
			1503 => x"06015840",
			1504 => x"06014a20",
			1505 => x"06014910",
			1506 => x"0207da08",
			1507 => x"06012d04",
			1508 => x"00021999",
			1509 => x"00bd1999",
			1510 => x"06013504",
			1511 => x"ffb71999",
			1512 => x"00131999",
			1513 => x"040b9d08",
			1514 => x"01006904",
			1515 => x"fef51999",
			1516 => x"00c51999",
			1517 => x"08035504",
			1518 => x"fd4c1999",
			1519 => x"ff841999",
			1520 => x"03056f10",
			1521 => x"01006508",
			1522 => x"03055304",
			1523 => x"002d1999",
			1524 => x"01431999",
			1525 => x"08037604",
			1526 => x"fdc11999",
			1527 => x"002d1999",
			1528 => x"0c04cb08",
			1529 => x"0e050704",
			1530 => x"00421999",
			1531 => x"01291999",
			1532 => x"06015604",
			1533 => x"00851999",
			1534 => x"fe7d1999",
			1535 => x"0803310c",
			1536 => x"0c04ed08",
			1537 => x"08031d04",
			1538 => x"ff0c1999",
			1539 => x"fbd11999",
			1540 => x"00901999",
			1541 => x"0a029204",
			1542 => x"035e1999",
			1543 => x"0704d408",
			1544 => x"0208a404",
			1545 => x"ff8b1999",
			1546 => x"01f21999",
			1547 => x"0d058e04",
			1548 => x"01581999",
			1549 => x"fefa1999",
			1550 => x"01005524",
			1551 => x"0d05421c",
			1552 => x"00052910",
			1553 => x"03046f08",
			1554 => x"0a02db04",
			1555 => x"ff351999",
			1556 => x"01f11999",
			1557 => x"06012b04",
			1558 => x"00001999",
			1559 => x"03131999",
			1560 => x"040eab04",
			1561 => x"fe471999",
			1562 => x"040fc604",
			1563 => x"01441999",
			1564 => x"fea21999",
			1565 => x"0e041604",
			1566 => x"fe511999",
			1567 => x"fffd1999",
			1568 => x"0c04b204",
			1569 => x"06ba1999",
			1570 => x"fee31999",
			1571 => x"06014f4c",
			1572 => x"0f07d528",
			1573 => x"0e057120",
			1574 => x"00045310",
			1575 => x"0b04b008",
			1576 => x"0c045c04",
			1577 => x"00001999",
			1578 => x"00e61999",
			1579 => x"0704c004",
			1580 => x"fd2b1999",
			1581 => x"fe6e1999",
			1582 => x"0704be08",
			1583 => x"0d054f04",
			1584 => x"ff681999",
			1585 => x"01161999",
			1586 => x"0704d804",
			1587 => x"fe121999",
			1588 => x"00241999",
			1589 => x"01006d04",
			1590 => x"02191999",
			1591 => x"ff3b1999",
			1592 => x"0e050d04",
			1593 => x"047d1999",
			1594 => x"0d05de10",
			1595 => x"0c04b208",
			1596 => x"08031204",
			1597 => x"01d01999",
			1598 => x"fe401999",
			1599 => x"00044a04",
			1600 => x"fc981999",
			1601 => x"fdc51999",
			1602 => x"06014d08",
			1603 => x"040a3a04",
			1604 => x"fff11999",
			1605 => x"fe581999",
			1606 => x"0208f904",
			1607 => x"019e1999",
			1608 => x"ff2d1999",
			1609 => x"06017d30",
			1610 => x"0f078110",
			1611 => x"06015308",
			1612 => x"03055f04",
			1613 => x"fe821999",
			1614 => x"01981999",
			1615 => x"01006f04",
			1616 => x"fe261999",
			1617 => x"00001999",
			1618 => x"08035b10",
			1619 => x"040b9108",
			1620 => x"0d05de04",
			1621 => x"01f11999",
			1622 => x"ffcf1999",
			1623 => x"0208c904",
			1624 => x"00b71999",
			1625 => x"fe7f1999",
			1626 => x"040c2408",
			1627 => x"0f084604",
			1628 => x"00951999",
			1629 => x"02281999",
			1630 => x"00047004",
			1631 => x"ff1a1999",
			1632 => x"00461999",
			1633 => x"0d060f08",
			1634 => x"02096004",
			1635 => x"ff6c1999",
			1636 => x"013d1999",
			1637 => x"fe5b1999",
			1638 => x"0c04d0ac",
			1639 => x"0c04b470",
			1640 => x"0208d638",
			1641 => x"01007520",
			1642 => x"0704c110",
			1643 => x"0704ad08",
			1644 => x"0704aa04",
			1645 => x"000e1c0d",
			1646 => x"ff571c0d",
			1647 => x"0e057104",
			1648 => x"00431c0d",
			1649 => x"01991c0d",
			1650 => x"0704c208",
			1651 => x"0a02bb04",
			1652 => x"fe981c0d",
			1653 => x"00f21c0d",
			1654 => x"08038204",
			1655 => x"ffe71c0d",
			1656 => x"00f91c0d",
			1657 => x"0900d610",
			1658 => x"0704ee08",
			1659 => x"040a4904",
			1660 => x"ff571c0d",
			1661 => x"01451c0d",
			1662 => x"0a029604",
			1663 => x"fea41c0d",
			1664 => x"00e91c0d",
			1665 => x"0e061e04",
			1666 => x"fe151c0d",
			1667 => x"00151c0d",
			1668 => x"0900b520",
			1669 => x"0f07ce10",
			1670 => x"0a02b608",
			1671 => x"08034a04",
			1672 => x"00d91c0d",
			1673 => x"fe691c0d",
			1674 => x"0e04e204",
			1675 => x"fe941c0d",
			1676 => x"00841c0d",
			1677 => x"0f080e08",
			1678 => x"0c049204",
			1679 => x"ffd11c0d",
			1680 => x"01931c0d",
			1681 => x"0f083904",
			1682 => x"fe411c0d",
			1683 => x"00001c0d",
			1684 => x"040b7808",
			1685 => x"040b4604",
			1686 => x"fef81c0d",
			1687 => x"019b1c0d",
			1688 => x"08036908",
			1689 => x"01007d04",
			1690 => x"fdf71c0d",
			1691 => x"00001c0d",
			1692 => x"040c6004",
			1693 => x"003f1c0d",
			1694 => x"fe4f1c0d",
			1695 => x"0c04b518",
			1696 => x"040bbd0c",
			1697 => x"03058004",
			1698 => x"feb31c0d",
			1699 => x"0e05a404",
			1700 => x"01dc1c0d",
			1701 => x"00401c0d",
			1702 => x"0b04f208",
			1703 => x"08037604",
			1704 => x"03801c0d",
			1705 => x"02321c0d",
			1706 => x"00e01c0d",
			1707 => x"0802fb10",
			1708 => x"0a024508",
			1709 => x"0900c804",
			1710 => x"fe831c0d",
			1711 => x"015f1c0d",
			1712 => x"01007804",
			1713 => x"010c1c0d",
			1714 => x"022a1c0d",
			1715 => x"0a026208",
			1716 => x"0a025e04",
			1717 => x"00681c0d",
			1718 => x"fcc31c0d",
			1719 => x"0a026a04",
			1720 => x"023e1c0d",
			1721 => x"08033104",
			1722 => x"ff8b1c0d",
			1723 => x"00481c0d",
			1724 => x"0c04d138",
			1725 => x"0704d60c",
			1726 => x"0704d204",
			1727 => x"fe811c0d",
			1728 => x"0f076504",
			1729 => x"00731c0d",
			1730 => x"020c1c0d",
			1731 => x"01007918",
			1732 => x"0208d610",
			1733 => x"0900b108",
			1734 => x"0b04f304",
			1735 => x"fe4c1c0d",
			1736 => x"fc941c0d",
			1737 => x"01007304",
			1738 => x"ffb11c0d",
			1739 => x"fd8b1c0d",
			1740 => x"05059304",
			1741 => x"fe4b1c0d",
			1742 => x"00001c0d",
			1743 => x"0e05e908",
			1744 => x"07050404",
			1745 => x"01c81c0d",
			1746 => x"ffb51c0d",
			1747 => x"0f087208",
			1748 => x"0003fb04",
			1749 => x"fcf91c0d",
			1750 => x"febe1c0d",
			1751 => x"008c1c0d",
			1752 => x"0c04d21c",
			1753 => x"05058608",
			1754 => x"05057604",
			1755 => x"01421c0d",
			1756 => x"02ac1c0d",
			1757 => x"0505a004",
			1758 => x"fef61c0d",
			1759 => x"0505df08",
			1760 => x"0e058e04",
			1761 => x"00ab1c0d",
			1762 => x"023a1c0d",
			1763 => x"0f085c04",
			1764 => x"fe441c0d",
			1765 => x"00bb1c0d",
			1766 => x"0c04ea1c",
			1767 => x"0c04e910",
			1768 => x"0e05d808",
			1769 => x"0704ee04",
			1770 => x"fff51c0d",
			1771 => x"fe8c1c0d",
			1772 => x"0208dd04",
			1773 => x"02281c0d",
			1774 => x"fe861c0d",
			1775 => x"0e056804",
			1776 => x"00101c0d",
			1777 => x"02093504",
			1778 => x"fdb11c0d",
			1779 => x"00381c0d",
			1780 => x"0c04ec10",
			1781 => x"0306c508",
			1782 => x"0e058704",
			1783 => x"ffdd1c0d",
			1784 => x"02031c0d",
			1785 => x"0100ad04",
			1786 => x"fe5f1c0d",
			1787 => x"010b1c0d",
			1788 => x"0c04ed08",
			1789 => x"02099504",
			1790 => x"fe6f1c0d",
			1791 => x"01991c0d",
			1792 => x"0505bd04",
			1793 => x"00ec1c0d",
			1794 => x"ffeb1c0d",
			1795 => x"0c04f1dc",
			1796 => x"0c047974",
			1797 => x"09008c40",
			1798 => x"03050020",
			1799 => x"09007e10",
			1800 => x"03049f08",
			1801 => x"0f069904",
			1802 => x"ffff1e59",
			1803 => x"fe761e59",
			1804 => x"05051104",
			1805 => x"00b91e59",
			1806 => x"ffbc1e59",
			1807 => x"040b6908",
			1808 => x"0e045304",
			1809 => x"ff1e1e59",
			1810 => x"01c01e59",
			1811 => x"0a029604",
			1812 => x"fe881e59",
			1813 => x"ffbf1e59",
			1814 => x"0f070510",
			1815 => x"0e048f08",
			1816 => x"07049304",
			1817 => x"ffd11e59",
			1818 => x"01b61e59",
			1819 => x"06012004",
			1820 => x"00001e59",
			1821 => x"02601e59",
			1822 => x"0a029e08",
			1823 => x"0e04c904",
			1824 => x"fee61e59",
			1825 => x"00711e59",
			1826 => x"0a02be04",
			1827 => x"015b1e59",
			1828 => x"fe8a1e59",
			1829 => x"05052d14",
			1830 => x"0b04ae0c",
			1831 => x"0c047808",
			1832 => x"0e04b404",
			1833 => x"fe0a1e59",
			1834 => x"fffe1e59",
			1835 => x"00fd1e59",
			1836 => x"09009504",
			1837 => x"fe8f1e59",
			1838 => x"fc9a1e59",
			1839 => x"0a027810",
			1840 => x"040ae808",
			1841 => x"0a025304",
			1842 => x"ff581e59",
			1843 => x"015c1e59",
			1844 => x"02081504",
			1845 => x"fdff1e59",
			1846 => x"ff6d1e59",
			1847 => x"0c047308",
			1848 => x"05055504",
			1849 => x"01aa1e59",
			1850 => x"fee01e59",
			1851 => x"02084404",
			1852 => x"00971e59",
			1853 => x"ff741e59",
			1854 => x"0c048f28",
			1855 => x"040b9114",
			1856 => x"0c047b0c",
			1857 => x"07049304",
			1858 => x"018a1e59",
			1859 => x"0704bc04",
			1860 => x"fddf1e59",
			1861 => x"00001e59",
			1862 => x"09009504",
			1863 => x"ffe11e59",
			1864 => x"02081e59",
			1865 => x"0b047104",
			1866 => x"fe481e59",
			1867 => x"02089808",
			1868 => x"0e049604",
			1869 => x"01021e59",
			1870 => x"028a1e59",
			1871 => x"0e050704",
			1872 => x"fee21e59",
			1873 => x"01491e59",
			1874 => x"03052520",
			1875 => x"09009510",
			1876 => x"0d056608",
			1877 => x"05054b04",
			1878 => x"ffff1e59",
			1879 => x"fee01e59",
			1880 => x"0f06ca04",
			1881 => x"01ca1e59",
			1882 => x"feca1e59",
			1883 => x"0f06ac08",
			1884 => x"03050004",
			1885 => x"fe841e59",
			1886 => x"00ad1e59",
			1887 => x"02082a04",
			1888 => x"fdac1e59",
			1889 => x"ffb71e59",
			1890 => x"09009c10",
			1891 => x"0c049608",
			1892 => x"0d058304",
			1893 => x"003d1e59",
			1894 => x"fd761e59",
			1895 => x"05053a04",
			1896 => x"02251e59",
			1897 => x"009b1e59",
			1898 => x"0e04e908",
			1899 => x"0a029804",
			1900 => x"fff11e59",
			1901 => x"fee91e59",
			1902 => x"0f074f04",
			1903 => x"006f1e59",
			1904 => x"fffa1e59",
			1905 => x"0f07ce18",
			1906 => x"0506160c",
			1907 => x"0e054408",
			1908 => x"040bd804",
			1909 => x"01201e59",
			1910 => x"fe7f1e59",
			1911 => x"fddf1e59",
			1912 => x"05061908",
			1913 => x"06014e04",
			1914 => x"00001e59",
			1915 => x"03011e59",
			1916 => x"feda1e59",
			1917 => x"06015c18",
			1918 => x"040b8a14",
			1919 => x"0208a408",
			1920 => x"0705a104",
			1921 => x"01b31e59",
			1922 => x"ffb91e59",
			1923 => x"09017604",
			1924 => x"fe5f1e59",
			1925 => x"0a021d04",
			1926 => x"ff2f1e59",
			1927 => x"01081e59",
			1928 => x"02f61e59",
			1929 => x"0a02cc10",
			1930 => x"0b057404",
			1931 => x"fe331e59",
			1932 => x"0900f704",
			1933 => x"01291e59",
			1934 => x"02092e04",
			1935 => x"fff11e59",
			1936 => x"fe9a1e59",
			1937 => x"0f083908",
			1938 => x"07053104",
			1939 => x"041f1e59",
			1940 => x"00001e59",
			1941 => x"feb11e59",
			1942 => x"09007b88",
			1943 => x"05051d48",
			1944 => x"05051440",
			1945 => x"02082a20",
			1946 => x"03049710",
			1947 => x"0b049d08",
			1948 => x"0a02dd04",
			1949 => x"001220bd",
			1950 => x"011120bd",
			1951 => x"06012b04",
			1952 => x"ffec20bd",
			1953 => x"fe7420bd",
			1954 => x"07047b08",
			1955 => x"0304be04",
			1956 => x"feca20bd",
			1957 => x"ffb420bd",
			1958 => x"0b048d04",
			1959 => x"01c320bd",
			1960 => x"00b020bd",
			1961 => x"01004710",
			1962 => x"0304be08",
			1963 => x"0c045c04",
			1964 => x"008e20bd",
			1965 => x"fe8c20bd",
			1966 => x"0304c004",
			1967 => x"021e20bd",
			1968 => x"000420bd",
			1969 => x"0b049008",
			1970 => x"08037e04",
			1971 => x"fdf620bd",
			1972 => x"ffab20bd",
			1973 => x"0c047a04",
			1974 => x"00c820bd",
			1975 => x"fec020bd",
			1976 => x"0f064a04",
			1977 => x"004920bd",
			1978 => x"fe3f20bd",
			1979 => x"06013424",
			1980 => x"0d051b0c",
			1981 => x"0c049308",
			1982 => x"08033904",
			1983 => x"013620bd",
			1984 => x"fe7c20bd",
			1985 => x"025120bd",
			1986 => x"01004710",
			1987 => x"08033108",
			1988 => x"0207b704",
			1989 => x"ff5920bd",
			1990 => x"023420bd",
			1991 => x"0208c004",
			1992 => x"fe5a20bd",
			1993 => x"002e20bd",
			1994 => x"0b04a204",
			1995 => x"fe3820bd",
			1996 => x"ff7520bd",
			1997 => x"0704c018",
			1998 => x"0e04360c",
			1999 => x"0f06d008",
			2000 => x"02080e04",
			2001 => x"002020bd",
			2002 => x"019a20bd",
			2003 => x"fe5220bd",
			2004 => x"0d051b04",
			2005 => x"005320bd",
			2006 => x"0d053304",
			2007 => x"02a520bd",
			2008 => x"016620bd",
			2009 => x"fead20bd",
			2010 => x"0305334c",
			2011 => x"03052f34",
			2012 => x"03052b20",
			2013 => x"09009b10",
			2014 => x"0c047808",
			2015 => x"0b04b004",
			2016 => x"ffd420bd",
			2017 => x"fefb20bd",
			2018 => x"0c049304",
			2019 => x"004d20bd",
			2020 => x"ffd220bd",
			2021 => x"09009d08",
			2022 => x"0a02ae04",
			2023 => x"fdf120bd",
			2024 => x"fff420bd",
			2025 => x"0f06e304",
			2026 => x"fffc20bd",
			2027 => x"fe3d20bd",
			2028 => x"0601410c",
			2029 => x"0c049608",
			2030 => x"0c048f04",
			2031 => x"004820bd",
			2032 => x"fe9620bd",
			2033 => x"015020bd",
			2034 => x"02088904",
			2035 => x"020120bd",
			2036 => x"00af20bd",
			2037 => x"0a028208",
			2038 => x"06013204",
			2039 => x"fea720bd",
			2040 => x"007720bd",
			2041 => x"0a02a908",
			2042 => x"0b04bf04",
			2043 => x"fe8220bd",
			2044 => x"fd8420bd",
			2045 => x"02087604",
			2046 => x"005720bd",
			2047 => x"fe5e20bd",
			2048 => x"09009330",
			2049 => x"0f071f14",
			2050 => x"0a026708",
			2051 => x"0f06d904",
			2052 => x"009720bd",
			2053 => x"ffb820bd",
			2054 => x"09008904",
			2055 => x"002220bd",
			2056 => x"0b04be04",
			2057 => x"014c20bd",
			2058 => x"024a20bd",
			2059 => x"05055710",
			2060 => x"0c047608",
			2061 => x"03054f04",
			2062 => x"023120bd",
			2063 => x"004f20bd",
			2064 => x"0c049804",
			2065 => x"ffc420bd",
			2066 => x"014520bd",
			2067 => x"09008d04",
			2068 => x"000020bd",
			2069 => x"0e04f904",
			2070 => x"fdab20bd",
			2071 => x"ff5e20bd",
			2072 => x"0c047414",
			2073 => x"09009804",
			2074 => x"fe6720bd",
			2075 => x"0f074908",
			2076 => x"0d056604",
			2077 => x"01dc20bd",
			2078 => x"ff4520bd",
			2079 => x"02088904",
			2080 => x"fdef20bd",
			2081 => x"000020bd",
			2082 => x"0c04760c",
			2083 => x"0704a804",
			2084 => x"ff5520bd",
			2085 => x"05056704",
			2086 => x"00f720bd",
			2087 => x"029520bd",
			2088 => x"03055308",
			2089 => x"03054f04",
			2090 => x"fff020bd",
			2091 => x"fea520bd",
			2092 => x"0900a804",
			2093 => x"005220bd",
			2094 => x"fffa20bd",
			2095 => x"0e053ba4",
			2096 => x"0f06d654",
			2097 => x"06012524",
			2098 => x"0d054e18",
			2099 => x"0304ef10",
			2100 => x"06011c08",
			2101 => x"0d052504",
			2102 => x"015d2341",
			2103 => x"ff7f2341",
			2104 => x"07047804",
			2105 => x"01ad2341",
			2106 => x"fedd2341",
			2107 => x"0e047104",
			2108 => x"00642341",
			2109 => x"02422341",
			2110 => x"0e04f004",
			2111 => x"fe452341",
			2112 => x"0e050d04",
			2113 => x"00002341",
			2114 => x"ff472341",
			2115 => x"03053320",
			2116 => x"02079b10",
			2117 => x"02077708",
			2118 => x"07049404",
			2119 => x"fe672341",
			2120 => x"009d2341",
			2121 => x"0f062f04",
			2122 => x"00602341",
			2123 => x"02242341",
			2124 => x"09009a08",
			2125 => x"03051b04",
			2126 => x"00162341",
			2127 => x"017a2341",
			2128 => x"0f06a504",
			2129 => x"008e2341",
			2130 => x"fe0e2341",
			2131 => x"0d05a90c",
			2132 => x"09009504",
			2133 => x"00032341",
			2134 => x"01006404",
			2135 => x"01562341",
			2136 => x"02622341",
			2137 => x"ffdd2341",
			2138 => x"0900bc3c",
			2139 => x"0305101c",
			2140 => x"0900820c",
			2141 => x"0704aa08",
			2142 => x"0304f704",
			2143 => x"ffc12341",
			2144 => x"00f12341",
			2145 => x"fdff2341",
			2146 => x"01005308",
			2147 => x"0f06ed04",
			2148 => x"ff942341",
			2149 => x"fde82341",
			2150 => x"0d054d04",
			2151 => x"001a2341",
			2152 => x"febc2341",
			2153 => x"09009810",
			2154 => x"0a029008",
			2155 => x"02082f04",
			2156 => x"00592341",
			2157 => x"ff772341",
			2158 => x"0208d004",
			2159 => x"00a42341",
			2160 => x"ffa32341",
			2161 => x"03054308",
			2162 => x"0f070904",
			2163 => x"ff812341",
			2164 => x"fde02341",
			2165 => x"0f074f04",
			2166 => x"00282341",
			2167 => x"ff922341",
			2168 => x"01007604",
			2169 => x"fd842341",
			2170 => x"0f077908",
			2171 => x"0e052604",
			2172 => x"fdee2341",
			2173 => x"ffea2341",
			2174 => x"020a0004",
			2175 => x"034e2341",
			2176 => x"00002341",
			2177 => x"0003ea54",
			2178 => x"040abb2c",
			2179 => x"0003d11c",
			2180 => x"0802f910",
			2181 => x"0a024108",
			2182 => x"040a0104",
			2183 => x"00382341",
			2184 => x"fe812341",
			2185 => x"0704ec04",
			2186 => x"01f12341",
			2187 => x"fff32341",
			2188 => x"0900c404",
			2189 => x"fce72341",
			2190 => x"0e065a04",
			2191 => x"00ba2341",
			2192 => x"fdef2341",
			2193 => x"040a5b04",
			2194 => x"fe632341",
			2195 => x"05058504",
			2196 => x"00292341",
			2197 => x"0208f204",
			2198 => x"023c2341",
			2199 => x"00002341",
			2200 => x"0704ed14",
			2201 => x"0505b110",
			2202 => x"0305b908",
			2203 => x"0802f804",
			2204 => x"fe842341",
			2205 => x"00912341",
			2206 => x"08030a04",
			2207 => x"fe342341",
			2208 => x"fc412341",
			2209 => x"007d2341",
			2210 => x"0505bd04",
			2211 => x"01ba2341",
			2212 => x"02090c08",
			2213 => x"040adc04",
			2214 => x"ff812341",
			2215 => x"fd9e2341",
			2216 => x"07064004",
			2217 => x"00e02341",
			2218 => x"fee42341",
			2219 => x"08031d14",
			2220 => x"040b560c",
			2221 => x"01006d08",
			2222 => x"0f079104",
			2223 => x"01d52341",
			2224 => x"00512341",
			2225 => x"02182341",
			2226 => x"00040804",
			2227 => x"fe372341",
			2228 => x"026e2341",
			2229 => x"0900c41c",
			2230 => x"0004100c",
			2231 => x"02088b08",
			2232 => x"0e054b04",
			2233 => x"fdd72341",
			2234 => x"00b12341",
			2235 => x"fdaf2341",
			2236 => x"0208eb08",
			2237 => x"0f07ce04",
			2238 => x"008c2341",
			2239 => x"01e02341",
			2240 => x"08036b04",
			2241 => x"ff2d2341",
			2242 => x"00732341",
			2243 => x"03061910",
			2244 => x"00041808",
			2245 => x"0f079104",
			2246 => x"01db2341",
			2247 => x"fff02341",
			2248 => x"040c9a04",
			2249 => x"fe932341",
			2250 => x"02772341",
			2251 => x"0f08f008",
			2252 => x"0d06af04",
			2253 => x"00512341",
			2254 => x"03112341",
			2255 => x"fe622341",
			2256 => x"050606c0",
			2257 => x"040c7f74",
			2258 => x"0e048834",
			2259 => x"03050014",
			2260 => x"00048e10",
			2261 => x"06013e08",
			2262 => x"0b048e04",
			2263 => x"01732555",
			2264 => x"00022555",
			2265 => x"00046304",
			2266 => x"04e42555",
			2267 => x"01782555",
			2268 => x"fe2e2555",
			2269 => x"09008f10",
			2270 => x"06013508",
			2271 => x"0207e504",
			2272 => x"03712555",
			2273 => x"fffc2555",
			2274 => x"0f06fb04",
			2275 => x"062a2555",
			2276 => x"022e2555",
			2277 => x"00043a08",
			2278 => x"0802fc04",
			2279 => x"ff102555",
			2280 => x"02a22555",
			2281 => x"03052b04",
			2282 => x"ff0c2555",
			2283 => x"01d32555",
			2284 => x"06012520",
			2285 => x"0802e810",
			2286 => x"0a023008",
			2287 => x"0c049304",
			2288 => x"ff0d2555",
			2289 => x"fe462555",
			2290 => x"040a6904",
			2291 => x"03b52555",
			2292 => x"fed92555",
			2293 => x"09009508",
			2294 => x"040b3604",
			2295 => x"055f2555",
			2296 => x"fe602555",
			2297 => x"0c049504",
			2298 => x"fe522555",
			2299 => x"ff862555",
			2300 => x"02085410",
			2301 => x"0e04d308",
			2302 => x"09009b04",
			2303 => x"037c2555",
			2304 => x"01a32555",
			2305 => x"06015a04",
			2306 => x"04462555",
			2307 => x"00982555",
			2308 => x"0e051d08",
			2309 => x"0c049304",
			2310 => x"02552555",
			2311 => x"00d52555",
			2312 => x"0b051204",
			2313 => x"03772555",
			2314 => x"019e2555",
			2315 => x"06013410",
			2316 => x"040ca704",
			2317 => x"02062555",
			2318 => x"01003904",
			2319 => x"fe412555",
			2320 => x"08037c04",
			2321 => x"fe552555",
			2322 => x"00f82555",
			2323 => x"0b04b920",
			2324 => x"02081b10",
			2325 => x"0b048e08",
			2326 => x"03046f04",
			2327 => x"005e2555",
			2328 => x"03eb2555",
			2329 => x"03048f04",
			2330 => x"fed52555",
			2331 => x"00c62555",
			2332 => x"09006f08",
			2333 => x"06014704",
			2334 => x"05412555",
			2335 => x"ff1f2555",
			2336 => x"0c04b304",
			2337 => x"01142555",
			2338 => x"06fc2555",
			2339 => x"0f082b10",
			2340 => x"02087608",
			2341 => x"0004ab04",
			2342 => x"01652555",
			2343 => x"fed02555",
			2344 => x"0a02c304",
			2345 => x"fe9e2555",
			2346 => x"ff982555",
			2347 => x"0b054308",
			2348 => x"03065004",
			2349 => x"ff6f2555",
			2350 => x"05012555",
			2351 => x"fe5c2555",
			2352 => x"0c054334",
			2353 => x"03066904",
			2354 => x"fe532555",
			2355 => x"06016414",
			2356 => x"06013104",
			2357 => x"fe5e2555",
			2358 => x"05061508",
			2359 => x"06015f04",
			2360 => x"01dd2555",
			2361 => x"ff452555",
			2362 => x"0b05d804",
			2363 => x"03912555",
			2364 => x"06af2555",
			2365 => x"06017910",
			2366 => x"02092008",
			2367 => x"09010604",
			2368 => x"fe452555",
			2369 => x"ffbf2555",
			2370 => x"02099a04",
			2371 => x"02522555",
			2372 => x"fe5f2555",
			2373 => x"0c04b904",
			2374 => x"ff862555",
			2375 => x"06017d04",
			2376 => x"fee12555",
			2377 => x"fe3f2555",
			2378 => x"0c054814",
			2379 => x"08035210",
			2380 => x"0803410c",
			2381 => x"0802c704",
			2382 => x"fe6b2555",
			2383 => x"08030804",
			2384 => x"00802555",
			2385 => x"fe962555",
			2386 => x"01aa2555",
			2387 => x"fe552555",
			2388 => x"fe422555",
			2389 => x"09008f80",
			2390 => x"01005a70",
			2391 => x"05055540",
			2392 => x"0b04af20",
			2393 => x"0803a310",
			2394 => x"040cf508",
			2395 => x"00049a04",
			2396 => x"00222759",
			2397 => x"ff7e2759",
			2398 => x"0f064204",
			2399 => x"fe722759",
			2400 => x"01492759",
			2401 => x"0f069908",
			2402 => x"02081d04",
			2403 => x"ff5c2759",
			2404 => x"01852759",
			2405 => x"01003904",
			2406 => x"00412759",
			2407 => x"fe152759",
			2408 => x"0e046110",
			2409 => x"09008208",
			2410 => x"0a02b004",
			2411 => x"ff6e2759",
			2412 => x"026d2759",
			2413 => x"07049304",
			2414 => x"00c62759",
			2415 => x"fee52759",
			2416 => x"02088508",
			2417 => x"06014104",
			2418 => x"01172759",
			2419 => x"02482759",
			2420 => x"06014604",
			2421 => x"feac2759",
			2422 => x"00bb2759",
			2423 => x"06014614",
			2424 => x"0d054e04",
			2425 => x"00522759",
			2426 => x"0704c008",
			2427 => x"040b2904",
			2428 => x"ff2b2759",
			2429 => x"fdcc2759",
			2430 => x"040bf104",
			2431 => x"003d2759",
			2432 => x"fdd92759",
			2433 => x"02084b0c",
			2434 => x"02080704",
			2435 => x"00002759",
			2436 => x"08056404",
			2437 => x"02882759",
			2438 => x"00002759",
			2439 => x"02090c08",
			2440 => x"02088b04",
			2441 => x"001b2759",
			2442 => x"fe502759",
			2443 => x"0a038504",
			2444 => x"03c32759",
			2445 => x"ffb12759",
			2446 => x"05053b04",
			2447 => x"ff6b2759",
			2448 => x"02085208",
			2449 => x"0b04bf04",
			2450 => x"02ac2759",
			2451 => x"00382759",
			2452 => x"03b62759",
			2453 => x"0100550c",
			2454 => x"0b04b908",
			2455 => x"07049504",
			2456 => x"fff32759",
			2457 => x"fdec2759",
			2458 => x"fcec2759",
			2459 => x"0e04963c",
			2460 => x"0b04b21c",
			2461 => x"040bec10",
			2462 => x"040b7008",
			2463 => x"0704a604",
			2464 => x"000a2759",
			2465 => x"fdad2759",
			2466 => x"01005904",
			2467 => x"01702759",
			2468 => x"034f2759",
			2469 => x"040c8c08",
			2470 => x"0f06f904",
			2471 => x"fdc62759",
			2472 => x"ff9a2759",
			2473 => x"00c22759",
			2474 => x"0f06c110",
			2475 => x"040c7208",
			2476 => x"0e047804",
			2477 => x"feae2759",
			2478 => x"002f2759",
			2479 => x"0a02d104",
			2480 => x"04d62759",
			2481 => x"fed12759",
			2482 => x"02080908",
			2483 => x"0f06ca04",
			2484 => x"fe6b2759",
			2485 => x"fd112759",
			2486 => x"040c1204",
			2487 => x"00002759",
			2488 => x"fe4e2759",
			2489 => x"0208091c",
			2490 => x"06012b10",
			2491 => x"0e04d308",
			2492 => x"040a8804",
			2493 => x"005c2759",
			2494 => x"fdc72759",
			2495 => x"0a023304",
			2496 => x"fee62759",
			2497 => x"01082759",
			2498 => x"040bb208",
			2499 => x"00042804",
			2500 => x"00ff2759",
			2501 => x"fe8e2759",
			2502 => x"02c22759",
			2503 => x"08037910",
			2504 => x"09009508",
			2505 => x"0f071d04",
			2506 => x"01122759",
			2507 => x"fff62759",
			2508 => x"0e04f004",
			2509 => x"ff812759",
			2510 => x"fffa2759",
			2511 => x"00047508",
			2512 => x"06016704",
			2513 => x"03102759",
			2514 => x"00622759",
			2515 => x"01008004",
			2516 => x"00582759",
			2517 => x"fea42759",
			2518 => x"0c059cac",
			2519 => x"0304a738",
			2520 => x"0f06c534",
			2521 => x"07047a18",
			2522 => x"08031d08",
			2523 => x"03045e04",
			2524 => x"014728b5",
			2525 => x"045b28b5",
			2526 => x"07047908",
			2527 => x"0c047404",
			2528 => x"ff4f28b5",
			2529 => x"017a28b5",
			2530 => x"0c047304",
			2531 => x"02e828b5",
			2532 => x"fea528b5",
			2533 => x"03047710",
			2534 => x"0a02d108",
			2535 => x"06012904",
			2536 => x"001f28b5",
			2537 => x"fe9a28b5",
			2538 => x"0a02f304",
			2539 => x"00bc28b5",
			2540 => x"fec528b5",
			2541 => x"0b047004",
			2542 => x"02cb28b5",
			2543 => x"040c4c04",
			2544 => x"ff4f28b5",
			2545 => x"007428b5",
			2546 => x"fe0c28b5",
			2547 => x"0f07053c",
			2548 => x"0505101c",
			2549 => x"0a02ab10",
			2550 => x"0d052808",
			2551 => x"0b049d04",
			2552 => x"00d128b5",
			2553 => x"feac28b5",
			2554 => x"0304d804",
			2555 => x"015028b5",
			2556 => x"046d28b5",
			2557 => x"05050f08",
			2558 => x"0c047304",
			2559 => x"030028b5",
			2560 => x"003728b5",
			2561 => x"049428b5",
			2562 => x"0304d810",
			2563 => x"0f064a08",
			2564 => x"0d055a04",
			2565 => x"04e228b5",
			2566 => x"ff8428b5",
			2567 => x"01005904",
			2568 => x"ff7c28b5",
			2569 => x"022b28b5",
			2570 => x"0d058e08",
			2571 => x"03052504",
			2572 => x"004c28b5",
			2573 => x"00ff28b5",
			2574 => x"03056104",
			2575 => x"fed928b5",
			2576 => x"000128b5",
			2577 => x"03053318",
			2578 => x"03052f10",
			2579 => x"03052b08",
			2580 => x"0d054c04",
			2581 => x"ffda28b5",
			2582 => x"fe8a28b5",
			2583 => x"0c049104",
			2584 => x"024728b5",
			2585 => x"ffd028b5",
			2586 => x"0f071f04",
			2587 => x"febf28b5",
			2588 => x"fd9328b5",
			2589 => x"08038810",
			2590 => x"040c4408",
			2591 => x"08036904",
			2592 => x"000b28b5",
			2593 => x"00a928b5",
			2594 => x"0a02b104",
			2595 => x"ff0a28b5",
			2596 => x"001f28b5",
			2597 => x"0208c008",
			2598 => x"06015704",
			2599 => x"048528b5",
			2600 => x"007128b5",
			2601 => x"040cbf04",
			2602 => x"013f28b5",
			2603 => x"ffc628b5",
			2604 => x"fe7128b5",
			2605 => x"0f0773e4",
			2606 => x"0e04616c",
			2607 => x"0b049134",
			2608 => x"01004d1c",
			2609 => x"09007910",
			2610 => x"0c047408",
			2611 => x"07047d04",
			2612 => x"00252ba3",
			2613 => x"ff442ba3",
			2614 => x"07046404",
			2615 => x"fdf52ba3",
			2616 => x"00a92ba3",
			2617 => x"0b049008",
			2618 => x"0c047304",
			2619 => x"ffa72ba3",
			2620 => x"fe272ba3",
			2621 => x"01002ba3",
			2622 => x"0c04770c",
			2623 => x"09007d04",
			2624 => x"01462ba3",
			2625 => x"0304c704",
			2626 => x"fe212ba3",
			2627 => x"00142ba3",
			2628 => x"0704a808",
			2629 => x"0d053204",
			2630 => x"02c42ba3",
			2631 => x"00e92ba3",
			2632 => x"ff592ba3",
			2633 => x"06014918",
			2634 => x"0208c710",
			2635 => x"09007308",
			2636 => x"01004704",
			2637 => x"ff802ba3",
			2638 => x"034d2ba3",
			2639 => x"0e043604",
			2640 => x"fede2ba3",
			2641 => x"ffbe2ba3",
			2642 => x"0208d004",
			2643 => x"07b22ba3",
			2644 => x"00002ba3",
			2645 => x"0f06a510",
			2646 => x"0f066608",
			2647 => x"02081d04",
			2648 => x"fe532ba3",
			2649 => x"018f2ba3",
			2650 => x"0704c104",
			2651 => x"023a2ba3",
			2652 => x"fe912ba3",
			2653 => x"0d056608",
			2654 => x"05051e04",
			2655 => x"00e22ba3",
			2656 => x"fe6f2ba3",
			2657 => x"09008e04",
			2658 => x"02612ba3",
			2659 => x"fedd2ba3",
			2660 => x"0d054f3c",
			2661 => x"0b04af20",
			2662 => x"03053910",
			2663 => x"0f071708",
			2664 => x"0c049904",
			2665 => x"00342ba3",
			2666 => x"02132ba3",
			2667 => x"07049204",
			2668 => x"00672ba3",
			2669 => x"febb2ba3",
			2670 => x"040be408",
			2671 => x"0f074904",
			2672 => x"00c92ba3",
			2673 => x"fe472ba3",
			2674 => x"040c3804",
			2675 => x"03042ba3",
			2676 => x"01652ba3",
			2677 => x"0a029010",
			2678 => x"0a028308",
			2679 => x"07049104",
			2680 => x"027b2ba3",
			2681 => x"00872ba3",
			2682 => x"02086004",
			2683 => x"ff042ba3",
			2684 => x"01162ba3",
			2685 => x"0f06e304",
			2686 => x"030e2ba3",
			2687 => x"0e048804",
			2688 => x"ff8a2ba3",
			2689 => x"017c2ba3",
			2690 => x"0e051620",
			2691 => x"0900a810",
			2692 => x"01005c08",
			2693 => x"09009304",
			2694 => x"001d2ba3",
			2695 => x"ff152ba3",
			2696 => x"0c04d104",
			2697 => x"00312ba3",
			2698 => x"02822ba3",
			2699 => x"040ba408",
			2700 => x"03056104",
			2701 => x"feb72ba3",
			2702 => x"00bd2ba3",
			2703 => x"06015704",
			2704 => x"fe7b2ba3",
			2705 => x"ffeb2ba3",
			2706 => x"0900ba10",
			2707 => x"0c049208",
			2708 => x"0c048f04",
			2709 => x"00782ba3",
			2710 => x"fea72ba3",
			2711 => x"0b04d004",
			2712 => x"01822ba3",
			2713 => x"009b2ba3",
			2714 => x"0a02b008",
			2715 => x"01007b04",
			2716 => x"ffb22ba3",
			2717 => x"00c32ba3",
			2718 => x"fdf32ba3",
			2719 => x"0704da5c",
			2720 => x"0a02b42c",
			2721 => x"040bde18",
			2722 => x"0c04cb0c",
			2723 => x"06013504",
			2724 => x"fde62ba3",
			2725 => x"0208c204",
			2726 => x"00592ba3",
			2727 => x"ff592ba3",
			2728 => x"0d05de08",
			2729 => x"0a029504",
			2730 => x"fd392ba3",
			2731 => x"ff192ba3",
			2732 => x"00e42ba3",
			2733 => x"0d053308",
			2734 => x"07047c04",
			2735 => x"fec02ba3",
			2736 => x"02672ba3",
			2737 => x"02089f04",
			2738 => x"00d62ba3",
			2739 => x"0c04d104",
			2740 => x"fedc2ba3",
			2741 => x"008a2ba3",
			2742 => x"0b050220",
			2743 => x"040c8510",
			2744 => x"05058208",
			2745 => x"0208e204",
			2746 => x"01712ba3",
			2747 => x"ff592ba3",
			2748 => x"06015b04",
			2749 => x"03022ba3",
			2750 => x"01932ba3",
			2751 => x"0704c008",
			2752 => x"0e04f004",
			2753 => x"fe552ba3",
			2754 => x"00af2ba3",
			2755 => x"0c049204",
			2756 => x"00002ba3",
			2757 => x"fe472ba3",
			2758 => x"0c04b104",
			2759 => x"01822ba3",
			2760 => x"0e055a04",
			2761 => x"ff452ba3",
			2762 => x"0505af04",
			2763 => x"fd672ba3",
			2764 => x"feb62ba3",
			2765 => x"0704eb1c",
			2766 => x"0f078104",
			2767 => x"fea42ba3",
			2768 => x"0100730c",
			2769 => x"0b04f004",
			2770 => x"00482ba3",
			2771 => x"01006c04",
			2772 => x"01a02ba3",
			2773 => x"02d22ba3",
			2774 => x"06016008",
			2775 => x"040b5d04",
			2776 => x"01082ba3",
			2777 => x"ff8e2ba3",
			2778 => x"01d72ba3",
			2779 => x"03059904",
			2780 => x"02832ba3",
			2781 => x"0900a708",
			2782 => x"0f079604",
			2783 => x"fead2ba3",
			2784 => x"fce62ba3",
			2785 => x"0c04b408",
			2786 => x"06015604",
			2787 => x"002b2ba3",
			2788 => x"fed92ba3",
			2789 => x"02084504",
			2790 => x"fe3d2ba3",
			2791 => x"00182ba3",
			2792 => x"05061674",
			2793 => x"07051c58",
			2794 => x"07051a3c",
			2795 => x"0704aa20",
			2796 => x"07049710",
			2797 => x"07049308",
			2798 => x"01006204",
			2799 => x"00142d15",
			2800 => x"01da2d15",
			2801 => x"0b049104",
			2802 => x"feaa2d15",
			2803 => x"ffbe2d15",
			2804 => x"05051408",
			2805 => x"0704a704",
			2806 => x"02332d15",
			2807 => x"00cc2d15",
			2808 => x"02090c04",
			2809 => x"003c2d15",
			2810 => x"02f92d15",
			2811 => x"0704ab0c",
			2812 => x"06012404",
			2813 => x"018c2d15",
			2814 => x"05056604",
			2815 => x"fe9f2d15",
			2816 => x"fff32d15",
			2817 => x"0a024708",
			2818 => x"02083304",
			2819 => x"ff862d15",
			2820 => x"fdcb2d15",
			2821 => x"0704be04",
			2822 => x"00442d15",
			2823 => x"fff92d15",
			2824 => x"0e05d80c",
			2825 => x"07051b08",
			2826 => x"08035004",
			2827 => x"016d2d15",
			2828 => x"04462d15",
			2829 => x"ff152d15",
			2830 => x"06015e04",
			2831 => x"fed32d15",
			2832 => x"0c04ea08",
			2833 => x"0b055404",
			2834 => x"feab2d15",
			2835 => x"008e2d15",
			2836 => x"02622d15",
			2837 => x"0a028b10",
			2838 => x"0c04ee04",
			2839 => x"fe2a2d15",
			2840 => x"0c050908",
			2841 => x"0a015104",
			2842 => x"00002d15",
			2843 => x"02c72d15",
			2844 => x"feff2d15",
			2845 => x"0f082b04",
			2846 => x"fe382d15",
			2847 => x"0306b904",
			2848 => x"009b2d15",
			2849 => x"fe732d15",
			2850 => x"0e07582c",
			2851 => x"0a02bf28",
			2852 => x"08035218",
			2853 => x"05066c0c",
			2854 => x"02092408",
			2855 => x"0a029e04",
			2856 => x"01382d15",
			2857 => x"fe872d15",
			2858 => x"fe572d15",
			2859 => x"05069808",
			2860 => x"0207ed04",
			2861 => x"00002d15",
			2862 => x"02862d15",
			2863 => x"00002d15",
			2864 => x"02094304",
			2865 => x"013d2d15",
			2866 => x"0f08bf08",
			2867 => x"07056104",
			2868 => x"03d72d15",
			2869 => x"00002d15",
			2870 => x"00002d15",
			2871 => x"fe9d2d15",
			2872 => x"0100b408",
			2873 => x"0208dd04",
			2874 => x"00842d15",
			2875 => x"fe562d15",
			2876 => x"0c05b810",
			2877 => x"0601800c",
			2878 => x"02091304",
			2879 => x"ff6d2d15",
			2880 => x"0c052704",
			2881 => x"020b2d15",
			2882 => x"006d2d15",
			2883 => x"feea2d15",
			2884 => x"fe9d2d15",
			2885 => x"07051b78",
			2886 => x"01002a08",
			2887 => x"06013904",
			2888 => x"fe4c2e79",
			2889 => x"012b2e79",
			2890 => x"08037140",
			2891 => x"06013d20",
			2892 => x"02087e10",
			2893 => x"0304d808",
			2894 => x"0b048104",
			2895 => x"01912e79",
			2896 => x"fff32e79",
			2897 => x"0a024504",
			2898 => x"00222e79",
			2899 => x"01ce2e79",
			2900 => x"08034f08",
			2901 => x"03056804",
			2902 => x"fe1c2e79",
			2903 => x"ff282e79",
			2904 => x"07049504",
			2905 => x"022e2e79",
			2906 => x"feaa2e79",
			2907 => x"0208f210",
			2908 => x"08035608",
			2909 => x"0c04d004",
			2910 => x"028a2e79",
			2911 => x"01732e79",
			2912 => x"0a029b04",
			2913 => x"ffe52e79",
			2914 => x"01d82e79",
			2915 => x"0e05a408",
			2916 => x"02090004",
			2917 => x"ff2a2e79",
			2918 => x"fddd2e79",
			2919 => x"0505df04",
			2920 => x"01a52e79",
			2921 => x"ff122e79",
			2922 => x"07047a14",
			2923 => x"0207d108",
			2924 => x"0b046d04",
			2925 => x"01652e79",
			2926 => x"ff692e79",
			2927 => x"01004b08",
			2928 => x"08038504",
			2929 => x"01c52e79",
			2930 => x"04d32e79",
			2931 => x"008b2e79",
			2932 => x"0803a310",
			2933 => x"03048f08",
			2934 => x"06014a04",
			2935 => x"fecd2e79",
			2936 => x"018b2e79",
			2937 => x"0704be04",
			2938 => x"01562e79",
			2939 => x"00592e79",
			2940 => x"06014104",
			2941 => x"02ce2e79",
			2942 => x"01005304",
			2943 => x"ffbe2e79",
			2944 => x"feae2e79",
			2945 => x"0c052a2c",
			2946 => x"03065910",
			2947 => x"03063a04",
			2948 => x"fe3c2e79",
			2949 => x"02089808",
			2950 => x"05063504",
			2951 => x"011f2e79",
			2952 => x"fe9e2e79",
			2953 => x"fe3d2e79",
			2954 => x"06017010",
			2955 => x"06013104",
			2956 => x"fe602e79",
			2957 => x"0f07dc04",
			2958 => x"04652e79",
			2959 => x"02091904",
			2960 => x"ffbb2e79",
			2961 => x"021c2e79",
			2962 => x"0d069f04",
			2963 => x"fe412e79",
			2964 => x"0209b104",
			2965 => x"05a22e79",
			2966 => x"fe5e2e79",
			2967 => x"0705730c",
			2968 => x"07056104",
			2969 => x"fe5d2e79",
			2970 => x"0c054804",
			2971 => x"01962e79",
			2972 => x"feda2e79",
			2973 => x"fe4d2e79",
			2974 => x"0c050b6c",
			2975 => x"040fc668",
			2976 => x"07050340",
			2977 => x"0e051620",
			2978 => x"0900a910",
			2979 => x"02087e08",
			2980 => x"0e048804",
			2981 => x"00682fa5",
			2982 => x"00eb2fa5",
			2983 => x"0a029e04",
			2984 => x"ff6f2fa5",
			2985 => x"006d2fa5",
			2986 => x"040ba408",
			2987 => x"03056104",
			2988 => x"fea62fa5",
			2989 => x"00ab2fa5",
			2990 => x"08034404",
			2991 => x"fd2a2fa5",
			2992 => x"ff522fa5",
			2993 => x"0900b510",
			2994 => x"040c9308",
			2995 => x"0a02c304",
			2996 => x"01302fa5",
			2997 => x"040a2fa5",
			2998 => x"0e056804",
			2999 => x"fea82fa5",
			3000 => x"00d92fa5",
			3001 => x"0e054b08",
			3002 => x"02086e04",
			3003 => x"00412fa5",
			3004 => x"fe912fa5",
			3005 => x"040bbf04",
			3006 => x"010b2fa5",
			3007 => x"003c2fa5",
			3008 => x"06017d20",
			3009 => x"02093d10",
			3010 => x"0a02b608",
			3011 => x"06012b04",
			3012 => x"fe3a2fa5",
			3013 => x"002a2fa5",
			3014 => x"0900bc04",
			3015 => x"006e2fa5",
			3016 => x"fe5b2fa5",
			3017 => x"00045b08",
			3018 => x"07051a04",
			3019 => x"fe112fa5",
			3020 => x"01992fa5",
			3021 => x"0b054304",
			3022 => x"04472fa5",
			3023 => x"00df2fa5",
			3024 => x"0b05a704",
			3025 => x"fe5b2fa5",
			3026 => x"00932fa5",
			3027 => x"fe602fa5",
			3028 => x"0c054818",
			3029 => x"0b061b14",
			3030 => x"0900dc04",
			3031 => x"fe382fa5",
			3032 => x"0900e004",
			3033 => x"02d12fa5",
			3034 => x"0b05b608",
			3035 => x"0d069f04",
			3036 => x"fef12fa5",
			3037 => x"02322fa5",
			3038 => x"fe592fa5",
			3039 => x"01d32fa5",
			3040 => x"0c05b810",
			3041 => x"0802c70c",
			3042 => x"0802bb04",
			3043 => x"fe702fa5",
			3044 => x"0c059f04",
			3045 => x"00c22fa5",
			3046 => x"030f2fa5",
			3047 => x"fe612fa5",
			3048 => x"fe5f2fa5",
			3049 => x"0c050b78",
			3050 => x"040fc674",
			3051 => x"0900cd3c",
			3052 => x"06015720",
			3053 => x"0f07a610",
			3054 => x"0e054b08",
			3055 => x"0900b504",
			3056 => x"007c3101",
			3057 => x"ff433101",
			3058 => x"0b051104",
			3059 => x"01543101",
			3060 => x"000d3101",
			3061 => x"06014a08",
			3062 => x"0f07d504",
			3063 => x"ff493101",
			3064 => x"fdbf3101",
			3065 => x"040bc404",
			3066 => x"016f3101",
			3067 => x"fff83101",
			3068 => x"0004a010",
			3069 => x"0900ab08",
			3070 => x"040c9304",
			3071 => x"02f33101",
			3072 => x"ff533101",
			3073 => x"0305f204",
			3074 => x"00883101",
			3075 => x"01c63101",
			3076 => x"06015a04",
			3077 => x"034e3101",
			3078 => x"0e057f04",
			3079 => x"fed33101",
			3080 => x"01403101",
			3081 => x"0e05ce1c",
			3082 => x"00042810",
			3083 => x"0f074608",
			3084 => x"0b054304",
			3085 => x"fcf33101",
			3086 => x"fe5a3101",
			3087 => x"0b052404",
			3088 => x"00003101",
			3089 => x"02c43101",
			3090 => x"03063a08",
			3091 => x"07051804",
			3092 => x"fd5b3101",
			3093 => x"fef93101",
			3094 => x"ffe83101",
			3095 => x"0c04af0c",
			3096 => x"040adc04",
			3097 => x"00ab3101",
			3098 => x"0b052004",
			3099 => x"fc8f3101",
			3100 => x"fee33101",
			3101 => x"0704ec08",
			3102 => x"0900e404",
			3103 => x"02513101",
			3104 => x"ff213101",
			3105 => x"0409ed04",
			3106 => x"01d43101",
			3107 => x"00043101",
			3108 => x"fe633101",
			3109 => x"0c054824",
			3110 => x"09010f10",
			3111 => x"07052f04",
			3112 => x"fe373101",
			3113 => x"07053104",
			3114 => x"012d3101",
			3115 => x"0b055404",
			3116 => x"00253101",
			3117 => x"fe5f3101",
			3118 => x"00038508",
			3119 => x"0f07e304",
			3120 => x"fef03101",
			3121 => x"025f3101",
			3122 => x"09012008",
			3123 => x"09011b04",
			3124 => x"ff423101",
			3125 => x"02373101",
			3126 => x"fe5d3101",
			3127 => x"0c05b810",
			3128 => x"0802c70c",
			3129 => x"0802bb04",
			3130 => x"fe7a3101",
			3131 => x"0c059f04",
			3132 => x"009e3101",
			3133 => x"02543101",
			3134 => x"fe643101",
			3135 => x"fe613101",
			3136 => x"0c04f178",
			3137 => x"09004204",
			3138 => x"fe503265",
			3139 => x"0e04bb38",
			3140 => x"0704c11c",
			3141 => x"0e04260c",
			3142 => x"0802d404",
			3143 => x"04693265",
			3144 => x"09006204",
			3145 => x"01763265",
			3146 => x"00113265",
			3147 => x"0f070508",
			3148 => x"0802d204",
			3149 => x"fe3b3265",
			3150 => x"01873265",
			3151 => x"0d054d04",
			3152 => x"00db3265",
			3153 => x"ff6b3265",
			3154 => x"03051b10",
			3155 => x"09008f08",
			3156 => x"0304c704",
			3157 => x"fe3b3265",
			3158 => x"00393265",
			3159 => x"0a026904",
			3160 => x"ff723265",
			3161 => x"fe213265",
			3162 => x"09008c04",
			3163 => x"036c3265",
			3164 => x"0f06b204",
			3165 => x"02403265",
			3166 => x"ffbb3265",
			3167 => x"02087e20",
			3168 => x"06012910",
			3169 => x"0b04d308",
			3170 => x"0d055c04",
			3171 => x"00033265",
			3172 => x"02ff3265",
			3173 => x"06012404",
			3174 => x"fe4b3265",
			3175 => x"ffa73265",
			3176 => x"0900a908",
			3177 => x"0f070504",
			3178 => x"03383265",
			3179 => x"02433265",
			3180 => x"08036304",
			3181 => x"01fd3265",
			3182 => x"fe1f3265",
			3183 => x"0306c510",
			3184 => x"0e054b08",
			3185 => x"0b04c004",
			3186 => x"018c3265",
			3187 => x"00283265",
			3188 => x"0704d504",
			3189 => x"02493265",
			3190 => x"012c3265",
			3191 => x"05065108",
			3192 => x"0d061f04",
			3193 => x"00483265",
			3194 => x"fe973265",
			3195 => x"015b3265",
			3196 => x"0c052a2c",
			3197 => x"0f07ce10",
			3198 => x"07050604",
			3199 => x"00003265",
			3200 => x"0f07a304",
			3201 => x"fe4a3265",
			3202 => x"0f07b204",
			3203 => x"00003265",
			3204 => x"fe403265",
			3205 => x"02099514",
			3206 => x"0d06ab0c",
			3207 => x"01009f08",
			3208 => x"0d065104",
			3209 => x"00213265",
			3210 => x"02663265",
			3211 => x"fe383265",
			3212 => x"0307b004",
			3213 => x"03a43265",
			3214 => x"00e63265",
			3215 => x"0a029b04",
			3216 => x"00d23265",
			3217 => x"fe5a3265",
			3218 => x"0705730c",
			3219 => x"07056104",
			3220 => x"fe613265",
			3221 => x"0c054804",
			3222 => x"015e3265",
			3223 => x"feef3265",
			3224 => x"fe523265",
			3225 => x"0c054378",
			3226 => x"040fc674",
			3227 => x"0208093c",
			3228 => x"0601251c",
			3229 => x"05053110",
			3230 => x"0304e708",
			3231 => x"0802fc04",
			3232 => x"01b93389",
			3233 => x"ff573389",
			3234 => x"07049304",
			3235 => x"00203389",
			3236 => x"03fb3389",
			3237 => x"0f069004",
			3238 => x"fe423389",
			3239 => x"0900b904",
			3240 => x"ff7a3389",
			3241 => x"02fa3389",
			3242 => x"0d052610",
			3243 => x"040c0408",
			3244 => x"08033004",
			3245 => x"005c3389",
			3246 => x"fef13389",
			3247 => x"0a029204",
			3248 => x"03273389",
			3249 => x"00373389",
			3250 => x"0a027d08",
			3251 => x"03051b04",
			3252 => x"ffeb3389",
			3253 => x"00ef3389",
			3254 => x"06013a04",
			3255 => x"02183389",
			3256 => x"00d33389",
			3257 => x"0a02bb1c",
			3258 => x"02080e0c",
			3259 => x"040b1604",
			3260 => x"fd4f3389",
			3261 => x"040b6b04",
			3262 => x"01c23389",
			3263 => x"fe8d3389",
			3264 => x"040c2c08",
			3265 => x"0a029304",
			3266 => x"00133389",
			3267 => x"00913389",
			3268 => x"01004104",
			3269 => x"014f3389",
			3270 => x"ffd33389",
			3271 => x"0f06990c",
			3272 => x"02081504",
			3273 => x"00003389",
			3274 => x"03048704",
			3275 => x"01353389",
			3276 => x"04a43389",
			3277 => x"0803a308",
			3278 => x"040d5504",
			3279 => x"00ad3389",
			3280 => x"03c23389",
			3281 => x"02086004",
			3282 => x"fe2f3389",
			3283 => x"ffa93389",
			3284 => x"fe6b3389",
			3285 => x"0c05b818",
			3286 => x"030a1210",
			3287 => x"0705730c",
			3288 => x"06016b04",
			3289 => x"fea83389",
			3290 => x"06017304",
			3291 => x"014e3389",
			3292 => x"fff23389",
			3293 => x"fe6c3389",
			3294 => x"040b9f04",
			3295 => x"03013389",
			3296 => x"00003389",
			3297 => x"fe663389",
			3298 => x"07053180",
			3299 => x"09004f08",
			3300 => x"06013e04",
			3301 => x"fe54350d",
			3302 => x"0154350d",
			3303 => x"040c2640",
			3304 => x"06013a20",
			3305 => x"02084d10",
			3306 => x"0f067408",
			3307 => x"0b04af04",
			3308 => x"00ab350d",
			3309 => x"fee2350d",
			3310 => x"03051004",
			3311 => x"00a5350d",
			3312 => x"0174350d",
			3313 => x"0003ed08",
			3314 => x"040abb04",
			3315 => x"0000350d",
			3316 => x"fdf6350d",
			3317 => x"03057904",
			3318 => x"ffab350d",
			3319 => x"0176350d",
			3320 => x"0b053110",
			3321 => x"040b9708",
			3322 => x"0a029304",
			3323 => x"020c350d",
			3324 => x"02e5350d",
			3325 => x"0a028a04",
			3326 => x"fff6350d",
			3327 => x"01ae350d",
			3328 => x"06016208",
			3329 => x"040a7b04",
			3330 => x"033a350d",
			3331 => x"00b1350d",
			3332 => x"0900fb04",
			3333 => x"ffe8350d",
			3334 => x"fea5350d",
			3335 => x"09008d1c",
			3336 => x"0207b510",
			3337 => x"06013508",
			3338 => x"06012d04",
			3339 => x"fe58350d",
			3340 => x"0564350d",
			3341 => x"07049104",
			3342 => x"fe31350d",
			3343 => x"ff84350d",
			3344 => x"0a028304",
			3345 => x"fe58350d",
			3346 => x"0c045404",
			3347 => x"042f350d",
			3348 => x"0113350d",
			3349 => x"0e04a50c",
			3350 => x"08038d08",
			3351 => x"0f06f304",
			3352 => x"0057350d",
			3353 => x"feb6350d",
			3354 => x"fe3a350d",
			3355 => x"040c9308",
			3356 => x"08037404",
			3357 => x"0000350d",
			3358 => x"018c350d",
			3359 => x"0704a704",
			3360 => x"01e0350d",
			3361 => x"ff94350d",
			3362 => x"0c05452c",
			3363 => x"0d069f18",
			3364 => x"0e061e04",
			3365 => x"fe4e350d",
			3366 => x"040b4a0c",
			3367 => x"0f07f208",
			3368 => x"0e064304",
			3369 => x"feba350d",
			3370 => x"0097350d",
			3371 => x"fe21350d",
			3372 => x"0c050a04",
			3373 => x"02bd350d",
			3374 => x"fe69350d",
			3375 => x"040c0c10",
			3376 => x"06017c08",
			3377 => x"00032c04",
			3378 => x"fe6e350d",
			3379 => x"0423350d",
			3380 => x"08035a04",
			3381 => x"fe63350d",
			3382 => x"00ce350d",
			3383 => x"fe55350d",
			3384 => x"0c05b814",
			3385 => x"07063d10",
			3386 => x"0705730c",
			3387 => x"07056104",
			3388 => x"fe78350d",
			3389 => x"0c054c04",
			3390 => x"00d2350d",
			3391 => x"fef1350d",
			3392 => x"fe5a350d",
			3393 => x"075a350d",
			3394 => x"fe52350d",
			3395 => x"0803a398",
			3396 => x"0a02d178",
			3397 => x"0a02933c",
			3398 => x"08034d20",
			3399 => x"09008c10",
			3400 => x"07047c08",
			3401 => x"08033f04",
			3402 => x"ffb836d9",
			3403 => x"fdb736d9",
			3404 => x"040bff04",
			3405 => x"002c36d9",
			3406 => x"014d36d9",
			3407 => x"09008e08",
			3408 => x"06013004",
			3409 => x"fdfb36d9",
			3410 => x"ff5c36d9",
			3411 => x"09008f04",
			3412 => x"00bc36d9",
			3413 => x"ffe636d9",
			3414 => x"040c2c10",
			3415 => x"0a029208",
			3416 => x"0c047804",
			3417 => x"fe9e36d9",
			3418 => x"003036d9",
			3419 => x"07049204",
			3420 => x"ff5736d9",
			3421 => x"fdf436d9",
			3422 => x"08035204",
			3423 => x"fe2d36d9",
			3424 => x"06013104",
			3425 => x"fea736d9",
			3426 => x"021136d9",
			3427 => x"040bf720",
			3428 => x"0d05b510",
			3429 => x"06013e08",
			3430 => x"09008d04",
			3431 => x"ffe036d9",
			3432 => x"fdf036d9",
			3433 => x"0f071f04",
			3434 => x"017636d9",
			3435 => x"009336d9",
			3436 => x"0f07ce08",
			3437 => x"0d05c204",
			3438 => x"fe6636d9",
			3439 => x"ffd336d9",
			3440 => x"0e05ac04",
			3441 => x"020836d9",
			3442 => x"004436d9",
			3443 => x"0c04760c",
			3444 => x"0f07a308",
			3445 => x"0c047404",
			3446 => x"001736d9",
			3447 => x"00e836d9",
			3448 => x"022d36d9",
			3449 => x"00045308",
			3450 => x"09009904",
			3451 => x"012236d9",
			3452 => x"fef536d9",
			3453 => x"0d05b604",
			3454 => x"ffd936d9",
			3455 => x"006936d9",
			3456 => x"09008e04",
			3457 => x"023d36d9",
			3458 => x"0b04e208",
			3459 => x"0e050d04",
			3460 => x"fe7236d9",
			3461 => x"ffb836d9",
			3462 => x"0900ba08",
			3463 => x"0e051d04",
			3464 => x"000036d9",
			3465 => x"024936d9",
			3466 => x"0f082b04",
			3467 => x"fe8336d9",
			3468 => x"01008604",
			3469 => x"01c336d9",
			3470 => x"fe8736d9",
			3471 => x"0c04751c",
			3472 => x"0004dd04",
			3473 => x"fea036d9",
			3474 => x"0b048e10",
			3475 => x"09005d0c",
			3476 => x"0f059f04",
			3477 => x"ff3436d9",
			3478 => x"0c045c04",
			3479 => x"015036d9",
			3480 => x"000036d9",
			3481 => x"fee236d9",
			3482 => x"0d050f04",
			3483 => x"ff5d36d9",
			3484 => x"02eb36d9",
			3485 => x"0704a814",
			3486 => x"040e6308",
			3487 => x"0d050004",
			3488 => x"ff4a36d9",
			3489 => x"fe2e36d9",
			3490 => x"06014608",
			3491 => x"00057a04",
			3492 => x"013636d9",
			3493 => x"000036d9",
			3494 => x"ff5836d9",
			3495 => x"01005410",
			3496 => x"0a02d704",
			3497 => x"fe8036d9",
			3498 => x"0a02e404",
			3499 => x"019c36d9",
			3500 => x"09007504",
			3501 => x"fecd36d9",
			3502 => x"005736d9",
			3503 => x"0004ab04",
			3504 => x"010336d9",
			3505 => x"0b04bf04",
			3506 => x"000336d9",
			3507 => x"040ca004",
			3508 => x"000036d9",
			3509 => x"fe5d36d9",
			3510 => x"0c05457c",
			3511 => x"040fc678",
			3512 => x"0c04b240",
			3513 => x"0c049620",
			3514 => x"0c049510",
			3515 => x"0704a708",
			3516 => x"0b04d004",
			3517 => x"00ac381d",
			3518 => x"0263381d",
			3519 => x"0704ad04",
			3520 => x"ffc6381d",
			3521 => x"0098381d",
			3522 => x"0704bf08",
			3523 => x"0704bc04",
			3524 => x"ff4c381d",
			3525 => x"0239381d",
			3526 => x"0704c404",
			3527 => x"fe24381d",
			3528 => x"ffba381d",
			3529 => x"0c049710",
			3530 => x"0704be08",
			3531 => x"0704ab04",
			3532 => x"01f0381d",
			3533 => x"ff72381d",
			3534 => x"0b04bf04",
			3535 => x"03c3381d",
			3536 => x"01ef381d",
			3537 => x"040c7208",
			3538 => x"0c049804",
			3539 => x"fee4381d",
			3540 => x"00d5381d",
			3541 => x"01004f04",
			3542 => x"0127381d",
			3543 => x"fed4381d",
			3544 => x"0c04b318",
			3545 => x"0d05b610",
			3546 => x"06014d08",
			3547 => x"02086c04",
			3548 => x"ff2c381d",
			3549 => x"fd6b381d",
			3550 => x"0e054b04",
			3551 => x"feff381d",
			3552 => x"0186381d",
			3553 => x"0d05cf04",
			3554 => x"fcf2381d",
			3555 => x"fe2d381d",
			3556 => x"06014210",
			3557 => x"040b4208",
			3558 => x"0a026504",
			3559 => x"ffa9381d",
			3560 => x"018f381d",
			3561 => x"0e053404",
			3562 => x"ff39381d",
			3563 => x"fd7f381d",
			3564 => x"0a028a08",
			3565 => x"040b9704",
			3566 => x"0117381d",
			3567 => x"ff20381d",
			3568 => x"0900c804",
			3569 => x"0072381d",
			3570 => x"ff92381d",
			3571 => x"fe64381d",
			3572 => x"0c05b824",
			3573 => x"07061318",
			3574 => x"0705fc10",
			3575 => x"0705730c",
			3576 => x"07056104",
			3577 => x"fec2381d",
			3578 => x"0c054c04",
			3579 => x"005a381d",
			3580 => x"fff7381d",
			3581 => x"fe66381d",
			3582 => x"0c059b04",
			3583 => x"0333381d",
			3584 => x"fe9e381d",
			3585 => x"040a8804",
			3586 => x"fee5381d",
			3587 => x"0a029504",
			3588 => x"03d3381d",
			3589 => x"ffeb381d",
			3590 => x"fe62381d",
			3591 => x"0c0548ac",
			3592 => x"0a027868",
			3593 => x"040b362c",
			3594 => x"040b3020",
			3595 => x"040acf10",
			3596 => x"08031708",
			3597 => x"0a023904",
			3598 => x"ffd43991",
			3599 => x"00ba3991",
			3600 => x"02081d04",
			3601 => x"00563991",
			3602 => x"fbf33991",
			3603 => x"0003e108",
			3604 => x"01006504",
			3605 => x"fffa3991",
			3606 => x"fdfa3991",
			3607 => x"0e04f904",
			3608 => x"ffd03991",
			3609 => x"00bf3991",
			3610 => x"0900a008",
			3611 => x"0b04ae04",
			3612 => x"03023991",
			3613 => x"fe843991",
			3614 => x"02a83991",
			3615 => x"0f06d91c",
			3616 => x"0100500c",
			3617 => x"0e046b08",
			3618 => x"0704aa04",
			3619 => x"00d03991",
			3620 => x"fe4e3991",
			3621 => x"03733991",
			3622 => x"0c049608",
			3623 => x"0f06c504",
			3624 => x"ffd83991",
			3625 => x"fe0e3991",
			3626 => x"08032104",
			3627 => x"004b3991",
			3628 => x"03253991",
			3629 => x"0d055a10",
			3630 => x"0b049008",
			3631 => x"00042004",
			3632 => x"fe443991",
			3633 => x"01b73991",
			3634 => x"0e04a904",
			3635 => x"fdb93991",
			3636 => x"fe973991",
			3637 => x"0c04ad08",
			3638 => x"0e055204",
			3639 => x"000e3991",
			3640 => x"fdb33991",
			3641 => x"0c04b404",
			3642 => x"fe093991",
			3643 => x"ffbb3991",
			3644 => x"0003ed14",
			3645 => x"0d05f704",
			3646 => x"fbba3991",
			3647 => x"0208c704",
			3648 => x"01bf3991",
			3649 => x"08031b08",
			3650 => x"08031804",
			3651 => x"fe583991",
			3652 => x"00b33991",
			3653 => x"fe3d3991",
			3654 => x"040b9f10",
			3655 => x"0004540c",
			3656 => x"01004904",
			3657 => x"fe2b3991",
			3658 => x"0c045c04",
			3659 => x"fed73991",
			3660 => x"00b33991",
			3661 => x"fdb43991",
			3662 => x"0704be10",
			3663 => x"0704ad08",
			3664 => x"0704aa04",
			3665 => x"00603991",
			3666 => x"ff593991",
			3667 => x"0f06d904",
			3668 => x"026c3991",
			3669 => x"00a93991",
			3670 => x"08034508",
			3671 => x"0f075d04",
			3672 => x"ff4a3991",
			3673 => x"fe523991",
			3674 => x"0704c204",
			3675 => x"ff9f3991",
			3676 => x"00493991",
			3677 => x"0c05b80c",
			3678 => x"00036308",
			3679 => x"00035304",
			3680 => x"feb13991",
			3681 => x"028c3991",
			3682 => x"fe743991",
			3683 => x"fe673991",
			3684 => x"0304d880",
			3685 => x"040c8c38",
			3686 => x"00048a28",
			3687 => x"0304cf18",
			3688 => x"02082410",
			3689 => x"0f06ac08",
			3690 => x"08036904",
			3691 => x"ff983b85",
			3692 => x"008f3b85",
			3693 => x"05050204",
			3694 => x"fee43b85",
			3695 => x"01bd3b85",
			3696 => x"0d050204",
			3697 => x"00f03b85",
			3698 => x"fe173b85",
			3699 => x"07047c04",
			3700 => x"00613b85",
			3701 => x"0f06ac08",
			3702 => x"0d053504",
			3703 => x"00813b85",
			3704 => x"fea83b85",
			3705 => x"fe173b85",
			3706 => x"06014504",
			3707 => x"fe383b85",
			3708 => x"0d051b04",
			3709 => x"01453b85",
			3710 => x"0d054e04",
			3711 => x"fe8e3b85",
			3712 => x"00003b85",
			3713 => x"040ca714",
			3714 => x"01005110",
			3715 => x"0a02bc0c",
			3716 => x"08037c08",
			3717 => x"06013904",
			3718 => x"02aa3b85",
			3719 => x"00ef3b85",
			3720 => x"ff213b85",
			3721 => x"02863b85",
			3722 => x"fe8a3b85",
			3723 => x"01003f1c",
			3724 => x"0f05ee10",
			3725 => x"0d04d908",
			3726 => x"0c045b04",
			3727 => x"fff13b85",
			3728 => x"00d73b85",
			3729 => x"0207ed04",
			3730 => x"fe6b3b85",
			3731 => x"00003b85",
			3732 => x"0c049208",
			3733 => x"0f06b504",
			3734 => x"01a83b85",
			3735 => x"00003b85",
			3736 => x"fec23b85",
			3737 => x"0207ed0c",
			3738 => x"03047708",
			3739 => x"0a02d704",
			3740 => x"fe833b85",
			3741 => x"00db3b85",
			3742 => x"02893b85",
			3743 => x"09008c08",
			3744 => x"040d5504",
			3745 => x"ff173b85",
			3746 => x"00223b85",
			3747 => x"02033b85",
			3748 => x"09007714",
			3749 => x"06012d04",
			3750 => x"fe3e3b85",
			3751 => x"06013904",
			3752 => x"027c3b85",
			3753 => x"06014104",
			3754 => x"00003b85",
			3755 => x"0304fe04",
			3756 => x"000a3b85",
			3757 => x"02273b85",
			3758 => x"0f06c12c",
			3759 => x"09008810",
			3760 => x"0100530c",
			3761 => x"05053c08",
			3762 => x"0704a804",
			3763 => x"005f3b85",
			3764 => x"01eb3b85",
			3765 => x"febf3b85",
			3766 => x"02a53b85",
			3767 => x"0d056710",
			3768 => x"0f06bb08",
			3769 => x"08031e04",
			3770 => x"fea13b85",
			3771 => x"00003b85",
			3772 => x"03050d04",
			3773 => x"01d43b85",
			3774 => x"00553b85",
			3775 => x"0c047e04",
			3776 => x"fea73b85",
			3777 => x"0d057504",
			3778 => x"01873b85",
			3779 => x"00333b85",
			3780 => x"06013520",
			3781 => x"03056810",
			3782 => x"05055508",
			3783 => x"040baa04",
			3784 => x"005a3b85",
			3785 => x"ff103b85",
			3786 => x"040ac904",
			3787 => x"001e3b85",
			3788 => x"fe6c3b85",
			3789 => x"0305b008",
			3790 => x"0c04ce04",
			3791 => x"00f33b85",
			3792 => x"fe2a3b85",
			3793 => x"01008604",
			3794 => x"fed83b85",
			3795 => x"00933b85",
			3796 => x"0207e50c",
			3797 => x"05056704",
			3798 => x"fd423b85",
			3799 => x"08030204",
			3800 => x"fe583b85",
			3801 => x"00a83b85",
			3802 => x"0d053508",
			3803 => x"02081b04",
			3804 => x"02853b85",
			3805 => x"00563b85",
			3806 => x"03051004",
			3807 => x"ff823b85",
			3808 => x"00153b85",
			3809 => x"0208d694",
			3810 => x"040d5554",
			3811 => x"0004b834",
			3812 => x"0504e714",
			3813 => x"0504e510",
			3814 => x"02081108",
			3815 => x"06013104",
			3816 => x"00aa3dc1",
			3817 => x"fe8e3dc1",
			3818 => x"03048f04",
			3819 => x"01113dc1",
			3820 => x"02de3dc1",
			3821 => x"031a3dc1",
			3822 => x"0b048010",
			3823 => x"040c3808",
			3824 => x"0d051904",
			3825 => x"fe743dc1",
			3826 => x"00003dc1",
			3827 => x"07047e04",
			3828 => x"00ef3dc1",
			3829 => x"febd3dc1",
			3830 => x"09007908",
			3831 => x"0304c004",
			3832 => x"002f3dc1",
			3833 => x"014a3dc1",
			3834 => x"06014104",
			3835 => x"ffee3dc1",
			3836 => x"002b3dc1",
			3837 => x"0e04b418",
			3838 => x"0b047d0c",
			3839 => x"0504e708",
			3840 => x"0504e204",
			3841 => x"fe473dc1",
			3842 => x"ff863dc1",
			3843 => x"01353dc1",
			3844 => x"0a02ed08",
			3845 => x"0704a904",
			3846 => x"fe313dc1",
			3847 => x"ff0f3dc1",
			3848 => x"00003dc1",
			3849 => x"0e04d304",
			3850 => x"03163dc1",
			3851 => x"fea83dc1",
			3852 => x"040e2324",
			3853 => x"0a02c90c",
			3854 => x"0b047f08",
			3855 => x"07046404",
			3856 => x"00003dc1",
			3857 => x"03403dc1",
			3858 => x"fe873dc1",
			3859 => x"0a02d708",
			3860 => x"0c049204",
			3861 => x"016c3dc1",
			3862 => x"035f3dc1",
			3863 => x"040da908",
			3864 => x"0803c704",
			3865 => x"fe663dc1",
			3866 => x"00e03dc1",
			3867 => x"02080204",
			3868 => x"025b3dc1",
			3869 => x"00b53dc1",
			3870 => x"0208300c",
			3871 => x"0504e508",
			3872 => x"0e02d904",
			3873 => x"fede3dc1",
			3874 => x"01683dc1",
			3875 => x"fe2f3dc1",
			3876 => x"0208830c",
			3877 => x"0e038e08",
			3878 => x"06014304",
			3879 => x"01033dc1",
			3880 => x"fee23dc1",
			3881 => x"021b3dc1",
			3882 => x"fe823dc1",
			3883 => x"06015340",
			3884 => x"05051e14",
			3885 => x"040d0008",
			3886 => x"00041404",
			3887 => x"00003dc1",
			3888 => x"02b73dc1",
			3889 => x"0004ab08",
			3890 => x"07047b04",
			3891 => x"00003dc1",
			3892 => x"00cf3dc1",
			3893 => x"fe7e3dc1",
			3894 => x"0704f118",
			3895 => x"0c04ca10",
			3896 => x"05059308",
			3897 => x"0b04e104",
			3898 => x"ff463dc1",
			3899 => x"fdba3dc1",
			3900 => x"0208eb04",
			3901 => x"01733dc1",
			3902 => x"ff1f3dc1",
			3903 => x"02090004",
			3904 => x"fd2f3dc1",
			3905 => x"fe993dc1",
			3906 => x"0004210c",
			3907 => x"0208f704",
			3908 => x"fdb53dc1",
			3909 => x"06015204",
			3910 => x"ff473dc1",
			3911 => x"01953dc1",
			3912 => x"040c9304",
			3913 => x"02133dc1",
			3914 => x"fe963dc1",
			3915 => x"0601550c",
			3916 => x"07052f04",
			3917 => x"02823dc1",
			3918 => x"09015a04",
			3919 => x"fe963dc1",
			3920 => x"00003dc1",
			3921 => x"08035a20",
			3922 => x"06015f10",
			3923 => x"040b8008",
			3924 => x"02090c04",
			3925 => x"00d83dc1",
			3926 => x"fe603dc1",
			3927 => x"02093d04",
			3928 => x"fd0d3dc1",
			3929 => x"ff593dc1",
			3930 => x"0306b908",
			3931 => x"0c04cc04",
			3932 => x"ffe43dc1",
			3933 => x"01e43dc1",
			3934 => x"05066c04",
			3935 => x"feb63dc1",
			3936 => x"00003dc1",
			3937 => x"040c1210",
			3938 => x"07050508",
			3939 => x"0c04cd04",
			3940 => x"00b43dc1",
			3941 => x"023d3dc1",
			3942 => x"08036104",
			3943 => x"02273dc1",
			3944 => x"fe933dc1",
			3945 => x"00046c08",
			3946 => x"02092004",
			3947 => x"fe223dc1",
			3948 => x"ff9f3dc1",
			3949 => x"040c6004",
			3950 => x"00cc3dc1",
			3951 => x"ffc13dc1",
			3952 => x"0c04f1b8",
			3953 => x"0c04796c",
			3954 => x"0c047640",
			3955 => x"0c047420",
			3956 => x"02089110",
			3957 => x"07049108",
			3958 => x"07048f04",
			3959 => x"ffc73fbd",
			3960 => x"00fc3fbd",
			3961 => x"02082a04",
			3962 => x"ffc63fbd",
			3963 => x"fecb3fbd",
			3964 => x"040cf508",
			3965 => x"0f072b04",
			3966 => x"033d3fbd",
			3967 => x"00ca3fbd",
			3968 => x"06014104",
			3969 => x"00003fbd",
			3970 => x"fe153fbd",
			3971 => x"0c047510",
			3972 => x"09008e08",
			3973 => x"0d050204",
			3974 => x"ff273fbd",
			3975 => x"02373fbd",
			3976 => x"0d056504",
			3977 => x"ff3f3fbd",
			3978 => x"025a3fbd",
			3979 => x"07048f08",
			3980 => x"07048004",
			3981 => x"00623fbd",
			3982 => x"030b3fbd",
			3983 => x"07049104",
			3984 => x"fdc43fbd",
			3985 => x"00293fbd",
			3986 => x"0c047710",
			3987 => x"07047a04",
			3988 => x"01163fbd",
			3989 => x"09009d08",
			3990 => x"03053704",
			3991 => x"ff083fbd",
			3992 => x"fd743fbd",
			3993 => x"007d3fbd",
			3994 => x"0704aa10",
			3995 => x"07047b08",
			3996 => x"01004304",
			3997 => x"006d3fbd",
			3998 => x"fdd33fbd",
			3999 => x"0207aa04",
			4000 => x"fe183fbd",
			4001 => x"007e3fbd",
			4002 => x"0704ad04",
			4003 => x"fded3fbd",
			4004 => x"0b04b204",
			4005 => x"00a13fbd",
			4006 => x"ff183fbd",
			4007 => x"0c048f20",
			4008 => x"0003cc04",
			4009 => x"fea43fbd",
			4010 => x"01005c10",
			4011 => x"0704ac08",
			4012 => x"0d052504",
			4013 => x"fffb3fbd",
			4014 => x"01463fbd",
			4015 => x"00043504",
			4016 => x"fda83fbd",
			4017 => x"ffe53fbd",
			4018 => x"0b04e008",
			4019 => x"03054304",
			4020 => x"029f3fbd",
			4021 => x"01da3fbd",
			4022 => x"00893fbd",
			4023 => x"01004310",
			4024 => x"03042608",
			4025 => x"0207d704",
			4026 => x"ff263fbd",
			4027 => x"02113fbd",
			4028 => x"0d053404",
			4029 => x"fe333fbd",
			4030 => x"ff883fbd",
			4031 => x"0d051a0c",
			4032 => x"0c049104",
			4033 => x"fe2f3fbd",
			4034 => x"02083104",
			4035 => x"01f53fbd",
			4036 => x"00213fbd",
			4037 => x"03052508",
			4038 => x"0d057504",
			4039 => x"ffdf3fbd",
			4040 => x"fdef3fbd",
			4041 => x"09009c04",
			4042 => x"006a3fbd",
			4043 => x"00023fbd",
			4044 => x"0f07ce0c",
			4045 => x"00042808",
			4046 => x"0b055404",
			4047 => x"00983fbd",
			4048 => x"fdfc3fbd",
			4049 => x"fe243fbd",
			4050 => x"0100951c",
			4051 => x"05063210",
			4052 => x"0a02cc0c",
			4053 => x"0a02ab08",
			4054 => x"0a029b04",
			4055 => x"fe3a3fbd",
			4056 => x"01fb3fbd",
			4057 => x"fe413fbd",
			4058 => x"026f3fbd",
			4059 => x"0b05a608",
			4060 => x"03065904",
			4061 => x"00003fbd",
			4062 => x"02f73fbd",
			4063 => x"00003fbd",
			4064 => x"00037010",
			4065 => x"0c05b80c",
			4066 => x"00031a04",
			4067 => x"00003fbd",
			4068 => x"01011704",
			4069 => x"01a03fbd",
			4070 => x"00003fbd",
			4071 => x"fec23fbd",
			4072 => x"07056104",
			4073 => x"fe483fbd",
			4074 => x"07057308",
			4075 => x"020a0004",
			4076 => x"01293fbd",
			4077 => x"00003fbd",
			4078 => x"fe8f3fbd",
			4079 => x"0a029990",
			4080 => x"08035870",
			4081 => x"00042538",
			4082 => x"0208dd20",
			4083 => x"0a027b10",
			4084 => x"06015808",
			4085 => x"01007904",
			4086 => x"fff441f9",
			4087 => x"00a041f9",
			4088 => x"0505f904",
			4089 => x"fdf441f9",
			4090 => x"000c41f9",
			4091 => x"06013d08",
			4092 => x"0e048804",
			4093 => x"ffa441f9",
			4094 => x"01fa41f9",
			4095 => x"03056104",
			4096 => x"feb441f9",
			4097 => x"006841f9",
			4098 => x"0f081608",
			4099 => x"0704d404",
			4100 => x"ff8341f9",
			4101 => x"fd5a41f9",
			4102 => x"0a028d08",
			4103 => x"0a028304",
			4104 => x"ff8841f9",
			4105 => x"017241f9",
			4106 => x"05066c04",
			4107 => x"fe7841f9",
			4108 => x"011541f9",
			4109 => x"0b04bf18",
			4110 => x"0b04be10",
			4111 => x"00043e08",
			4112 => x"08034104",
			4113 => x"000941f9",
			4114 => x"014a41f9",
			4115 => x"08035504",
			4116 => x"ff9941f9",
			4117 => x"010341f9",
			4118 => x"08034204",
			4119 => x"000041f9",
			4120 => x"02de41f9",
			4121 => x"0e04c910",
			4122 => x"0d056908",
			4123 => x"02085204",
			4124 => x"ffb441f9",
			4125 => x"fe5541f9",
			4126 => x"06014504",
			4127 => x"fdf941f9",
			4128 => x"00f641f9",
			4129 => x"0900c008",
			4130 => x"0d057304",
			4131 => x"ff6241f9",
			4132 => x"002d41f9",
			4133 => x"0b054304",
			4134 => x"fe6041f9",
			4135 => x"003841f9",
			4136 => x"0d052814",
			4137 => x"05050f10",
			4138 => x"01003f08",
			4139 => x"0004ab04",
			4140 => x"020741f9",
			4141 => x"000041f9",
			4142 => x"00046b04",
			4143 => x"ff2b41f9",
			4144 => x"fdec41f9",
			4145 => x"00de41f9",
			4146 => x"0704bc04",
			4147 => x"fd9541f9",
			4148 => x"0f074104",
			4149 => x"ff8c41f9",
			4150 => x"fe4041f9",
			4151 => x"03046f34",
			4152 => x"0a02d418",
			4153 => x"09006210",
			4154 => x"0f05fc04",
			4155 => x"fe5b41f9",
			4156 => x"0504e708",
			4157 => x"03041f04",
			4158 => x"000041f9",
			4159 => x"01ff41f9",
			4160 => x"ffae41f9",
			4161 => x"0f05e004",
			4162 => x"002141f9",
			4163 => x"fe3b41f9",
			4164 => x"06015318",
			4165 => x"00052908",
			4166 => x"0803be04",
			4167 => x"004a41f9",
			4168 => x"023541f9",
			4169 => x"03045608",
			4170 => x"05050104",
			4171 => x"001f41f9",
			4172 => x"fe4241f9",
			4173 => x"0208d404",
			4174 => x"013841f9",
			4175 => x"000041f9",
			4176 => x"fe6c41f9",
			4177 => x"02081d28",
			4178 => x"0004a718",
			4179 => x"0e03da08",
			4180 => x"0207eb04",
			4181 => x"039941f9",
			4182 => x"007e41f9",
			4183 => x"08038208",
			4184 => x"01005004",
			4185 => x"ffd641f9",
			4186 => x"00f841f9",
			4187 => x"0f069904",
			4188 => x"02c641f9",
			4189 => x"ffe541f9",
			4190 => x"03049f08",
			4191 => x"01004704",
			4192 => x"ffd741f9",
			4193 => x"fe4b41f9",
			4194 => x"01005604",
			4195 => x"016041f9",
			4196 => x"fe9941f9",
			4197 => x"02082a14",
			4198 => x"06014508",
			4199 => x"02082404",
			4200 => x"fda741f9",
			4201 => x"ff8041f9",
			4202 => x"01005104",
			4203 => x"015b41f9",
			4204 => x"01005a04",
			4205 => x"fe0c41f9",
			4206 => x"ffef41f9",
			4207 => x"0d052610",
			4208 => x"0e048508",
			4209 => x"07047d04",
			4210 => x"006441f9",
			4211 => x"ff8741f9",
			4212 => x"03051b04",
			4213 => x"fda141f9",
			4214 => x"ff6b41f9",
			4215 => x"09009d08",
			4216 => x"03053304",
			4217 => x"001641f9",
			4218 => x"00ae41f9",
			4219 => x"01006204",
			4220 => x"ff2541f9",
			4221 => x"001041f9",
			4222 => x"0a0288ac",
			4223 => x"0c049250",
			4224 => x"0704a820",
			4225 => x"05055818",
			4226 => x"0601360c",
			4227 => x"0704a708",
			4228 => x"0704a604",
			4229 => x"001b441d",
			4230 => x"fe86441d",
			4231 => x"0269441d",
			4232 => x"0b04be08",
			4233 => x"040b7804",
			4234 => x"fd7d441d",
			4235 => x"ff41441d",
			4236 => x"0016441d",
			4237 => x"0704a504",
			4238 => x"009a441d",
			4239 => x"027a441d",
			4240 => x"0c049120",
			4241 => x"01006310",
			4242 => x"040ba408",
			4243 => x"00040804",
			4244 => x"ff88441d",
			4245 => x"00ad441d",
			4246 => x"040bb204",
			4247 => x"fd3d441d",
			4248 => x"ff3d441d",
			4249 => x"0b04e108",
			4250 => x"06014204",
			4251 => x"fe29441d",
			4252 => x"0041441d",
			4253 => x"0704c404",
			4254 => x"ff64441d",
			4255 => x"017a441d",
			4256 => x"0704bf08",
			4257 => x"01005e04",
			4258 => x"fe9f441d",
			4259 => x"fd11441d",
			4260 => x"0b04d204",
			4261 => x"004f441d",
			4262 => x"fe3b441d",
			4263 => x"0c049424",
			4264 => x"01005410",
			4265 => x"0b04a008",
			4266 => x"09007e04",
			4267 => x"ff8b441d",
			4268 => x"fdf1441d",
			4269 => x"0704a904",
			4270 => x"024c441d",
			4271 => x"fe37441d",
			4272 => x"0b04e20c",
			4273 => x"03056f08",
			4274 => x"0304fe04",
			4275 => x"023e441d",
			4276 => x"fffa441d",
			4277 => x"0246441d",
			4278 => x"0704d304",
			4279 => x"0095441d",
			4280 => x"fe27441d",
			4281 => x"0207b718",
			4282 => x"0304cf08",
			4283 => x"0d054004",
			4284 => x"fe4c441d",
			4285 => x"0000441d",
			4286 => x"0a023308",
			4287 => x"03067804",
			4288 => x"fe36441d",
			4289 => x"0080441d",
			4290 => x"0c04b004",
			4291 => x"00f3441d",
			4292 => x"0262441d",
			4293 => x"0207e510",
			4294 => x"0207da08",
			4295 => x"0207d704",
			4296 => x"ff92441d",
			4297 => x"0169441d",
			4298 => x"0a025304",
			4299 => x"0000441d",
			4300 => x"fd86441d",
			4301 => x"0d058308",
			4302 => x"01006204",
			4303 => x"ffda441d",
			4304 => x"0105441d",
			4305 => x"05058304",
			4306 => x"fe99441d",
			4307 => x"0016441d",
			4308 => x"0a028a18",
			4309 => x"0c048f04",
			4310 => x"feaa441d",
			4311 => x"0d055904",
			4312 => x"03e6441d",
			4313 => x"040bcc0c",
			4314 => x"06014604",
			4315 => x"0079441d",
			4316 => x"0003ed04",
			4317 => x"0000441d",
			4318 => x"0265441d",
			4319 => x"fe26441d",
			4320 => x"0c044018",
			4321 => x"0207b504",
			4322 => x"fecd441d",
			4323 => x"06012d04",
			4324 => x"ff53441d",
			4325 => x"0c043a08",
			4326 => x"01001804",
			4327 => x"0000441d",
			4328 => x"00b6441d",
			4329 => x"00057a04",
			4330 => x"026d441d",
			4331 => x"0000441d",
			4332 => x"03049f1c",
			4333 => x"040c7210",
			4334 => x"0c045e08",
			4335 => x"0c045a04",
			4336 => x"feab441d",
			4337 => x"010c441d",
			4338 => x"0a02b004",
			4339 => x"fe97441d",
			4340 => x"fff0441d",
			4341 => x"00048604",
			4342 => x"01ee441d",
			4343 => x"040c9a04",
			4344 => x"fe4c441d",
			4345 => x"0025441d",
			4346 => x"08032b0c",
			4347 => x"040aa908",
			4348 => x"05061604",
			4349 => x"0000441d",
			4350 => x"014e441d",
			4351 => x"fd39441d",
			4352 => x"02081108",
			4353 => x"02080e04",
			4354 => x"0061441d",
			4355 => x"021b441d",
			4356 => x"040bf704",
			4357 => x"0043441d",
			4358 => x"000c441d",
			4359 => x"0b0543bc",
			4360 => x"040c6060",
			4361 => x"0e047824",
			4362 => x"0409c704",
			4363 => x"e7f24661",
			4364 => x"06013510",
			4365 => x"06012108",
			4366 => x"0b048d04",
			4367 => x"e0fb4661",
			4368 => x"de734661",
			4369 => x"03049704",
			4370 => x"df134661",
			4371 => x"e0b04661",
			4372 => x"00043a08",
			4373 => x"09008204",
			4374 => x"ea294661",
			4375 => x"e3544661",
			4376 => x"05054b04",
			4377 => x"e14a4661",
			4378 => x"de534661",
			4379 => x"0601251c",
			4380 => x"0802ee10",
			4381 => x"0a023008",
			4382 => x"06011204",
			4383 => x"de0c4661",
			4384 => x"def14661",
			4385 => x"040a9504",
			4386 => x"e39e4661",
			4387 => x"dea74661",
			4388 => x"09009508",
			4389 => x"040b3604",
			4390 => x"e80a4661",
			4391 => x"e0324661",
			4392 => x"de284661",
			4393 => x"040bcc10",
			4394 => x"06013908",
			4395 => x"0207ed04",
			4396 => x"e7704661",
			4397 => x"e3b34661",
			4398 => x"07050404",
			4399 => x"e81a4661",
			4400 => x"e2634661",
			4401 => x"0704aa08",
			4402 => x"06014f04",
			4403 => x"e5434661",
			4404 => x"e94e4661",
			4405 => x"0e054404",
			4406 => x"e25e4661",
			4407 => x"e4784661",
			4408 => x"0601341c",
			4409 => x"040ca70c",
			4410 => x"00045f04",
			4411 => x"de254661",
			4412 => x"00048604",
			4413 => x"e59e4661",
			4414 => x"e0624661",
			4415 => x"01003904",
			4416 => x"de074661",
			4417 => x"040ce104",
			4418 => x"de304661",
			4419 => x"09006c04",
			4420 => x"e0324661",
			4421 => x"de3c4661",
			4422 => x"09008620",
			4423 => x"0004a010",
			4424 => x"0304fe08",
			4425 => x"040ca004",
			4426 => x"e1564661",
			4427 => x"e4664661",
			4428 => x"0704a604",
			4429 => x"e8dd4661",
			4430 => x"e4334661",
			4431 => x"040cf508",
			4432 => x"0304c704",
			4433 => x"dec64661",
			4434 => x"e11c4661",
			4435 => x"040fc604",
			4436 => x"e2354661",
			4437 => x"de174661",
			4438 => x"0e054b10",
			4439 => x"05054b08",
			4440 => x"00048a04",
			4441 => x"e23e4661",
			4442 => x"df944661",
			4443 => x"02081d04",
			4444 => x"e20a4661",
			4445 => x"dee94661",
			4446 => x"040c7f08",
			4447 => x"08037e04",
			4448 => x"dfe04661",
			4449 => x"e7d44661",
			4450 => x"0f082b04",
			4451 => x"dffb4661",
			4452 => x"e3234661",
			4453 => x"0705323c",
			4454 => x"06017428",
			4455 => x"03065010",
			4456 => x"0505db04",
			4457 => x"e1ba4661",
			4458 => x"03061904",
			4459 => x"de0a4661",
			4460 => x"07051b04",
			4461 => x"e1f14661",
			4462 => x"de214661",
			4463 => x"0a026108",
			4464 => x"06013d04",
			4465 => x"e3404661",
			4466 => x"e90c4661",
			4467 => x"0900fb08",
			4468 => x"0b057404",
			4469 => x"e1554661",
			4470 => x"e5bb4661",
			4471 => x"00040b04",
			4472 => x"de3c4661",
			4473 => x"df8e4661",
			4474 => x"06017910",
			4475 => x"07050304",
			4476 => x"e1964661",
			4477 => x"0f087204",
			4478 => x"de134661",
			4479 => x"01009d04",
			4480 => x"de3c4661",
			4481 => x"e09c4661",
			4482 => x"de0a4661",
			4483 => x"0705751c",
			4484 => x"0e062e0c",
			4485 => x"0b056308",
			4486 => x"05060604",
			4487 => x"de334661",
			4488 => x"df6c4661",
			4489 => x"de084661",
			4490 => x"0209810c",
			4491 => x"00033e04",
			4492 => x"de114661",
			4493 => x"0b059904",
			4494 => x"df994661",
			4495 => x"e83b4661",
			4496 => x"de0e4661",
			4497 => x"0802c70c",
			4498 => x"0a021d04",
			4499 => x"de074661",
			4500 => x"0802bb04",
			4501 => x"de2e4661",
			4502 => x"de684661",
			4503 => x"de074661",
			4504 => x"080329a8",
			4505 => x"08031d64",
			4506 => x"0d05332c",
			4507 => x"0704921c",
			4508 => x"0c047510",
			4509 => x"03049f08",
			4510 => x"07046c04",
			4511 => x"000048b5",
			4512 => x"02df48b5",
			4513 => x"0304f704",
			4514 => x"ff4648b5",
			4515 => x"01e148b5",
			4516 => x"0d052608",
			4517 => x"09007104",
			4518 => x"000048b5",
			4519 => x"fe2648b5",
			4520 => x"007548b5",
			4521 => x"0207c50c",
			4522 => x"03049704",
			4523 => x"000b48b5",
			4524 => x"0e044b04",
			4525 => x"037e48b5",
			4526 => x"013748b5",
			4527 => x"ff7548b5",
			4528 => x"0e04e918",
			4529 => x"07049008",
			4530 => x"01005104",
			4531 => x"ff5948b5",
			4532 => x"02db48b5",
			4533 => x"0b04b008",
			4534 => x"00040b04",
			4535 => x"fe1948b5",
			4536 => x"ff8148b5",
			4537 => x"0b04b904",
			4538 => x"009648b5",
			4539 => x"ff6d48b5",
			4540 => x"0704a910",
			4541 => x"02081b08",
			4542 => x"05055904",
			4543 => x"000048b5",
			4544 => x"017248b5",
			4545 => x"040b4a04",
			4546 => x"020448b5",
			4547 => x"031948b5",
			4548 => x"040b5008",
			4549 => x"0003e204",
			4550 => x"ffd148b5",
			4551 => x"00c848b5",
			4552 => x"0d05a904",
			4553 => x"ffa648b5",
			4554 => x"fd3648b5",
			4555 => x"02084524",
			4556 => x"0a026f10",
			4557 => x"0004200c",
			4558 => x"0a026904",
			4559 => x"000048b5",
			4560 => x"0b04c204",
			4561 => x"fdc348b5",
			4562 => x"ff1c48b5",
			4563 => x"005d48b5",
			4564 => x"0003ee04",
			4565 => x"fd6148b5",
			4566 => x"03054308",
			4567 => x"0207f804",
			4568 => x"008a48b5",
			4569 => x"fee148b5",
			4570 => x"0c04ae04",
			4571 => x"020448b5",
			4572 => x"001248b5",
			4573 => x"01007910",
			4574 => x"0e05b30c",
			4575 => x"0e057808",
			4576 => x"0208a604",
			4577 => x"fe6e48b5",
			4578 => x"01f448b5",
			4579 => x"01ef48b5",
			4580 => x"fc6948b5",
			4581 => x"0a028d0c",
			4582 => x"02090908",
			4583 => x"0e05e004",
			4584 => x"fefa48b5",
			4585 => x"016048b5",
			4586 => x"fdc948b5",
			4587 => x"fd7c48b5",
			4588 => x"08032e2c",
			4589 => x"0208911c",
			4590 => x"0c045b04",
			4591 => x"02d648b5",
			4592 => x"0a027508",
			4593 => x"0a027204",
			4594 => x"000a48b5",
			4595 => x"fe3c48b5",
			4596 => x"05055908",
			4597 => x"01006104",
			4598 => x"012d48b5",
			4599 => x"feb848b5",
			4600 => x"0d059d04",
			4601 => x"023748b5",
			4602 => x"011748b5",
			4603 => x"0208f708",
			4604 => x"01007b04",
			4605 => x"fff448b5",
			4606 => x"fccb48b5",
			4607 => x"07054504",
			4608 => x"01f748b5",
			4609 => x"ffc148b5",
			4610 => x"08033118",
			4611 => x"00042514",
			4612 => x"040bb00c",
			4613 => x"0e04ad04",
			4614 => x"011a48b5",
			4615 => x"0e056804",
			4616 => x"fdec48b5",
			4617 => x"001248b5",
			4618 => x"00041d04",
			4619 => x"000048b5",
			4620 => x"03f348b5",
			4621 => x"fdc948b5",
			4622 => x"00043920",
			4623 => x"08033410",
			4624 => x"0a028308",
			4625 => x"01006304",
			4626 => x"ffaf48b5",
			4627 => x"fd2848b5",
			4628 => x"040ba404",
			4629 => x"015a48b5",
			4630 => x"ff3f48b5",
			4631 => x"02087608",
			4632 => x"040b5604",
			4633 => x"ffa548b5",
			4634 => x"011248b5",
			4635 => x"040baa04",
			4636 => x"008048b5",
			4637 => x"ff0b48b5",
			4638 => x"05054a10",
			4639 => x"01005e08",
			4640 => x"09009a04",
			4641 => x"002f48b5",
			4642 => x"fe8248b5",
			4643 => x"0c049404",
			4644 => x"01e648b5",
			4645 => x"000048b5",
			4646 => x"040c6608",
			4647 => x"0e04f704",
			4648 => x"ffbf48b5",
			4649 => x"003248b5",
			4650 => x"08035304",
			4651 => x"045a48b5",
			4652 => x"ff5e48b5",
			4653 => x"0c0548cc",
			4654 => x"0a029e60",
			4655 => x"0207da2c",
			4656 => x"0207d720",
			4657 => x"0a023910",
			4658 => x"0b049e08",
			4659 => x"0f064a04",
			4660 => x"02584a69",
			4661 => x"fee74a69",
			4662 => x"0f070f04",
			4663 => x"fe884a69",
			4664 => x"00824a69",
			4665 => x"02077708",
			4666 => x"0802e604",
			4667 => x"02104a69",
			4668 => x"ff104a69",
			4669 => x"0f064a04",
			4670 => x"01dc4a69",
			4671 => x"00904a69",
			4672 => x"05051d04",
			4673 => x"ff974a69",
			4674 => x"0d054004",
			4675 => x"03de4a69",
			4676 => x"01da4a69",
			4677 => x"0505f91c",
			4678 => x"02089010",
			4679 => x"0e04bb08",
			4680 => x"09008c04",
			4681 => x"000f4a69",
			4682 => x"ff6c4a69",
			4683 => x"08032504",
			4684 => x"ffea4a69",
			4685 => x"00884a69",
			4686 => x"0c04ef08",
			4687 => x"00043e04",
			4688 => x"ff2f4a69",
			4689 => x"ffd74a69",
			4690 => x"01fa4a69",
			4691 => x"0e065a0c",
			4692 => x"0c050708",
			4693 => x"03066904",
			4694 => x"01544a69",
			4695 => x"04014a69",
			4696 => x"005f4a69",
			4697 => x"01008a04",
			4698 => x"fe3b4a69",
			4699 => x"00037d04",
			4700 => x"02074a69",
			4701 => x"00364a69",
			4702 => x"040c1840",
			4703 => x"0900c620",
			4704 => x"02089110",
			4705 => x"09009508",
			4706 => x"00046b04",
			4707 => x"02994a69",
			4708 => x"00984a69",
			4709 => x"00044304",
			4710 => x"02154a69",
			4711 => x"ffb14a69",
			4712 => x"0b050108",
			4713 => x"0900b704",
			4714 => x"01624a69",
			4715 => x"ffaf4a69",
			4716 => x"08035b04",
			4717 => x"00794a69",
			4718 => x"02884a69",
			4719 => x"02091910",
			4720 => x"00044708",
			4721 => x"0d060304",
			4722 => x"01784a69",
			4723 => x"ff214a69",
			4724 => x"03062104",
			4725 => x"fe1b4a69",
			4726 => x"ffd74a69",
			4727 => x"0b054508",
			4728 => x"0505ce04",
			4729 => x"009a4a69",
			4730 => x"029d4a69",
			4731 => x"0a02a504",
			4732 => x"02c44a69",
			4733 => x"ff204a69",
			4734 => x"03041f0c",
			4735 => x"00051504",
			4736 => x"fe214a69",
			4737 => x"040fc604",
			4738 => x"00ab4a69",
			4739 => x"fe764a69",
			4740 => x"0f06a510",
			4741 => x"0304df08",
			4742 => x"09008704",
			4743 => x"00b04a69",
			4744 => x"fe414a69",
			4745 => x"01005a04",
			4746 => x"05254a69",
			4747 => x"030e4a69",
			4748 => x"0c047208",
			4749 => x"0c045b04",
			4750 => x"00134a69",
			4751 => x"02104a69",
			4752 => x"0304c004",
			4753 => x"fed14a69",
			4754 => x"001e4a69",
			4755 => x"0c05b80c",
			4756 => x"00036308",
			4757 => x"00035304",
			4758 => x"febc4a69",
			4759 => x"02514a69",
			4760 => x"fe774a69",
			4761 => x"fe684a69",
			4762 => x"0f06fb84",
			4763 => x"03054358",
			4764 => x"0d057434",
			4765 => x"05056520",
			4766 => x"0b04cf10",
			4767 => x"01005c08",
			4768 => x"05055704",
			4769 => x"00134cc5",
			4770 => x"ff074cc5",
			4771 => x"0900a004",
			4772 => x"00ea4cc5",
			4773 => x"fec04cc5",
			4774 => x"040b2908",
			4775 => x"01005804",
			4776 => x"fed04cc5",
			4777 => x"01564cc5",
			4778 => x"01005604",
			4779 => x"00004cc5",
			4780 => x"fe854cc5",
			4781 => x"040ae204",
			4782 => x"fdf54cc5",
			4783 => x"040be908",
			4784 => x"040b9d04",
			4785 => x"009a4cc5",
			4786 => x"02784cc5",
			4787 => x"040c2404",
			4788 => x"fe584cc5",
			4789 => x"00e84cc5",
			4790 => x"0f06e31c",
			4791 => x"0d058d10",
			4792 => x"03052508",
			4793 => x"0704bf04",
			4794 => x"002b4cc5",
			4795 => x"fe4b4cc5",
			4796 => x"06013404",
			4797 => x"ff9f4cc5",
			4798 => x"018c4cc5",
			4799 => x"0b050404",
			4800 => x"fe484cc5",
			4801 => x"06014504",
			4802 => x"fff04cc5",
			4803 => x"00f14cc5",
			4804 => x"01005704",
			4805 => x"00004cc5",
			4806 => x"fdad4cc5",
			4807 => x"0704bc10",
			4808 => x"07049404",
			4809 => x"feb04cc5",
			4810 => x"06012b04",
			4811 => x"00764cc5",
			4812 => x"0e04e204",
			4813 => x"02ee4cc5",
			4814 => x"01a84cc5",
			4815 => x"09009c0c",
			4816 => x"0f06ca04",
			4817 => x"fe884cc5",
			4818 => x"03055304",
			4819 => x"025f4cc5",
			4820 => x"010b4cc5",
			4821 => x"0b04c104",
			4822 => x"fddd4cc5",
			4823 => x"03054804",
			4824 => x"026d4cc5",
			4825 => x"06013e04",
			4826 => x"00594cc5",
			4827 => x"feea4cc5",
			4828 => x"03055334",
			4829 => x"03054f28",
			4830 => x"05057620",
			4831 => x"05055710",
			4832 => x"0b04d008",
			4833 => x"0d056704",
			4834 => x"ffe34cc5",
			4835 => x"fe934cc5",
			4836 => x"0704c004",
			4837 => x"ffed4cc5",
			4838 => x"02d54cc5",
			4839 => x"01006308",
			4840 => x"0e04a904",
			4841 => x"fde24cc5",
			4842 => x"ff1e4cc5",
			4843 => x"0704d304",
			4844 => x"01c44cc5",
			4845 => x"fe584cc5",
			4846 => x"0704d504",
			4847 => x"02da4cc5",
			4848 => x"ff7c4cc5",
			4849 => x"0900a008",
			4850 => x"0d054104",
			4851 => x"00004cc5",
			4852 => x"fded4cc5",
			4853 => x"fff94cc5",
			4854 => x"040bfa38",
			4855 => x"01006920",
			4856 => x"00041810",
			4857 => x"06013008",
			4858 => x"0d057504",
			4859 => x"01854cc5",
			4860 => x"ff754cc5",
			4861 => x"03056f04",
			4862 => x"00484cc5",
			4863 => x"ff494cc5",
			4864 => x"01005e08",
			4865 => x"0b04ae04",
			4866 => x"01ae4cc5",
			4867 => x"ff8e4cc5",
			4868 => x"0b04c104",
			4869 => x"002a4cc5",
			4870 => x"01254cc5",
			4871 => x"0b04d20c",
			4872 => x"0305d908",
			4873 => x"0d057604",
			4874 => x"ffa64cc5",
			4875 => x"fde64cc5",
			4876 => x"010f4cc5",
			4877 => x"0d057504",
			4878 => x"02b84cc5",
			4879 => x"00046704",
			4880 => x"000d4cc5",
			4881 => x"fe834cc5",
			4882 => x"08036120",
			4883 => x"0b04e010",
			4884 => x"01006008",
			4885 => x"0d053304",
			4886 => x"014a4cc5",
			4887 => x"fe264cc5",
			4888 => x"0d057404",
			4889 => x"011f4cc5",
			4890 => x"ffd84cc5",
			4891 => x"0a029008",
			4892 => x"08033704",
			4893 => x"ffcb4cc5",
			4894 => x"01094cc5",
			4895 => x"00045304",
			4896 => x"fe2e4cc5",
			4897 => x"ff1d4cc5",
			4898 => x"040c6010",
			4899 => x"06016308",
			4900 => x"0704ea04",
			4901 => x"00284cc5",
			4902 => x"00f74cc5",
			4903 => x"0f07c704",
			4904 => x"fe524cc5",
			4905 => x"ffe64cc5",
			4906 => x"0a02c408",
			4907 => x"05054b04",
			4908 => x"00954cc5",
			4909 => x"feeb4cc5",
			4910 => x"0f076b04",
			4911 => x"018f4cc5",
			4912 => x"00184cc5",
			4913 => x"0a0283ac",
			4914 => x"08031b58",
			4915 => x"08030f30",
			4916 => x"040b0214",
			4917 => x"0003f310",
			4918 => x"040aef08",
			4919 => x"040ac204",
			4920 => x"003e4f29",
			4921 => x"ff914f29",
			4922 => x"0b04e104",
			4923 => x"01fc4f29",
			4924 => x"ffae4f29",
			4925 => x"fe3a4f29",
			4926 => x"0a026710",
			4927 => x"0a025c08",
			4928 => x"0e04d304",
			4929 => x"ff184f29",
			4930 => x"009e4f29",
			4931 => x"040b7604",
			4932 => x"fe264f29",
			4933 => x"00944f29",
			4934 => x"0a026c08",
			4935 => x"0003d904",
			4936 => x"00004f29",
			4937 => x"02004f29",
			4938 => x"fe4d4f29",
			4939 => x"040aa108",
			4940 => x"0d05ed04",
			4941 => x"fded4f29",
			4942 => x"00004f29",
			4943 => x"040b6310",
			4944 => x"00040808",
			4945 => x"00040304",
			4946 => x"00f14f29",
			4947 => x"ff384f29",
			4948 => x"0e048804",
			4949 => x"00714f29",
			4950 => x"026b4f29",
			4951 => x"0704a708",
			4952 => x"0304f704",
			4953 => x"ff114f29",
			4954 => x"02254f29",
			4955 => x"0b04b904",
			4956 => x"003b4f29",
			4957 => x"feac4f29",
			4958 => x"0a027020",
			4959 => x"0c04760c",
			4960 => x"00041404",
			4961 => x"fe314f29",
			4962 => x"05050f04",
			4963 => x"ff0c4f29",
			4964 => x"01be4f29",
			4965 => x"0704be10",
			4966 => x"09008f08",
			4967 => x"09008704",
			4968 => x"fe304f29",
			4969 => x"00004f29",
			4970 => x"0c049204",
			4971 => x"fe494f29",
			4972 => x"fd1b4f29",
			4973 => x"ffe84f29",
			4974 => x"0d058318",
			4975 => x"00042e0c",
			4976 => x"040aef04",
			4977 => x"fe414f29",
			4978 => x"040b2204",
			4979 => x"01d94f29",
			4980 => x"00484f29",
			4981 => x"040b8a04",
			4982 => x"fd9b4f29",
			4983 => x"0c049604",
			4984 => x"ff814f29",
			4985 => x"01544f29",
			4986 => x"0505840c",
			4987 => x"0704a604",
			4988 => x"004f4f29",
			4989 => x"0704bf04",
			4990 => x"fc2d4f29",
			4991 => x"fe7c4f29",
			4992 => x"0505bd08",
			4993 => x"01007104",
			4994 => x"ffed4f29",
			4995 => x"01394f29",
			4996 => x"040b5b04",
			4997 => x"000e4f29",
			4998 => x"fdd84f29",
			4999 => x"040b914c",
			5000 => x"00040c18",
			5001 => x"02086004",
			5002 => x"fd8e4f29",
			5003 => x"040b6b10",
			5004 => x"040b1608",
			5005 => x"03063204",
			5006 => x"fe4e4f29",
			5007 => x"00004f29",
			5008 => x"0900ef04",
			5009 => x"01c24f29",
			5010 => x"fe914f29",
			5011 => x"fd624f29",
			5012 => x"0004391c",
			5013 => x"0d05dc10",
			5014 => x"0a029008",
			5015 => x"040b8004",
			5016 => x"01094f29",
			5017 => x"ffc74f29",
			5018 => x"040b5604",
			5019 => x"01044f29",
			5020 => x"01f84f29",
			5021 => x"0505bf04",
			5022 => x"fe9d4f29",
			5023 => x"0c04e904",
			5024 => x"01514f29",
			5025 => x"ffca4f29",
			5026 => x"02085908",
			5027 => x"0a029304",
			5028 => x"fd804f29",
			5029 => x"ff734f29",
			5030 => x"0704ed08",
			5031 => x"08035304",
			5032 => x"01d04f29",
			5033 => x"00004f29",
			5034 => x"00043f04",
			5035 => x"ff964f29",
			5036 => x"fe394f29",
			5037 => x"00042108",
			5038 => x"08033e04",
			5039 => x"feb14f29",
			5040 => x"fdb74f29",
			5041 => x"0b055220",
			5042 => x"0900b310",
			5043 => x"0b051108",
			5044 => x"0e053e04",
			5045 => x"000c4f29",
			5046 => x"008f4f29",
			5047 => x"0305cc04",
			5048 => x"023e4f29",
			5049 => x"ffed4f29",
			5050 => x"0e055a08",
			5051 => x"00044e04",
			5052 => x"ffc94f29",
			5053 => x"fea34f29",
			5054 => x"0c04af04",
			5055 => x"ff484f29",
			5056 => x"00344f29",
			5057 => x"02099a10",
			5058 => x"0c050b08",
			5059 => x"0e05ce04",
			5060 => x"038c4f29",
			5061 => x"011e4f29",
			5062 => x"0900e904",
			5063 => x"ff1a4f29",
			5064 => x"015e4f29",
			5065 => x"fe904f29",
			5066 => x"0900b7c4",
			5067 => x"0704c458",
			5068 => x"0704c140",
			5069 => x"0704ad20",
			5070 => x"0704ac10",
			5071 => x"0704aa08",
			5072 => x"0c04b404",
			5073 => x"00155165",
			5074 => x"01875165",
			5075 => x"08039604",
			5076 => x"ff445165",
			5077 => x"01ad5165",
			5078 => x"09008a08",
			5079 => x"0b04b004",
			5080 => x"fe295165",
			5081 => x"00d85165",
			5082 => x"0e046804",
			5083 => x"ff8a5165",
			5084 => x"fdc75165",
			5085 => x"09009c10",
			5086 => x"01005c08",
			5087 => x"0b04b004",
			5088 => x"01205165",
			5089 => x"000a5165",
			5090 => x"02083304",
			5091 => x"020d5165",
			5092 => x"00a45165",
			5093 => x"0704be08",
			5094 => x"08032104",
			5095 => x"ff985165",
			5096 => x"00a15165",
			5097 => x"00042804",
			5098 => x"00ae5165",
			5099 => x"ff1d5165",
			5100 => x"01006d14",
			5101 => x"0f07c710",
			5102 => x"06014f08",
			5103 => x"0c049804",
			5104 => x"fe6b5165",
			5105 => x"ff745165",
			5106 => x"0c049504",
			5107 => x"03565165",
			5108 => x"ffad5165",
			5109 => x"fd315165",
			5110 => x"fcde5165",
			5111 => x"0e04f030",
			5112 => x"0b04cf18",
			5113 => x"0704d710",
			5114 => x"0e046108",
			5115 => x"0207e504",
			5116 => x"01a65165",
			5117 => x"feee5165",
			5118 => x"0f071f04",
			5119 => x"02cb5165",
			5120 => x"00655165",
			5121 => x"06014904",
			5122 => x"fd3a5165",
			5123 => x"ffe95165",
			5124 => x"03052508",
			5125 => x"08032c04",
			5126 => x"00005165",
			5127 => x"fe365165",
			5128 => x"0f06c108",
			5129 => x"03053f04",
			5130 => x"02955165",
			5131 => x"00955165",
			5132 => x"0900a204",
			5133 => x"001b5165",
			5134 => x"fefa5165",
			5135 => x"0900a420",
			5136 => x"08036610",
			5137 => x"0704d508",
			5138 => x"0e051004",
			5139 => x"02465165",
			5140 => x"00d15165",
			5141 => x"0704d804",
			5142 => x"fe595165",
			5143 => x"01325165",
			5144 => x"040c6c08",
			5145 => x"0c04af04",
			5146 => x"01fd5165",
			5147 => x"038b5165",
			5148 => x"0305b904",
			5149 => x"ff505165",
			5150 => x"02b15165",
			5151 => x"0c049710",
			5152 => x"06014f08",
			5153 => x"0f071d04",
			5154 => x"030b5165",
			5155 => x"009e5165",
			5156 => x"0f078e04",
			5157 => x"00e15165",
			5158 => x"030a5165",
			5159 => x"0c049c04",
			5160 => x"fd985165",
			5161 => x"01006804",
			5162 => x"ffa65165",
			5163 => x"00a65165",
			5164 => x"0f06f310",
			5165 => x"0802ae0c",
			5166 => x"03061904",
			5167 => x"fe4c5165",
			5168 => x"0e05ce04",
			5169 => x"00005165",
			5170 => x"ffb45165",
			5171 => x"037a5165",
			5172 => x"0305a914",
			5173 => x"01006f04",
			5174 => x"ffe75165",
			5175 => x"02083304",
			5176 => x"ff995165",
			5177 => x"040b9104",
			5178 => x"fc545165",
			5179 => x"0704ed04",
			5180 => x"fdd75165",
			5181 => x"fee95165",
			5182 => x"0c049618",
			5183 => x"0c049108",
			5184 => x"0208db04",
			5185 => x"01c25165",
			5186 => x"ff005165",
			5187 => x"0704d408",
			5188 => x"0704c204",
			5189 => x"fea55165",
			5190 => x"011d5165",
			5191 => x"0b051104",
			5192 => x"fd195165",
			5193 => x"ffc25165",
			5194 => x"0704d410",
			5195 => x"0e058e08",
			5196 => x"0305d904",
			5197 => x"00515165",
			5198 => x"fe4d5165",
			5199 => x"06014a04",
			5200 => x"005e5165",
			5201 => x"01df5165",
			5202 => x"06013a08",
			5203 => x"02083104",
			5204 => x"00185165",
			5205 => x"fe005165",
			5206 => x"040b5b04",
			5207 => x"00555165",
			5208 => x"ffc85165",
			5209 => x"0c0548d0",
			5210 => x"0a029e6c",
			5211 => x"0207da30",
			5212 => x"0207d11c",
			5213 => x"0a02390c",
			5214 => x"0b048d04",
			5215 => x"024f5321",
			5216 => x"06012404",
			5217 => x"fe565321",
			5218 => x"fffd5321",
			5219 => x"02077708",
			5220 => x"0802e604",
			5221 => x"024b5321",
			5222 => x"fef95321",
			5223 => x"040c1204",
			5224 => x"00ae5321",
			5225 => x"02f15321",
			5226 => x"0c04b310",
			5227 => x"08033a08",
			5228 => x"040b8a04",
			5229 => x"024c5321",
			5230 => x"05485321",
			5231 => x"040bff04",
			5232 => x"ff185321",
			5233 => x"042d5321",
			5234 => x"ff6d5321",
			5235 => x"06014a20",
			5236 => x"02089810",
			5237 => x"0a029d08",
			5238 => x"06013504",
			5239 => x"ffb25321",
			5240 => x"00325321",
			5241 => x"0c049304",
			5242 => x"fdbe5321",
			5243 => x"ffe45321",
			5244 => x"01006708",
			5245 => x"01006304",
			5246 => x"ff155321",
			5247 => x"00f75321",
			5248 => x"02089f04",
			5249 => x"00335321",
			5250 => x"fe075321",
			5251 => x"0900a90c",
			5252 => x"08035808",
			5253 => x"040bf104",
			5254 => x"01db5321",
			5255 => x"00a95321",
			5256 => x"ff545321",
			5257 => x"040bd808",
			5258 => x"0003ea04",
			5259 => x"ff965321",
			5260 => x"008f5321",
			5261 => x"0b055204",
			5262 => x"fee05321",
			5263 => x"02d75321",
			5264 => x"040c1840",
			5265 => x"0900c620",
			5266 => x"02089110",
			5267 => x"0900a008",
			5268 => x"08037104",
			5269 => x"01c45321",
			5270 => x"ff985321",
			5271 => x"00045204",
			5272 => x"014c5321",
			5273 => x"fee75321",
			5274 => x"0c04b308",
			5275 => x"0c04b104",
			5276 => x"014a5321",
			5277 => x"ff585321",
			5278 => x"05059104",
			5279 => x"012a5321",
			5280 => x"02fe5321",
			5281 => x"02093510",
			5282 => x"00044708",
			5283 => x"0d060304",
			5284 => x"01aa5321",
			5285 => x"ff2f5321",
			5286 => x"0e05bb04",
			5287 => x"fdd95321",
			5288 => x"ffba5321",
			5289 => x"0e070108",
			5290 => x"040b9d04",
			5291 => x"058e5321",
			5292 => x"01ac5321",
			5293 => x"07054904",
			5294 => x"fe725321",
			5295 => x"01d85321",
			5296 => x"0a031020",
			5297 => x"08035e10",
			5298 => x"0704bd08",
			5299 => x"09008404",
			5300 => x"fea85321",
			5301 => x"026f5321",
			5302 => x"08035604",
			5303 => x"00335321",
			5304 => x"fdd95321",
			5305 => x"00045b08",
			5306 => x"08036804",
			5307 => x"fde35321",
			5308 => x"00055321",
			5309 => x"0e03e704",
			5310 => x"ffb35321",
			5311 => x"00625321",
			5312 => x"fe655321",
			5313 => x"0c05b80c",
			5314 => x"00036308",
			5315 => x"00035304",
			5316 => x"fea65321",
			5317 => x"02c75321",
			5318 => x"fe715321",
			5319 => x"fe665321",
			5320 => x"0f0773d0",
			5321 => x"03050068",
			5322 => x"09008230",
			5323 => x"01004d1c",
			5324 => x"0d054010",
			5325 => x"0304ef08",
			5326 => x"0f06ed04",
			5327 => x"000c55cd",
			5328 => x"ff3755cd",
			5329 => x"0c045704",
			5330 => x"fe0b55cd",
			5331 => x"018355cd",
			5332 => x"01004708",
			5333 => x"0e041604",
			5334 => x"fecc55cd",
			5335 => x"018255cd",
			5336 => x"fe4455cd",
			5337 => x"0208620c",
			5338 => x"0e047108",
			5339 => x"08036e04",
			5340 => x"000055cd",
			5341 => x"015a55cd",
			5342 => x"028c55cd",
			5343 => x"0304d604",
			5344 => x"002d55cd",
			5345 => x"fe2655cd",
			5346 => x"01005318",
			5347 => x"07048f08",
			5348 => x"05051e04",
			5349 => x"fea555cd",
			5350 => x"023f55cd",
			5351 => x"0c049608",
			5352 => x"06011904",
			5353 => x"004f55cd",
			5354 => x"fe6e55cd",
			5355 => x"0704ad04",
			5356 => x"009755cd",
			5357 => x"fe2d55cd",
			5358 => x"0c047810",
			5359 => x"0c047608",
			5360 => x"0f06d004",
			5361 => x"001a55cd",
			5362 => x"fe3655cd",
			5363 => x"0304e704",
			5364 => x"ff3d55cd",
			5365 => x"fe0e55cd",
			5366 => x"05054908",
			5367 => x"08036b04",
			5368 => x"010155cd",
			5369 => x"ff9055cd",
			5370 => x"0704bb04",
			5371 => x"fe1c55cd",
			5372 => x"000055cd",
			5373 => x"0704902c",
			5374 => x"0100571c",
			5375 => x"040b8a0c",
			5376 => x"040b3008",
			5377 => x"0c045b04",
			5378 => x"013755cd",
			5379 => x"ff5b55cd",
			5380 => x"fd2c55cd",
			5381 => x"02089108",
			5382 => x"0a02a904",
			5383 => x"00e255cd",
			5384 => x"02c055cd",
			5385 => x"08037604",
			5386 => x"fe8055cd",
			5387 => x"007f55cd",
			5388 => x"02083f0c",
			5389 => x"0d054d04",
			5390 => x"ff1055cd",
			5391 => x"05055504",
			5392 => x"01f455cd",
			5393 => x"00be55cd",
			5394 => x"024c55cd",
			5395 => x"0704ee20",
			5396 => x"0c04d110",
			5397 => x"0c04d008",
			5398 => x"0c04af04",
			5399 => x"000b55cd",
			5400 => x"006e55cd",
			5401 => x"0a02a804",
			5402 => x"fe2455cd",
			5403 => x"009055cd",
			5404 => x"05058408",
			5405 => x"0d058004",
			5406 => x"010655cd",
			5407 => x"02cb55cd",
			5408 => x"0e052004",
			5409 => x"ff6255cd",
			5410 => x"014a55cd",
			5411 => x"08035210",
			5412 => x"0505b108",
			5413 => x"0e054b04",
			5414 => x"ffbb55cd",
			5415 => x"022f55cd",
			5416 => x"0c04b604",
			5417 => x"fdf755cd",
			5418 => x"ffcb55cd",
			5419 => x"0900ad08",
			5420 => x"05059504",
			5421 => x"fea455cd",
			5422 => x"006555cd",
			5423 => x"fe2855cd",
			5424 => x"0e059d50",
			5425 => x"0f07ce30",
			5426 => x"0f07a61c",
			5427 => x"0208740c",
			5428 => x"02086808",
			5429 => x"06014504",
			5430 => x"ff4955cd",
			5431 => x"00b455cd",
			5432 => x"fd0d55cd",
			5433 => x"0704bf08",
			5434 => x"03056804",
			5435 => x"ff5855cd",
			5436 => x"00d055cd",
			5437 => x"0704d804",
			5438 => x"ff2955cd",
			5439 => x"003e55cd",
			5440 => x"07050310",
			5441 => x"06015708",
			5442 => x"0900b104",
			5443 => x"ff9355cd",
			5444 => x"fe4c55cd",
			5445 => x"0208e204",
			5446 => x"00c555cd",
			5447 => x"ff2355cd",
			5448 => x"fdab55cd",
			5449 => x"0208e204",
			5450 => x"022955cd",
			5451 => x"0900b50c",
			5452 => x"040d0008",
			5453 => x"01006c04",
			5454 => x"008f55cd",
			5455 => x"021155cd",
			5456 => x"fe8155cd",
			5457 => x"0c04ce08",
			5458 => x"040c4c04",
			5459 => x"fd8855cd",
			5460 => x"ff5f55cd",
			5461 => x"07050304",
			5462 => x"009255cd",
			5463 => x"fe6955cd",
			5464 => x"0e05ac1c",
			5465 => x"0c04cf14",
			5466 => x"0505af10",
			5467 => x"0305e908",
			5468 => x"0305d104",
			5469 => x"00f855cd",
			5470 => x"fe7055cd",
			5471 => x"02090504",
			5472 => x"01fc55cd",
			5473 => x"009755cd",
			5474 => x"fdfc55cd",
			5475 => x"0900cb04",
			5476 => x"028855cd",
			5477 => x"ff4255cd",
			5478 => x"0704aa04",
			5479 => x"01b755cd",
			5480 => x"01006908",
			5481 => x"040c0c04",
			5482 => x"ff1d55cd",
			5483 => x"fda655cd",
			5484 => x"0f087208",
			5485 => x"0f07d504",
			5486 => x"004b55cd",
			5487 => x"ffb155cd",
			5488 => x"0f08bf04",
			5489 => x"00fa55cd",
			5490 => x"ff9255cd",
			5491 => x"0c059cd4",
			5492 => x"0f074958",
			5493 => x"0d05d140",
			5494 => x"0e047820",
			5495 => x"0704c110",
			5496 => x"01005c08",
			5497 => x"05053104",
			5498 => x"0023577b",
			5499 => x"ff7c577b",
			5500 => x"0b04b904",
			5501 => x"0353577b",
			5502 => x"0042577b",
			5503 => x"05054908",
			5504 => x"0a02d104",
			5505 => x"fe18577b",
			5506 => x"0087577b",
			5507 => x"09008f04",
			5508 => x"0149577b",
			5509 => x"fe9b577b",
			5510 => x"040ca010",
			5511 => x"09008c08",
			5512 => x"0d053404",
			5513 => x"0010577b",
			5514 => x"0171577b",
			5515 => x"01005504",
			5516 => x"feaa577b",
			5517 => x"0043577b",
			5518 => x"02087608",
			5519 => x"0a02cc04",
			5520 => x"0405577b",
			5521 => x"fea4577b",
			5522 => x"0f073904",
			5523 => x"ff87577b",
			5524 => x"0283577b",
			5525 => x"01006e08",
			5526 => x"0d060304",
			5527 => x"fc05577b",
			5528 => x"feaf577b",
			5529 => x"040b830c",
			5530 => x"0a026c08",
			5531 => x"040a4904",
			5532 => x"fff1577b",
			5533 => x"fd37577b",
			5534 => x"01aa577b",
			5535 => x"fdda577b",
			5536 => x"06014e3c",
			5537 => x"0e052020",
			5538 => x"09009310",
			5539 => x"0a028808",
			5540 => x"0e050004",
			5541 => x"fdb6577b",
			5542 => x"0000577b",
			5543 => x"0208bb04",
			5544 => x"00ef577b",
			5545 => x"ff4b577b",
			5546 => x"01005e08",
			5547 => x"02088504",
			5548 => x"fc2e577b",
			5549 => x"fde4577b",
			5550 => x"0900aa04",
			5551 => x"0006577b",
			5552 => x"fe79577b",
			5553 => x"0208dd10",
			5554 => x"0d058108",
			5555 => x"0c045b04",
			5556 => x"fabb577b",
			5557 => x"00f3577b",
			5558 => x"06014d04",
			5559 => x"fff3577b",
			5560 => x"fd71577b",
			5561 => x"0c048f04",
			5562 => x"000b577b",
			5563 => x"0003ff04",
			5564 => x"ffdc577b",
			5565 => x"fe0f577b",
			5566 => x"0900b520",
			5567 => x"040c9310",
			5568 => x"0a02b808",
			5569 => x"0d05bd04",
			5570 => x"0031577b",
			5571 => x"0240577b",
			5572 => x"0b04e304",
			5573 => x"00f7577b",
			5574 => x"0254577b",
			5575 => x"09009708",
			5576 => x"0208f004",
			5577 => x"ff45577b",
			5578 => x"01b5577b",
			5579 => x"06016304",
			5580 => x"feb4577b",
			5581 => x"0034577b",
			5582 => x"02094310",
			5583 => x"00047108",
			5584 => x"0c049604",
			5585 => x"ff0e577b",
			5586 => x"0025577b",
			5587 => x"0b04f104",
			5588 => x"00b0577b",
			5589 => x"ff09577b",
			5590 => x"02094908",
			5591 => x"0e05f704",
			5592 => x"0325577b",
			5593 => x"0162577b",
			5594 => x"040d0004",
			5595 => x"00ae577b",
			5596 => x"fe77577b",
			5597 => x"fe77577b",
			5598 => x"07057374",
			5599 => x"040f0268",
			5600 => x"00049630",
			5601 => x"06010710",
			5602 => x"03043504",
			5603 => x"02915885",
			5604 => x"03047f08",
			5605 => x"03046704",
			5606 => x"fece5885",
			5607 => x"00715885",
			5608 => x"fe5d5885",
			5609 => x"0704c110",
			5610 => x"03051b08",
			5611 => x"07047804",
			5612 => x"02a85885",
			5613 => x"009d5885",
			5614 => x"02085904",
			5615 => x"01ac5885",
			5616 => x"00ef5885",
			5617 => x"0704c208",
			5618 => x"0d058e04",
			5619 => x"ff615885",
			5620 => x"fd6f5885",
			5621 => x"06012b04",
			5622 => x"fe865885",
			5623 => x"00cc5885",
			5624 => x"06015a20",
			5625 => x"0a02c910",
			5626 => x"0504e708",
			5627 => x"02080704",
			5628 => x"ffc25885",
			5629 => x"02e75885",
			5630 => x"0f06ca04",
			5631 => x"ff155885",
			5632 => x"00315885",
			5633 => x"040d6e08",
			5634 => x"0803a304",
			5635 => x"01b95885",
			5636 => x"feca5885",
			5637 => x"06014f04",
			5638 => x"03515885",
			5639 => x"00275885",
			5640 => x"0209200c",
			5641 => x"08038d04",
			5642 => x"003d5885",
			5643 => x"0d05e904",
			5644 => x"fe755885",
			5645 => x"00005885",
			5646 => x"0b052208",
			5647 => x"01006e04",
			5648 => x"002a5885",
			5649 => x"04955885",
			5650 => x"fe4b5885",
			5651 => x"040f7008",
			5652 => x"06010e04",
			5653 => x"febb5885",
			5654 => x"00295885",
			5655 => x"fe5a5885",
			5656 => x"0a024510",
			5657 => x"020a180c",
			5658 => x"07058d08",
			5659 => x"0801e404",
			5660 => x"fea35885",
			5661 => x"01965885",
			5662 => x"fe5c5885",
			5663 => x"054a5885",
			5664 => x"fe5a5885",
			5665 => x"0207da54",
			5666 => x"0100794c",
			5667 => x"0e04e238",
			5668 => x"05056420",
			5669 => x"0e045310",
			5670 => x"0d053508",
			5671 => x"0f069004",
			5672 => x"00685a01",
			5673 => x"feba5a01",
			5674 => x"0304df04",
			5675 => x"ffb55a01",
			5676 => x"fe2c5a01",
			5677 => x"08032508",
			5678 => x"06013004",
			5679 => x"00d55a01",
			5680 => x"fefe5a01",
			5681 => x"0704ac04",
			5682 => x"02a45a01",
			5683 => x"012b5a01",
			5684 => x"0f06870c",
			5685 => x"040be408",
			5686 => x"02077704",
			5687 => x"fef85a01",
			5688 => x"014c5a01",
			5689 => x"fe5b5a01",
			5690 => x"05056704",
			5691 => x"fd775a01",
			5692 => x"0d057504",
			5693 => x"00895a01",
			5694 => x"feac5a01",
			5695 => x"0a022b0c",
			5696 => x"04095908",
			5697 => x"01006104",
			5698 => x"00005a01",
			5699 => x"00ff5a01",
			5700 => x"fe8b5a01",
			5701 => x"0f06f904",
			5702 => x"01f15a01",
			5703 => x"00d95a01",
			5704 => x"0f075704",
			5705 => x"fdb95a01",
			5706 => x"00005a01",
			5707 => x"0207df14",
			5708 => x"0704aa0c",
			5709 => x"0e045308",
			5710 => x"07046c04",
			5711 => x"01315a01",
			5712 => x"fe335a01",
			5713 => x"00875a01",
			5714 => x"05060804",
			5715 => x"fdef5a01",
			5716 => x"00005a01",
			5717 => x"03048f28",
			5718 => x"040d000c",
			5719 => x"06013108",
			5720 => x"01004104",
			5721 => x"016b5a01",
			5722 => x"fe885a01",
			5723 => x"fe525a01",
			5724 => x"07049110",
			5725 => x"02084d08",
			5726 => x"03046f04",
			5727 => x"00635a01",
			5728 => x"02215a01",
			5729 => x"0f068704",
			5730 => x"001b5a01",
			5731 => x"fe665a01",
			5732 => x"02085404",
			5733 => x"fe515a01",
			5734 => x"0e03a604",
			5735 => x"00005a01",
			5736 => x"00ee5a01",
			5737 => x"0d050d14",
			5738 => x"07049410",
			5739 => x"0f070f08",
			5740 => x"040be404",
			5741 => x"ffe25a01",
			5742 => x"01955a01",
			5743 => x"02089f04",
			5744 => x"fe345a01",
			5745 => x"00ba5a01",
			5746 => x"fe965a01",
			5747 => x"0f067a0c",
			5748 => x"0f067408",
			5749 => x"0d054004",
			5750 => x"fe4b5a01",
			5751 => x"01c75a01",
			5752 => x"02f85a01",
			5753 => x"03050d08",
			5754 => x"0f06ed04",
			5755 => x"ffee5a01",
			5756 => x"ff445a01",
			5757 => x"09008f04",
			5758 => x"006b5a01",
			5759 => x"fff25a01",
			5760 => x"0c050b68",
			5761 => x"040fc664",
			5762 => x"07050340",
			5763 => x"0e04f720",
			5764 => x"0f070510",
			5765 => x"0d058308",
			5766 => x"03051b04",
			5767 => x"007c5b25",
			5768 => x"013c5b25",
			5769 => x"01007104",
			5770 => x"fed85b25",
			5771 => x"02aa5b25",
			5772 => x"0a027208",
			5773 => x"05057604",
			5774 => x"fe915b25",
			5775 => x"00cd5b25",
			5776 => x"00042104",
			5777 => x"02065b25",
			5778 => x"001c5b25",
			5779 => x"0900b510",
			5780 => x"0704c408",
			5781 => x"0704c004",
			5782 => x"00d85b25",
			5783 => x"ffb05b25",
			5784 => x"040c9304",
			5785 => x"01815b25",
			5786 => x"ffcb5b25",
			5787 => x"0e054b08",
			5788 => x"01007104",
			5789 => x"fe275b25",
			5790 => x"ffbc5b25",
			5791 => x"040bbf04",
			5792 => x"00ee5b25",
			5793 => x"00355b25",
			5794 => x"05059504",
			5795 => x"01d35b25",
			5796 => x"0305f910",
			5797 => x"0505cc08",
			5798 => x"0f078704",
			5799 => x"fdd35b25",
			5800 => x"ffac5b25",
			5801 => x"0305d104",
			5802 => x"02c25b25",
			5803 => x"fe815b25",
			5804 => x"06016c08",
			5805 => x"0f082b04",
			5806 => x"00015b25",
			5807 => x"01695b25",
			5808 => x"0a028d04",
			5809 => x"019e5b25",
			5810 => x"feff5b25",
			5811 => x"fe615b25",
			5812 => x"0c054818",
			5813 => x"0b061b14",
			5814 => x"0900dc04",
			5815 => x"fe3f5b25",
			5816 => x"0900e004",
			5817 => x"024e5b25",
			5818 => x"0b05b608",
			5819 => x"0d069f04",
			5820 => x"ff045b25",
			5821 => x"01f65b25",
			5822 => x"fe5d5b25",
			5823 => x"01985b25",
			5824 => x"0c05b810",
			5825 => x"0a024c0c",
			5826 => x"0a023c04",
			5827 => x"fe755b25",
			5828 => x"0c058504",
			5829 => x"ffa85b25",
			5830 => x"024b5b25",
			5831 => x"fe635b25",
			5832 => x"fe605b25",
			5833 => x"0e061e8c",
			5834 => x"0900cd54",
			5835 => x"0b053540",
			5836 => x"01004d20",
			5837 => x"09007710",
			5838 => x"0304c708",
			5839 => x"0f06c504",
			5840 => x"00175ce9",
			5841 => x"ff1c5ce9",
			5842 => x"05052d04",
			5843 => x"014d5ce9",
			5844 => x"fe8a5ce9",
			5845 => x"05052d08",
			5846 => x"0a02a104",
			5847 => x"fed45ce9",
			5848 => x"ff9b5ce9",
			5849 => x"0e045304",
			5850 => x"ff1d5ce9",
			5851 => x"014f5ce9",
			5852 => x"0f068710",
			5853 => x"0f067408",
			5854 => x"0b049e04",
			5855 => x"016e5ce9",
			5856 => x"ffe05ce9",
			5857 => x"0b04b204",
			5858 => x"00625ce9",
			5859 => x"01b95ce9",
			5860 => x"05051008",
			5861 => x"0c047804",
			5862 => x"fff45ce9",
			5863 => x"01ad5ce9",
			5864 => x"0b049d04",
			5865 => x"ff4a5ce9",
			5866 => x"00055ce9",
			5867 => x"0505ea0c",
			5868 => x"0505ce04",
			5869 => x"003e5ce9",
			5870 => x"03060104",
			5871 => x"fff25ce9",
			5872 => x"03335ce9",
			5873 => x"0900c804",
			5874 => x"fe925ce9",
			5875 => x"014f5ce9",
			5876 => x"00044f20",
			5877 => x"01007d04",
			5878 => x"fe025ce9",
			5879 => x"0704f10c",
			5880 => x"0a028e08",
			5881 => x"03062104",
			5882 => x"fd765ce9",
			5883 => x"ffee5ce9",
			5884 => x"006d5ce9",
			5885 => x"0900d608",
			5886 => x"0c050904",
			5887 => x"01905ce9",
			5888 => x"fe505ce9",
			5889 => x"0a029204",
			5890 => x"005b5ce9",
			5891 => x"fefa5ce9",
			5892 => x"0900ec10",
			5893 => x"06017404",
			5894 => x"fe355ce9",
			5895 => x"0505f604",
			5896 => x"feec5ce9",
			5897 => x"01008604",
			5898 => x"01885ce9",
			5899 => x"00005ce9",
			5900 => x"0b058504",
			5901 => x"018e5ce9",
			5902 => x"00005ce9",
			5903 => x"06017944",
			5904 => x"0a02b830",
			5905 => x"0c04d018",
			5906 => x"06016c0c",
			5907 => x"03064804",
			5908 => x"ffa45ce9",
			5909 => x"0c04b404",
			5910 => x"00b85ce9",
			5911 => x"01e55ce9",
			5912 => x"0100a108",
			5913 => x"00042004",
			5914 => x"ff3f5ce9",
			5915 => x"fdb55ce9",
			5916 => x"016a5ce9",
			5917 => x"01008408",
			5918 => x"01008004",
			5919 => x"ff4f5ce9",
			5920 => x"fe0a5ce9",
			5921 => x"06017808",
			5922 => x"0e068d04",
			5923 => x"00a95ce9",
			5924 => x"ff9a5ce9",
			5925 => x"05061604",
			5926 => x"002a5ce9",
			5927 => x"02a75ce9",
			5928 => x"0f085c08",
			5929 => x"0c04d104",
			5930 => x"01545ce9",
			5931 => x"fe405ce9",
			5932 => x"0f08bf08",
			5933 => x"0c050c04",
			5934 => x"02a05ce9",
			5935 => x"ffae5ce9",
			5936 => x"feb65ce9",
			5937 => x"01009208",
			5938 => x"0b054304",
			5939 => x"010b5ce9",
			5940 => x"fea65ce9",
			5941 => x"06018c04",
			5942 => x"fe5a5ce9",
			5943 => x"0f08bf04",
			5944 => x"016c5ce9",
			5945 => x"fead5ce9",
			5946 => x"07051b98",
			5947 => x"0207da48",
			5948 => x"0100431c",
			5949 => x"05051118",
			5950 => x"0505020c",
			5951 => x"0504f208",
			5952 => x"03041f04",
			5953 => x"ff4b5e95",
			5954 => x"01585e95",
			5955 => x"fe435e95",
			5956 => x"03043e04",
			5957 => x"fe9a5e95",
			5958 => x"00044604",
			5959 => x"00895e95",
			5960 => x"032c5e95",
			5961 => x"fe4b5e95",
			5962 => x"09007110",
			5963 => x"07049008",
			5964 => x"03046704",
			5965 => x"ff425e95",
			5966 => x"03105e95",
			5967 => x"05051004",
			5968 => x"03945e95",
			5969 => x"06a25e95",
			5970 => x"06012110",
			5971 => x"0e044b08",
			5972 => x"040a9504",
			5973 => x"01ae5e95",
			5974 => x"fe3c5e95",
			5975 => x"0a024504",
			5976 => x"ff195e95",
			5977 => x"01c05e95",
			5978 => x"03046704",
			5979 => x"fe5a5e95",
			5980 => x"0704aa04",
			5981 => x"014e5e95",
			5982 => x"007b5e95",
			5983 => x"0f087238",
			5984 => x"0900d620",
			5985 => x"0a026510",
			5986 => x"040acf08",
			5987 => x"02083304",
			5988 => x"00bc5e95",
			5989 => x"ff285e95",
			5990 => x"0b04bf04",
			5991 => x"00185e95",
			5992 => x"fe815e95",
			5993 => x"040b0f08",
			5994 => x"0003ea04",
			5995 => x"00215e95",
			5996 => x"01625e95",
			5997 => x"0a028304",
			5998 => x"ffe05e95",
			5999 => x"00405e95",
			6000 => x"0004200c",
			6001 => x"0f078704",
			6002 => x"fe0e5e95",
			6003 => x"06016204",
			6004 => x"01395e95",
			6005 => x"ff805e95",
			6006 => x"0a029d04",
			6007 => x"fcaf5e95",
			6008 => x"0e060f04",
			6009 => x"fde25e95",
			6010 => x"ff545e95",
			6011 => x"03075414",
			6012 => x"09010f10",
			6013 => x"08036508",
			6014 => x"040b7804",
			6015 => x"01265e95",
			6016 => x"fe235e95",
			6017 => x"040c7204",
			6018 => x"034a5e95",
			6019 => x"ff9c5e95",
			6020 => x"06355e95",
			6021 => x"fe8c5e95",
			6022 => x"03067810",
			6023 => x"0f08390c",
			6024 => x"0b055204",
			6025 => x"fdd25e95",
			6026 => x"0b055404",
			6027 => x"00005e95",
			6028 => x"fe615e95",
			6029 => x"02455e95",
			6030 => x"0900f718",
			6031 => x"01007d04",
			6032 => x"fe7b5e95",
			6033 => x"02091108",
			6034 => x"0208d404",
			6035 => x"01f45e95",
			6036 => x"fe495e95",
			6037 => x"0f088b08",
			6038 => x"06017404",
			6039 => x"03345e95",
			6040 => x"ff475e95",
			6041 => x"feac5e95",
			6042 => x"07064014",
			6043 => x"05080410",
			6044 => x"0b059908",
			6045 => x"040a1504",
			6046 => x"00c75e95",
			6047 => x"fe275e95",
			6048 => x"07054504",
			6049 => x"024e5e95",
			6050 => x"ff3c5e95",
			6051 => x"02495e95",
			6052 => x"fe6a5e95",
			6053 => x"0c054578",
			6054 => x"040fc674",
			6055 => x"0c04b23c",
			6056 => x"0c04961c",
			6057 => x"0c049410",
			6058 => x"0a029308",
			6059 => x"02084d04",
			6060 => x"00705fd1",
			6061 => x"ff9c5fd1",
			6062 => x"040c0a04",
			6063 => x"015c5fd1",
			6064 => x"00715fd1",
			6065 => x"040d6e08",
			6066 => x"040a5b04",
			6067 => x"fc755fd1",
			6068 => x"ffbd5fd1",
			6069 => x"03555fd1",
			6070 => x"0c049710",
			6071 => x"03051008",
			6072 => x"0d053f04",
			6073 => x"01b55fd1",
			6074 => x"febb5fd1",
			6075 => x"0d057604",
			6076 => x"02435fd1",
			6077 => x"01105fd1",
			6078 => x"040c7208",
			6079 => x"08037f04",
			6080 => x"00905fd1",
			6081 => x"02ca5fd1",
			6082 => x"01004f04",
			6083 => x"00ee5fd1",
			6084 => x"fee15fd1",
			6085 => x"0c04b318",
			6086 => x"0d05b610",
			6087 => x"08033608",
			6088 => x"0207ed04",
			6089 => x"00005fd1",
			6090 => x"fd825fd1",
			6091 => x"05059204",
			6092 => x"ff215fd1",
			6093 => x"01db5fd1",
			6094 => x"0d05cf04",
			6095 => x"fd2c5fd1",
			6096 => x"fe5b5fd1",
			6097 => x"0e050710",
			6098 => x"0f069f08",
			6099 => x"0e043604",
			6100 => x"ff3d5fd1",
			6101 => x"024b5fd1",
			6102 => x"05053a04",
			6103 => x"013d5fd1",
			6104 => x"ff5c5fd1",
			6105 => x"0900ab08",
			6106 => x"0c04e904",
			6107 => x"016b5fd1",
			6108 => x"fe035fd1",
			6109 => x"040c1804",
			6110 => x"00595fd1",
			6111 => x"ffba5fd1",
			6112 => x"fe675fd1",
			6113 => x"0c05b824",
			6114 => x"07061318",
			6115 => x"0705fc10",
			6116 => x"0705730c",
			6117 => x"07056104",
			6118 => x"fed55fd1",
			6119 => x"0c054c04",
			6120 => x"006b5fd1",
			6121 => x"00005fd1",
			6122 => x"fe695fd1",
			6123 => x"0c059b04",
			6124 => x"02585fd1",
			6125 => x"feb45fd1",
			6126 => x"07061504",
			6127 => x"06235fd1",
			6128 => x"040abb04",
			6129 => x"ff2e5fd1",
			6130 => x"016b5fd1",
			6131 => x"fe645fd1",
			6132 => x"0c04f19c",
			6133 => x"040c605c",
			6134 => x"0304d82c",
			6135 => x"0b049014",
			6136 => x"040ac904",
			6137 => x"063c6175",
			6138 => x"03045e08",
			6139 => x"0b048d04",
			6140 => x"fe306175",
			6141 => x"00006175",
			6142 => x"09006204",
			6143 => x"05b76175",
			6144 => x"00c86175",
			6145 => x"0e04360c",
			6146 => x"0c045a04",
			6147 => x"02206175",
			6148 => x"00046304",
			6149 => x"ff696175",
			6150 => x"fe606175",
			6151 => x"0a026c04",
			6152 => x"fe386175",
			6153 => x"0f068a04",
			6154 => x"05966175",
			6155 => x"006b6175",
			6156 => x"0306c51c",
			6157 => x"0a02450c",
			6158 => x"06013908",
			6159 => x"06010e04",
			6160 => x"fe536175",
			6161 => x"00336175",
			6162 => x"045d6175",
			6163 => x"040b4a08",
			6164 => x"03051b04",
			6165 => x"01206175",
			6166 => x"03476175",
			6167 => x"08031704",
			6168 => x"ffa76175",
			6169 => x"022b6175",
			6170 => x"0003b704",
			6171 => x"03fc6175",
			6172 => x"00044f08",
			6173 => x"0b058504",
			6174 => x"fe996175",
			6175 => x"01656175",
			6176 => x"01009b04",
			6177 => x"02de6175",
			6178 => x"fe6b6175",
			6179 => x"09004204",
			6180 => x"fe466175",
			6181 => x"0208bb1c",
			6182 => x"0b047d0c",
			6183 => x"06012b04",
			6184 => x"fe626175",
			6185 => x"0207d104",
			6186 => x"003a6175",
			6187 => x"047a6175",
			6188 => x"0004a708",
			6189 => x"08039304",
			6190 => x"00ba6175",
			6191 => x"04e26175",
			6192 => x"040d5504",
			6193 => x"ff616175",
			6194 => x"011d6175",
			6195 => x"040cd810",
			6196 => x"0a02c108",
			6197 => x"0c047504",
			6198 => x"02096175",
			6199 => x"fef66175",
			6200 => x"0900dc04",
			6201 => x"01d66175",
			6202 => x"fe396175",
			6203 => x"0e056108",
			6204 => x"0a033404",
			6205 => x"fe716175",
			6206 => x"00006175",
			6207 => x"03060904",
			6208 => x"02d56175",
			6209 => x"fe7e6175",
			6210 => x"0c052a2c",
			6211 => x"0f07ce0c",
			6212 => x"0305d108",
			6213 => x"0505df04",
			6214 => x"00a46175",
			6215 => x"fe6b6175",
			6216 => x"fe576175",
			6217 => x"02099518",
			6218 => x"0b059910",
			6219 => x"01009508",
			6220 => x"0b057404",
			6221 => x"000b6175",
			6222 => x"03fc6175",
			6223 => x"0b057604",
			6224 => x"ffac6175",
			6225 => x"fe336175",
			6226 => x"05069104",
			6227 => x"03c86175",
			6228 => x"00ad6175",
			6229 => x"0a029b04",
			6230 => x"010f6175",
			6231 => x"fe546175",
			6232 => x"0c059908",
			6233 => x"0c058504",
			6234 => x"fe5c6175",
			6235 => x"ff766175",
			6236 => x"fe456175",
			6237 => x"07054588",
			6238 => x"01003208",
			6239 => x"06014604",
			6240 => x"fe5762d9",
			6241 => x"012162d9",
			6242 => x"09008240",
			6243 => x"0304d820",
			6244 => x"09007e10",
			6245 => x"03049708",
			6246 => x"0a024c04",
			6247 => x"031862d9",
			6248 => x"fff362d9",
			6249 => x"09007504",
			6250 => x"01af62d9",
			6251 => x"005562d9",
			6252 => x"01004f08",
			6253 => x"05050f04",
			6254 => x"ff5c62d9",
			6255 => x"fe1b62d9",
			6256 => x"01005004",
			6257 => x"037f62d9",
			6258 => x"ffdd62d9",
			6259 => x"0f06ed10",
			6260 => x"08030a08",
			6261 => x"0b049e04",
			6262 => x"fe5462d9",
			6263 => x"000d62d9",
			6264 => x"0a02b004",
			6265 => x"028d62d9",
			6266 => x"058562d9",
			6267 => x"0304f708",
			6268 => x"09007504",
			6269 => x"01fe62d9",
			6270 => x"fed062d9",
			6271 => x"07049404",
			6272 => x"01f462d9",
			6273 => x"002f62d9",
			6274 => x"0e04e220",
			6275 => x"09009510",
			6276 => x"03051008",
			6277 => x"0f06ed04",
			6278 => x"003362d9",
			6279 => x"feb462d9",
			6280 => x"0b04d304",
			6281 => x"00a762d9",
			6282 => x"031b62d9",
			6283 => x"0f074908",
			6284 => x"05053d04",
			6285 => x"013062d9",
			6286 => x"ffa862d9",
			6287 => x"040c7904",
			6288 => x"fdbd62d9",
			6289 => x"ff7162d9",
			6290 => x"0900af10",
			6291 => x"0208d008",
			6292 => x"0a02b804",
			6293 => x"00e862d9",
			6294 => x"026962d9",
			6295 => x"08037604",
			6296 => x"ff0962d9",
			6297 => x"009662d9",
			6298 => x"0e057808",
			6299 => x"02085b04",
			6300 => x"003a62d9",
			6301 => x"ff8962d9",
			6302 => x"0900cd04",
			6303 => x"00db62d9",
			6304 => x"000662d9",
			6305 => x"07058d18",
			6306 => x"0b05a704",
			6307 => x"fe5262d9",
			6308 => x"02098e10",
			6309 => x"0208c004",
			6310 => x"fe9362d9",
			6311 => x"040aef04",
			6312 => x"005962d9",
			6313 => x"03076c04",
			6314 => x"00d362d9",
			6315 => x"035662d9",
			6316 => x"fe7562d9",
			6317 => x"0a024c10",
			6318 => x"020a3a0c",
			6319 => x"0705a408",
			6320 => x"0f06c104",
			6321 => x"ffc462d9",
			6322 => x"00bb62d9",
			6323 => x"fe6862d9",
			6324 => x"038962d9",
			6325 => x"fe6562d9",
			6326 => x"0004b8a4",
			6327 => x"0207a140",
			6328 => x"0207671c",
			6329 => x"0003c414",
			6330 => x"0b049e04",
			6331 => x"01e864b5",
			6332 => x"0c049c08",
			6333 => x"00033e04",
			6334 => x"000064b5",
			6335 => x"fecb64b5",
			6336 => x"06011004",
			6337 => x"000064b5",
			6338 => x"017f64b5",
			6339 => x"0c045c04",
			6340 => x"000064b5",
			6341 => x"fe5e64b5",
			6342 => x"0b048e10",
			6343 => x"0d050d0c",
			6344 => x"0f063b08",
			6345 => x"0f060a04",
			6346 => x"019964b5",
			6347 => x"fe8f64b5",
			6348 => x"01b564b5",
			6349 => x"fe5a64b5",
			6350 => x"00046c10",
			6351 => x"0a026708",
			6352 => x"0003cc04",
			6353 => x"002064b5",
			6354 => x"01e764b5",
			6355 => x"0a027504",
			6356 => x"fde864b5",
			6357 => x"007b64b5",
			6358 => x"029c64b5",
			6359 => x"0a02be34",
			6360 => x"05063220",
			6361 => x"0208f210",
			6362 => x"0f07c008",
			6363 => x"0f07ac04",
			6364 => x"fff864b5",
			6365 => x"ff7564b5",
			6366 => x"0e05a404",
			6367 => x"014064b5",
			6368 => x"000b64b5",
			6369 => x"0505b108",
			6370 => x"05053b04",
			6371 => x"01a464b5",
			6372 => x"ff0d64b5",
			6373 => x"0900dc04",
			6374 => x"00ab64b5",
			6375 => x"feda64b5",
			6376 => x"0900f704",
			6377 => x"01e164b5",
			6378 => x"0b056908",
			6379 => x"07050804",
			6380 => x"000064b5",
			6381 => x"020564b5",
			6382 => x"09010f04",
			6383 => x"fed064b5",
			6384 => x"00a264b5",
			6385 => x"05052e14",
			6386 => x"06014a08",
			6387 => x"0004a704",
			6388 => x"012a64b5",
			6389 => x"fe6764b5",
			6390 => x"05051404",
			6391 => x"000764b5",
			6392 => x"09008404",
			6393 => x"02ed64b5",
			6394 => x"00b164b5",
			6395 => x"0c04920c",
			6396 => x"040c9a08",
			6397 => x"0e04bb04",
			6398 => x"fed164b5",
			6399 => x"011664b5",
			6400 => x"fe3d64b5",
			6401 => x"0900a608",
			6402 => x"03057904",
			6403 => x"005264b5",
			6404 => x"01f564b5",
			6405 => x"06016304",
			6406 => x"ff8264b5",
			6407 => x"005a64b5",
			6408 => x"0208c22c",
			6409 => x"0e04b428",
			6410 => x"0c049418",
			6411 => x"0304d610",
			6412 => x"03049f08",
			6413 => x"0a02d104",
			6414 => x"fe6664b5",
			6415 => x"000a64b5",
			6416 => x"0a02cf04",
			6417 => x"028964b5",
			6418 => x"006b64b5",
			6419 => x"0a02d404",
			6420 => x"fe5064b5",
			6421 => x"000064b5",
			6422 => x"02087c04",
			6423 => x"fe4f64b5",
			6424 => x"02088308",
			6425 => x"06015204",
			6426 => x"000064b5",
			6427 => x"018064b5",
			6428 => x"fe9764b5",
			6429 => x"015464b5",
			6430 => x"05056604",
			6431 => x"fe4764b5",
			6432 => x"0900890c",
			6433 => x"02090c04",
			6434 => x"000064b5",
			6435 => x"00065804",
			6436 => x"01c464b5",
			6437 => x"000064b5",
			6438 => x"0c050708",
			6439 => x"0e062e04",
			6440 => x"fe6d64b5",
			6441 => x"008564b5",
			6442 => x"0305e104",
			6443 => x"017d64b5",
			6444 => x"000064b5",
			6445 => x"09008f88",
			6446 => x"09008e60",
			6447 => x"00044e24",
			6448 => x"09008c14",
			6449 => x"0f074f10",
			6450 => x"040bd808",
			6451 => x"00043e04",
			6452 => x"007166a1",
			6453 => x"ff7d66a1",
			6454 => x"0f072504",
			6455 => x"015966a1",
			6456 => x"fe4e66a1",
			6457 => x"fdeb66a1",
			6458 => x"00043f0c",
			6459 => x"02082f08",
			6460 => x"06013004",
			6461 => x"fe3066a1",
			6462 => x"003e66a1",
			6463 => x"fd6d66a1",
			6464 => x"009666a1",
			6465 => x"03052520",
			6466 => x"0f06ed10",
			6467 => x"0304d808",
			6468 => x"08035504",
			6469 => x"ff3366a1",
			6470 => x"fff766a1",
			6471 => x"0f06b204",
			6472 => x"01e166a1",
			6473 => x"002466a1",
			6474 => x"0704a508",
			6475 => x"02085b04",
			6476 => x"fe7c66a1",
			6477 => x"ffe366a1",
			6478 => x"0c047b04",
			6479 => x"ff6266a1",
			6480 => x"fe5866a1",
			6481 => x"0c04900c",
			6482 => x"0a02be08",
			6483 => x"09008604",
			6484 => x"015d66a1",
			6485 => x"ffe266a1",
			6486 => x"fe6566a1",
			6487 => x"01005108",
			6488 => x"0c04ad04",
			6489 => x"00c566a1",
			6490 => x"fddc66a1",
			6491 => x"0c049904",
			6492 => x"028466a1",
			6493 => x"00fc66a1",
			6494 => x"0601491c",
			6495 => x"02081108",
			6496 => x"08030804",
			6497 => x"013466a1",
			6498 => x"feac66a1",
			6499 => x"03051f08",
			6500 => x"00046304",
			6501 => x"01f066a1",
			6502 => x"031566a1",
			6503 => x"0d054f08",
			6504 => x"03053704",
			6505 => x"024d66a1",
			6506 => x"006866a1",
			6507 => x"003866a1",
			6508 => x"02084504",
			6509 => x"016c66a1",
			6510 => x"02089d04",
			6511 => x"fdf466a1",
			6512 => x"00d866a1",
			6513 => x"0100550c",
			6514 => x"0c047804",
			6515 => x"ff8666a1",
			6516 => x"00044f04",
			6517 => x"fd1e66a1",
			6518 => x"fe4a66a1",
			6519 => x"03053938",
			6520 => x"0c04ac1c",
			6521 => x"00045f10",
			6522 => x"040adc08",
			6523 => x"040ab204",
			6524 => x"000066a1",
			6525 => x"fd6566a1",
			6526 => x"01005e04",
			6527 => x"ffed66a1",
			6528 => x"00d366a1",
			6529 => x"0d054004",
			6530 => x"007866a1",
			6531 => x"0704d604",
			6532 => x"fecd66a1",
			6533 => x"00ae66a1",
			6534 => x"0f06ca0c",
			6535 => x"0c04af04",
			6536 => x"fdf966a1",
			6537 => x"0c04ce04",
			6538 => x"004e66a1",
			6539 => x"fe3366a1",
			6540 => x"0f071f08",
			6541 => x"03053704",
			6542 => x"fe7e66a1",
			6543 => x"fd5166a1",
			6544 => x"06014d04",
			6545 => x"003b66a1",
			6546 => x"feab66a1",
			6547 => x"03053f10",
			6548 => x"02085908",
			6549 => x"02081504",
			6550 => x"022e66a1",
			6551 => x"fe8a66a1",
			6552 => x"0a02a604",
			6553 => x"02e166a1",
			6554 => x"003166a1",
			6555 => x"0305430c",
			6556 => x"040bd604",
			6557 => x"fd9666a1",
			6558 => x"0e04a504",
			6559 => x"fe2a66a1",
			6560 => x"002166a1",
			6561 => x"0c047408",
			6562 => x"0f073b04",
			6563 => x"003166a1",
			6564 => x"fec366a1",
			6565 => x"01005904",
			6566 => x"00e866a1",
			6567 => x"000066a1",
			6568 => x"0c050b70",
			6569 => x"040f706c",
			6570 => x"0004963c",
			6571 => x"0704a71c",
			6572 => x"05052d10",
			6573 => x"0c047608",
			6574 => x"09005504",
			6575 => x"fe6b680d",
			6576 => x"015c680d",
			6577 => x"040c9a04",
			6578 => x"004b680d",
			6579 => x"0321680d",
			6580 => x"02077704",
			6581 => x"fe4b680d",
			6582 => x"09008004",
			6583 => x"0330680d",
			6584 => x"016b680d",
			6585 => x"06012510",
			6586 => x"0b04ce08",
			6587 => x"040b0204",
			6588 => x"0173680d",
			6589 => x"fe71680d",
			6590 => x"09010604",
			6591 => x"fe7c680d",
			6592 => x"02db680d",
			6593 => x"040b9708",
			6594 => x"06013a04",
			6595 => x"007c680d",
			6596 => x"0132680d",
			6597 => x"0a028d04",
			6598 => x"ffbc680d",
			6599 => x"00a5680d",
			6600 => x"06015a14",
			6601 => x"06015710",
			6602 => x"0004e908",
			6603 => x"03048f04",
			6604 => x"ff6d680d",
			6605 => x"0056680d",
			6606 => x"0f069904",
			6607 => x"027d680d",
			6608 => x"0000680d",
			6609 => x"043f680d",
			6610 => x"02092010",
			6611 => x"0004a308",
			6612 => x"01006a04",
			6613 => x"01e3680d",
			6614 => x"fe3b680d",
			6615 => x"0d05dc04",
			6616 => x"fe78680d",
			6617 => x"0022680d",
			6618 => x"040ce104",
			6619 => x"0301680d",
			6620 => x"0f07fe04",
			6621 => x"fe59680d",
			6622 => x"0030680d",
			6623 => x"fe5c680d",
			6624 => x"0c054528",
			6625 => x"03064804",
			6626 => x"fe40680d",
			6627 => x"02094914",
			6628 => x"040b8010",
			6629 => x"09010f08",
			6630 => x"0c052804",
			6631 => x"fe3c680d",
			6632 => x"0000680d",
			6633 => x"0b05b704",
			6634 => x"01be680d",
			6635 => x"fe6c680d",
			6636 => x"02f8680d",
			6637 => x"0d07550c",
			6638 => x"06017804",
			6639 => x"fe42680d",
			6640 => x"0100a304",
			6641 => x"007d680d",
			6642 => x"fe82680d",
			6643 => x"013e680d",
			6644 => x"0c05b81c",
			6645 => x"07063d18",
			6646 => x"0705730c",
			6647 => x"00043108",
			6648 => x"07056104",
			6649 => x"feef680d",
			6650 => x"0154680d",
			6651 => x"fe7a680d",
			6652 => x"0705fc04",
			6653 => x"fe5e680d",
			6654 => x"0705fd04",
			6655 => x"00dd680d",
			6656 => x"fe72680d",
			6657 => x"024e680d",
			6658 => x"fe5c680d",
			6659 => x"0c0543ac",
			6660 => x"09008f64",
			6661 => x"0c04963c",
			6662 => x"0207df1c",
			6663 => x"0e045310",
			6664 => x"0704aa08",
			6665 => x"03040e04",
			6666 => x"ff456979",
			6667 => x"00a96979",
			6668 => x"0a029604",
			6669 => x"fe386979",
			6670 => x"01666979",
			6671 => x"00041008",
			6672 => x"0b04af04",
			6673 => x"ffa56979",
			6674 => x"01b26979",
			6675 => x"037f6979",
			6676 => x"0a028310",
			6677 => x"02084d08",
			6678 => x"08033004",
			6679 => x"00436979",
			6680 => x"ff0c6979",
			6681 => x"00044304",
			6682 => x"fdd16979",
			6683 => x"01516979",
			6684 => x"040baa08",
			6685 => x"02084604",
			6686 => x"02846979",
			6687 => x"00256979",
			6688 => x"0d056804",
			6689 => x"00286979",
			6690 => x"02746979",
			6691 => x"01005a20",
			6692 => x"0e047110",
			6693 => x"0d053408",
			6694 => x"0b04a104",
			6695 => x"003e6979",
			6696 => x"03776979",
			6697 => x"02083004",
			6698 => x"00336979",
			6699 => x"feaf6979",
			6700 => x"02089008",
			6701 => x"0a02c304",
			6702 => x"018e6979",
			6703 => x"059b6979",
			6704 => x"0704ac04",
			6705 => x"00d86979",
			6706 => x"fe086979",
			6707 => x"0c04af04",
			6708 => x"01626979",
			6709 => x"05106979",
			6710 => x"0100550c",
			6711 => x"0208a408",
			6712 => x"0704a804",
			6713 => x"fe5b6979",
			6714 => x"fcb46979",
			6715 => x"ff626979",
			6716 => x"0305791c",
			6717 => x"0900a910",
			6718 => x"0704c408",
			6719 => x"0704a704",
			6720 => x"00516979",
			6721 => x"ffaa6979",
			6722 => x"03050d04",
			6723 => x"fe2b6979",
			6724 => x"00be6979",
			6725 => x"0e052608",
			6726 => x"0b04d304",
			6727 => x"fdf26979",
			6728 => x"ffc26979",
			6729 => x"fbbe6979",
			6730 => x"0900a410",
			6731 => x"0c04b408",
			6732 => x"0208d604",
			6733 => x"01526979",
			6734 => x"ff716979",
			6735 => x"01006404",
			6736 => x"01c56979",
			6737 => x"04536979",
			6738 => x"03058708",
			6739 => x"0900b504",
			6740 => x"01646979",
			6741 => x"fde96979",
			6742 => x"0e052004",
			6743 => x"ff696979",
			6744 => x"002e6979",
			6745 => x"0c05b808",
			6746 => x"0507d904",
			6747 => x"fe716979",
			6748 => x"023e6979",
			6749 => x"fe6a6979",
			6750 => x"0c0543bc",
			6751 => x"0900a95c",
			6752 => x"0704ad34",
			6753 => x"0704aa18",
			6754 => x"0c04b410",
			6755 => x"02080208",
			6756 => x"00048a04",
			6757 => x"00996b05",
			6758 => x"ff726b05",
			6759 => x"0a027004",
			6760 => x"feda6b05",
			6761 => x"00146b05",
			6762 => x"040c2604",
			6763 => x"ffc76b05",
			6764 => x"03306b05",
			6765 => x"0a02b110",
			6766 => x"0c049808",
			6767 => x"0f06d904",
			6768 => x"feff6b05",
			6769 => x"fddf6b05",
			6770 => x"0207eb04",
			6771 => x"fdc96b05",
			6772 => x"00c86b05",
			6773 => x"0c047904",
			6774 => x"fe426b05",
			6775 => x"05054804",
			6776 => x"01656b05",
			6777 => x"ffa66b05",
			6778 => x"0a02490c",
			6779 => x"01006508",
			6780 => x"0704bd04",
			6781 => x"fef26b05",
			6782 => x"fdf06b05",
			6783 => x"01446b05",
			6784 => x"040ba410",
			6785 => x"0c047808",
			6786 => x"0e04d304",
			6787 => x"feef6b05",
			6788 => x"00e86b05",
			6789 => x"09009b04",
			6790 => x"01a66b05",
			6791 => x"00b96b05",
			6792 => x"0d051a04",
			6793 => x"04606b05",
			6794 => x"0e04c304",
			6795 => x"ffe06b05",
			6796 => x"00816b05",
			6797 => x"0e054b30",
			6798 => x"01006810",
			6799 => x"040b3c04",
			6800 => x"fccd6b05",
			6801 => x"02085904",
			6802 => x"01136b05",
			6803 => x"040bd604",
			6804 => x"fced6b05",
			6805 => x"fecf6b05",
			6806 => x"0d05c210",
			6807 => x"0f076b08",
			6808 => x"0e051604",
			6809 => x"ffa16b05",
			6810 => x"00bc6b05",
			6811 => x"08034d04",
			6812 => x"fe266b05",
			6813 => x"fff76b05",
			6814 => x"0c04ee08",
			6815 => x"0f079104",
			6816 => x"fe156b05",
			6817 => x"00006b05",
			6818 => x"08036b04",
			6819 => x"fee86b05",
			6820 => x"04126b05",
			6821 => x"0900af18",
			6822 => x"0208e90c",
			6823 => x"0f07b908",
			6824 => x"0c04ae04",
			6825 => x"01ee6b05",
			6826 => x"00746b05",
			6827 => x"02bc6b05",
			6828 => x"08037704",
			6829 => x"fe396b05",
			6830 => x"0b04f104",
			6831 => x"ffae6b05",
			6832 => x"01ed6b05",
			6833 => x"0f072b0c",
			6834 => x"0c04af04",
			6835 => x"00f06b05",
			6836 => x"0f071d04",
			6837 => x"fef16b05",
			6838 => x"fb286b05",
			6839 => x"0f073904",
			6840 => x"01fe6b05",
			6841 => x"0e057104",
			6842 => x"ff8b6b05",
			6843 => x"00286b05",
			6844 => x"0a024c08",
			6845 => x"020a3a04",
			6846 => x"fe846b05",
			6847 => x"01be6b05",
			6848 => x"fe6e6b05",
			6849 => x"0c0543c0",
			6850 => x"0f06e350",
			6851 => x"03052528",
			6852 => x"09009718",
			6853 => x"01005e10",
			6854 => x"09008d08",
			6855 => x"0304d804",
			6856 => x"00186c99",
			6857 => x"00d26c99",
			6858 => x"0d054d04",
			6859 => x"008b6c99",
			6860 => x"ff3f6c99",
			6861 => x"0c049504",
			6862 => x"03c26c99",
			6863 => x"00786c99",
			6864 => x"0e047804",
			6865 => x"fdf56c99",
			6866 => x"02081108",
			6867 => x"0d057304",
			6868 => x"017d6c99",
			6869 => x"fe9b6c99",
			6870 => x"fd9e6c99",
			6871 => x"0d05ab1c",
			6872 => x"040bb20c",
			6873 => x"08033908",
			6874 => x"0f069f04",
			6875 => x"021b6c99",
			6876 => x"00b56c99",
			6877 => x"fd096c99",
			6878 => x"02081d08",
			6879 => x"0f06d004",
			6880 => x"039f6c99",
			6881 => x"02056c99",
			6882 => x"0e048f04",
			6883 => x"ff446c99",
			6884 => x"03036c99",
			6885 => x"0e052d04",
			6886 => x"fda36c99",
			6887 => x"0600fb04",
			6888 => x"ff0a6c99",
			6889 => x"02636c99",
			6890 => x"06014140",
			6891 => x"0305b920",
			6892 => x"0e051610",
			6893 => x"08032108",
			6894 => x"03053304",
			6895 => x"fdf46c99",
			6896 => x"ff776c99",
			6897 => x"0e050004",
			6898 => x"000d6c99",
			6899 => x"fe126c99",
			6900 => x"0d05a708",
			6901 => x"08032004",
			6902 => x"01cd6c99",
			6903 => x"ffe26c99",
			6904 => x"0f073b04",
			6905 => x"fd4c6c99",
			6906 => x"ff3f6c99",
			6907 => x"0e058e10",
			6908 => x"02083d08",
			6909 => x"02081504",
			6910 => x"fdb66c99",
			6911 => x"00cd6c99",
			6912 => x"0900af04",
			6913 => x"ff966c99",
			6914 => x"fd606c99",
			6915 => x"0a024708",
			6916 => x"040a0104",
			6917 => x"ffef6c99",
			6918 => x"fd2d6c99",
			6919 => x"02088904",
			6920 => x"01bb6c99",
			6921 => x"ff1e6c99",
			6922 => x"0c045b14",
			6923 => x"06014608",
			6924 => x"02086e04",
			6925 => x"fe346c99",
			6926 => x"00856c99",
			6927 => x"02087c04",
			6928 => x"ffa06c99",
			6929 => x"0d054204",
			6930 => x"fe696c99",
			6931 => x"fc996c99",
			6932 => x"0c04720c",
			6933 => x"0208ab08",
			6934 => x"0a02b004",
			6935 => x"016e6c99",
			6936 => x"ff326c99",
			6937 => x"02fa6c99",
			6938 => x"0802fb08",
			6939 => x"0208b404",
			6940 => x"01e86c99",
			6941 => x"ffc06c99",
			6942 => x"0003cc04",
			6943 => x"fe656c99",
			6944 => x"001f6c99",
			6945 => x"0a024c08",
			6946 => x"020a3a04",
			6947 => x"fe896c99",
			6948 => x"01976c99",
			6949 => x"fe706c99",
			6950 => x"0803a39c",
			6951 => x"0a02d178",
			6952 => x"09007e3c",
			6953 => x"05051f20",
			6954 => x"00044b10",
			6955 => x"07047808",
			6956 => x"0504e704",
			6957 => x"01716e55",
			6958 => x"fe146e55",
			6959 => x"0a028204",
			6960 => x"004d6e55",
			6961 => x"01796e55",
			6962 => x"00045208",
			6963 => x"0c047804",
			6964 => x"fe526e55",
			6965 => x"ff8c6e55",
			6966 => x"0e03f104",
			6967 => x"ff9e6e55",
			6968 => x"003a6e55",
			6969 => x"0a028310",
			6970 => x"09007708",
			6971 => x"09007304",
			6972 => x"febb6e55",
			6973 => x"016b6e55",
			6974 => x"0e044b04",
			6975 => x"fe296e55",
			6976 => x"001b6e55",
			6977 => x"01004504",
			6978 => x"ff716e55",
			6979 => x"00046b04",
			6980 => x"02946e55",
			6981 => x"010b6e55",
			6982 => x"0100511c",
			6983 => x"05052d10",
			6984 => x"05051108",
			6985 => x"06014104",
			6986 => x"ff896e55",
			6987 => x"01826e55",
			6988 => x"0f070904",
			6989 => x"ff5f6e55",
			6990 => x"fe406e55",
			6991 => x"07048f04",
			6992 => x"02066e55",
			6993 => x"0e045304",
			6994 => x"fecd6e55",
			6995 => x"00486e55",
			6996 => x"09008b10",
			6997 => x"07049708",
			6998 => x"09008a04",
			6999 => x"000f6e55",
			7000 => x"fdbb6e55",
			7001 => x"09008a04",
			7002 => x"00656e55",
			7003 => x"01d76e55",
			7004 => x"0e04a908",
			7005 => x"06013104",
			7006 => x"ff1f6e55",
			7007 => x"ffde6e55",
			7008 => x"0a02c404",
			7009 => x"fffe6e55",
			7010 => x"009a6e55",
			7011 => x"09008a04",
			7012 => x"032a6e55",
			7013 => x"0b04e208",
			7014 => x"0004b004",
			7015 => x"00726e55",
			7016 => x"fe626e55",
			7017 => x"0505a108",
			7018 => x"0e051d04",
			7019 => x"00006e55",
			7020 => x"028c6e55",
			7021 => x"0f082b08",
			7022 => x"06017404",
			7023 => x"fe686e55",
			7024 => x"00006e55",
			7025 => x"01008604",
			7026 => x"021f6e55",
			7027 => x"fe836e55",
			7028 => x"02093040",
			7029 => x"0208f22c",
			7030 => x"0f068a18",
			7031 => x"0e03cb10",
			7032 => x"0c045a08",
			7033 => x"0207d704",
			7034 => x"00006e55",
			7035 => x"016a6e55",
			7036 => x"06014704",
			7037 => x"ff9e6e55",
			7038 => x"fe3e6e55",
			7039 => x"01005004",
			7040 => x"01436e55",
			7041 => x"fe8f6e55",
			7042 => x"0704a608",
			7043 => x"02088304",
			7044 => x"fdf56e55",
			7045 => x"ff816e55",
			7046 => x"0b04bf08",
			7047 => x"0d054104",
			7048 => x"fef56e55",
			7049 => x"00f66e55",
			7050 => x"fe6f6e55",
			7051 => x"05056604",
			7052 => x"fea76e55",
			7053 => x"06015308",
			7054 => x"0705b804",
			7055 => x"03916e55",
			7056 => x"00006e55",
			7057 => x"06017004",
			7058 => x"ff476e55",
			7059 => x"01986e55",
			7060 => x"fe4d6e55",
			7061 => x"0c050dc8",
			7062 => x"0207da58",
			7063 => x"0100432c",
			7064 => x"0c04761c",
			7065 => x"07046c0c",
			7066 => x"0b045e08",
			7067 => x"01001d04",
			7068 => x"febc7021",
			7069 => x"003c7021",
			7070 => x"fe0b7021",
			7071 => x"07047a08",
			7072 => x"0b047e04",
			7073 => x"02c67021",
			7074 => x"ff6e7021",
			7075 => x"0c047404",
			7076 => x"ff807021",
			7077 => x"04077021",
			7078 => x"0704a808",
			7079 => x"07046c04",
			7080 => x"ff797021",
			7081 => x"fe457021",
			7082 => x"0b048f04",
			7083 => x"01f27021",
			7084 => x"fea67021",
			7085 => x"09007110",
			7086 => x"07049008",
			7087 => x"00046704",
			7088 => x"022a7021",
			7089 => x"ff467021",
			7090 => x"05051004",
			7091 => x"02ac7021",
			7092 => x"04567021",
			7093 => x"06012110",
			7094 => x"0d055b08",
			7095 => x"0f06b504",
			7096 => x"ffc67021",
			7097 => x"02017021",
			7098 => x"0409db04",
			7099 => x"ffbc7021",
			7100 => x"fe437021",
			7101 => x"01006f08",
			7102 => x"0d059004",
			7103 => x"00bb7021",
			7104 => x"febe7021",
			7105 => x"02597021",
			7106 => x"0f082b40",
			7107 => x"0d05cf20",
			7108 => x"0c049610",
			7109 => x"0c049408",
			7110 => x"0704c404",
			7111 => x"00197021",
			7112 => x"00c87021",
			7113 => x"0d05ab04",
			7114 => x"ff8d7021",
			7115 => x"fd277021",
			7116 => x"0b04bf08",
			7117 => x"06012b04",
			7118 => x"ff307021",
			7119 => x"01127021",
			7120 => x"0b04c104",
			7121 => x"ff397021",
			7122 => x"00487021",
			7123 => x"040b0910",
			7124 => x"0003d108",
			7125 => x"0409b304",
			7126 => x"01fa7021",
			7127 => x"ff657021",
			7128 => x"0a028b04",
			7129 => x"01757021",
			7130 => x"ffc97021",
			7131 => x"0003fb08",
			7132 => x"02089304",
			7133 => x"fcce7021",
			7134 => x"feb17021",
			7135 => x"0900d604",
			7136 => x"ffcd7021",
			7137 => x"fecb7021",
			7138 => x"0803551c",
			7139 => x"0003f310",
			7140 => x"0c04d408",
			7141 => x"0c04d004",
			7142 => x"011d7021",
			7143 => x"076a7021",
			7144 => x"0b059904",
			7145 => x"fe317021",
			7146 => x"01b47021",
			7147 => x"0c050908",
			7148 => x"040b3604",
			7149 => x"fdef7021",
			7150 => x"ff737021",
			7151 => x"01c67021",
			7152 => x"040d0e10",
			7153 => x"06016608",
			7154 => x"06015f04",
			7155 => x"00c17021",
			7156 => x"02cd7021",
			7157 => x"0f086404",
			7158 => x"fffe7021",
			7159 => x"018f7021",
			7160 => x"fe527021",
			7161 => x"0c05b81c",
			7162 => x"0507d918",
			7163 => x"0c054314",
			7164 => x"02093a0c",
			7165 => x"0208f008",
			7166 => x"0c052804",
			7167 => x"fe597021",
			7168 => x"00007021",
			7169 => x"00f17021",
			7170 => x"0b060604",
			7171 => x"fe5a7021",
			7172 => x"00007021",
			7173 => x"fe747021",
			7174 => x"02147021",
			7175 => x"fe6b7021",
			7176 => x"0c04f1d4",
			7177 => x"0c047968",
			7178 => x"09008a3c",
			7179 => x"03050020",
			7180 => x"0704a810",
			7181 => x"00040208",
			7182 => x"05051404",
			7183 => x"02f67245",
			7184 => x"ff487245",
			7185 => x"0304a704",
			7186 => x"ff9c7245",
			7187 => x"00297245",
			7188 => x"0f067408",
			7189 => x"03049704",
			7190 => x"febc7245",
			7191 => x"017d7245",
			7192 => x"0304d804",
			7193 => x"fe297245",
			7194 => x"ff5a7245",
			7195 => x"0f07010c",
			7196 => x"09007f04",
			7197 => x"00007245",
			7198 => x"0f06de04",
			7199 => x"029a7245",
			7200 => x"019b7245",
			7201 => x"05051e08",
			7202 => x"02089304",
			7203 => x"00187245",
			7204 => x"024d7245",
			7205 => x"0a02a004",
			7206 => x"ff0e7245",
			7207 => x"00aa7245",
			7208 => x"05052d10",
			7209 => x"0b04b00c",
			7210 => x"0e04e208",
			7211 => x"0f071d04",
			7212 => x"ff197245",
			7213 => x"fd517245",
			7214 => x"00577245",
			7215 => x"fce87245",
			7216 => x"0c04720c",
			7217 => x"0a027004",
			7218 => x"fed57245",
			7219 => x"0c045b04",
			7220 => x"ffdd7245",
			7221 => x"02317245",
			7222 => x"0704c408",
			7223 => x"0e050704",
			7224 => x"ff397245",
			7225 => x"001d7245",
			7226 => x"05056804",
			7227 => x"026b7245",
			7228 => x"00007245",
			7229 => x"0c048f2c",
			7230 => x"0a027a14",
			7231 => x"07049304",
			7232 => x"02257245",
			7233 => x"0c047b08",
			7234 => x"0f06e304",
			7235 => x"fdc67245",
			7236 => x"feaf7245",
			7237 => x"09009804",
			7238 => x"ff577245",
			7239 => x"02357245",
			7240 => x"02089810",
			7241 => x"07049008",
			7242 => x"0b047104",
			7243 => x"fe237245",
			7244 => x"00517245",
			7245 => x"09006804",
			7246 => x"febc7245",
			7247 => x"024c7245",
			7248 => x"06014f04",
			7249 => x"ff017245",
			7250 => x"01777245",
			7251 => x"03052520",
			7252 => x"09009510",
			7253 => x"0c049308",
			7254 => x"0c049104",
			7255 => x"ff6c7245",
			7256 => x"00dd7245",
			7257 => x"0f06ca04",
			7258 => x"001c7245",
			7259 => x"ff7d7245",
			7260 => x"08032e08",
			7261 => x"0d057504",
			7262 => x"00b07245",
			7263 => x"fddf7245",
			7264 => x"0f06ed04",
			7265 => x"fde47245",
			7266 => x"00007245",
			7267 => x"09009c10",
			7268 => x"03057908",
			7269 => x"0f074904",
			7270 => x"00a67245",
			7271 => x"ff977245",
			7272 => x"0c049204",
			7273 => x"ffe47245",
			7274 => x"01fe7245",
			7275 => x"0b04c308",
			7276 => x"0c04b304",
			7277 => x"ff377245",
			7278 => x"00ff7245",
			7279 => x"03053904",
			7280 => x"fec67245",
			7281 => x"00147245",
			7282 => x"0f07ce18",
			7283 => x"0506160c",
			7284 => x"0e054408",
			7285 => x"00044604",
			7286 => x"01367245",
			7287 => x"fe757245",
			7288 => x"fdce7245",
			7289 => x"05061908",
			7290 => x"02084404",
			7291 => x"00007245",
			7292 => x"03777245",
			7293 => x"fecc7245",
			7294 => x"0900d308",
			7295 => x"06016204",
			7296 => x"02c77245",
			7297 => x"fe827245",
			7298 => x"0b057404",
			7299 => x"fe5e7245",
			7300 => x"0f088b10",
			7301 => x"0208f008",
			7302 => x"0d069f04",
			7303 => x"feaa7245",
			7304 => x"013b7245",
			7305 => x"0900f704",
			7306 => x"02d67245",
			7307 => x"ff207245",
			7308 => x"0a024108",
			7309 => x"0705bb04",
			7310 => x"012f7245",
			7311 => x"ff2e7245",
			7312 => x"fe7b7245",
			7313 => x"0209abc4",
			7314 => x"0a02b168",
			7315 => x"00048540",
			7316 => x"0207da20",
			7317 => x"06012110",
			7318 => x"0c047508",
			7319 => x"0003e204",
			7320 => x"01b373e1",
			7321 => x"000073e1",
			7322 => x"03050004",
			7323 => x"feb173e1",
			7324 => x"ffd273e1",
			7325 => x"0c047508",
			7326 => x"03047f04",
			7327 => x"fe9173e1",
			7328 => x"001673e1",
			7329 => x"0f065904",
			7330 => x"01ac73e1",
			7331 => x"008073e1",
			7332 => x"01004710",
			7333 => x"0d051a08",
			7334 => x"0b048d04",
			7335 => x"00d173e1",
			7336 => x"ff4973e1",
			7337 => x"07049504",
			7338 => x"01fd73e1",
			7339 => x"fef673e1",
			7340 => x"0304ef08",
			7341 => x"0b048e04",
			7342 => x"004d73e1",
			7343 => x"ff1d73e1",
			7344 => x"0f071f04",
			7345 => x"003573e1",
			7346 => x"ffea73e1",
			7347 => x"0b04a220",
			7348 => x"06013d10",
			7349 => x"040cb608",
			7350 => x"0d052504",
			7351 => x"fe3b73e1",
			7352 => x"ffcb73e1",
			7353 => x"08037304",
			7354 => x"fe3873e1",
			7355 => x"010773e1",
			7356 => x"06014208",
			7357 => x"040c7904",
			7358 => x"ff3c73e1",
			7359 => x"01fa73e1",
			7360 => x"02086204",
			7361 => x"ffa273e1",
			7362 => x"fe0b73e1",
			7363 => x"040cc604",
			7364 => x"fe1873e1",
			7365 => x"ff9773e1",
			7366 => x"040c1224",
			7367 => x"0209351c",
			7368 => x"0b050410",
			7369 => x"0f073b08",
			7370 => x"040bfa04",
			7371 => x"fdd373e1",
			7372 => x"ff2173e1",
			7373 => x"0c04b304",
			7374 => x"015273e1",
			7375 => x"ff3173e1",
			7376 => x"00043a04",
			7377 => x"00ea73e1",
			7378 => x"0f080e04",
			7379 => x"fdec73e1",
			7380 => x"ff7973e1",
			7381 => x"0d062d04",
			7382 => x"028673e1",
			7383 => x"feb873e1",
			7384 => x"0004961c",
			7385 => x"0f06ed0c",
			7386 => x"040c4404",
			7387 => x"ffe273e1",
			7388 => x"0b04b104",
			7389 => x"016a73e1",
			7390 => x"030673e1",
			7391 => x"040c4408",
			7392 => x"040c3804",
			7393 => x"00a973e1",
			7394 => x"021b73e1",
			7395 => x"07051804",
			7396 => x"001073e1",
			7397 => x"019f73e1",
			7398 => x"040c790c",
			7399 => x"08039004",
			7400 => x"fdff73e1",
			7401 => x"0004a304",
			7402 => x"010173e1",
			7403 => x"fe1b73e1",
			7404 => x"0704ab08",
			7405 => x"040cc604",
			7406 => x"ff4373e1",
			7407 => x"001f73e1",
			7408 => x"0d052804",
			7409 => x"035b73e1",
			7410 => x"006773e1",
			7411 => x"0a024c08",
			7412 => x"0c05ba04",
			7413 => x"017573e1",
			7414 => x"ff9673e1",
			7415 => x"fe5973e1",
			7416 => x"0207a154",
			7417 => x"0601464c",
			7418 => x"06012d24",
			7419 => x"08031014",
			7420 => x"02079210",
			7421 => x"05052d08",
			7422 => x"0003e604",
			7423 => x"015375fd",
			7424 => x"ff3c75fd",
			7425 => x"0f06bb04",
			7426 => x"ff0975fd",
			7427 => x"010e75fd",
			7428 => x"019d75fd",
			7429 => x"0b04910c",
			7430 => x"07049508",
			7431 => x"0b046c04",
			7432 => x"01f475fd",
			7433 => x"feda75fd",
			7434 => x"02c375fd",
			7435 => x"fe6375fd",
			7436 => x"0b048010",
			7437 => x"0601360c",
			7438 => x"0f060308",
			7439 => x"0c045a04",
			7440 => x"000075fd",
			7441 => x"025775fd",
			7442 => x"feba75fd",
			7443 => x"fe6e75fd",
			7444 => x"0c047608",
			7445 => x"08036f04",
			7446 => x"ffd675fd",
			7447 => x"017675fd",
			7448 => x"05054908",
			7449 => x"01004504",
			7450 => x"00d075fd",
			7451 => x"025a75fd",
			7452 => x"0c04ac04",
			7453 => x"ff7575fd",
			7454 => x"017775fd",
			7455 => x"0f05da04",
			7456 => x"000075fd",
			7457 => x"fe6b75fd",
			7458 => x"0900826c",
			7459 => x"0304c73c",
			7460 => x"0f06b51c",
			7461 => x"040bb20c",
			7462 => x"09007908",
			7463 => x"08033004",
			7464 => x"009b75fd",
			7465 => x"fe6b75fd",
			7466 => x"fe3e75fd",
			7467 => x"0e041608",
			7468 => x"08034404",
			7469 => x"015075fd",
			7470 => x"ffdf75fd",
			7471 => x"08038204",
			7472 => x"009e75fd",
			7473 => x"023f75fd",
			7474 => x"0b048d10",
			7475 => x"0b047f08",
			7476 => x"01004304",
			7477 => x"000075fd",
			7478 => x"fe5c75fd",
			7479 => x"07047e04",
			7480 => x"02bd75fd",
			7481 => x"ffab75fd",
			7482 => x"09006f08",
			7483 => x"06013d04",
			7484 => x"ff1a75fd",
			7485 => x"014775fd",
			7486 => x"00049204",
			7487 => x"fe1175fd",
			7488 => x"feef75fd",
			7489 => x"0f070518",
			7490 => x"08031508",
			7491 => x"0304f704",
			7492 => x"fe4875fd",
			7493 => x"004e75fd",
			7494 => x"040d1b08",
			7495 => x"040ce104",
			7496 => x"00c675fd",
			7497 => x"027075fd",
			7498 => x"0304d804",
			7499 => x"000075fd",
			7500 => x"fecc75fd",
			7501 => x"08038a10",
			7502 => x"08037408",
			7503 => x"040be904",
			7504 => x"013075fd",
			7505 => x"ff5c75fd",
			7506 => x"07049304",
			7507 => x"01e675fd",
			7508 => x"000775fd",
			7509 => x"0704ad04",
			7510 => x"fe2a75fd",
			7511 => x"000075fd",
			7512 => x"0100572c",
			7513 => x"0505100c",
			7514 => x"0c047504",
			7515 => x"ff5f75fd",
			7516 => x"09008704",
			7517 => x"029f75fd",
			7518 => x"005275fd",
			7519 => x"0c047610",
			7520 => x"02080208",
			7521 => x"040b5604",
			7522 => x"ffb175fd",
			7523 => x"01ec75fd",
			7524 => x"03050004",
			7525 => x"fe5275fd",
			7526 => x"003475fd",
			7527 => x"0c049608",
			7528 => x"0004d204",
			7529 => x"ff3375fd",
			7530 => x"00d075fd",
			7531 => x"0c04b004",
			7532 => x"008675fd",
			7533 => x"ff1175fd",
			7534 => x"0304c704",
			7535 => x"01fc75fd",
			7536 => x"0c047810",
			7537 => x"05053a08",
			7538 => x"05051f04",
			7539 => x"007475fd",
			7540 => x"fe2b75fd",
			7541 => x"08031204",
			7542 => x"fed175fd",
			7543 => x"000b75fd",
			7544 => x"0b04bf08",
			7545 => x"0704c004",
			7546 => x"002f75fd",
			7547 => x"010675fd",
			7548 => x"0304fe04",
			7549 => x"fe9a75fd",
			7550 => x"fff375fd",
			7551 => x"0803a3c8",
			7552 => x"06015f74",
			7553 => x"0c04ac38",
			7554 => x"0c049820",
			7555 => x"0c049410",
			7556 => x"0704c408",
			7557 => x"0704c104",
			7558 => x"00157819",
			7559 => x"fefd7819",
			7560 => x"0208ab04",
			7561 => x"01137819",
			7562 => x"ff707819",
			7563 => x"0c049608",
			7564 => x"040abb04",
			7565 => x"fe2e7819",
			7566 => x"ff967819",
			7567 => x"0d055b04",
			7568 => x"00cf7819",
			7569 => x"ffc57819",
			7570 => x"0704ac0c",
			7571 => x"040c0c08",
			7572 => x"0704a904",
			7573 => x"007b7819",
			7574 => x"027e7819",
			7575 => x"02c87819",
			7576 => x"0e055208",
			7577 => x"02085404",
			7578 => x"00ec7819",
			7579 => x"ff327819",
			7580 => x"01fb7819",
			7581 => x"0c04af1c",
			7582 => x"0208090c",
			7583 => x"01006a08",
			7584 => x"0704bd04",
			7585 => x"00ec7819",
			7586 => x"fe637819",
			7587 => x"01b87819",
			7588 => x"0a026d08",
			7589 => x"01006f04",
			7590 => x"fced7819",
			7591 => x"feef7819",
			7592 => x"040b9d04",
			7593 => x"00647819",
			7594 => x"fefa7819",
			7595 => x"0c04b110",
			7596 => x"0e057108",
			7597 => x"0d058e04",
			7598 => x"00b47819",
			7599 => x"ff477819",
			7600 => x"0d05a704",
			7601 => x"00007819",
			7602 => x"01fa7819",
			7603 => x"0c04b408",
			7604 => x"06012b04",
			7605 => x"fe877819",
			7606 => x"ff9f7819",
			7607 => x"0c04b604",
			7608 => x"00f47819",
			7609 => x"ffea7819",
			7610 => x"0704ec20",
			7611 => x"0d05900c",
			7612 => x"040c5e08",
			7613 => x"03059904",
			7614 => x"00007819",
			7615 => x"01dc7819",
			7616 => x"fe317819",
			7617 => x"0900b508",
			7618 => x"0b04e304",
			7619 => x"00007819",
			7620 => x"02c77819",
			7621 => x"01006f04",
			7622 => x"feaf7819",
			7623 => x"0e05b304",
			7624 => x"00427819",
			7625 => x"01507819",
			7626 => x"0208c214",
			7627 => x"00043d0c",
			7628 => x"03067804",
			7629 => x"01477819",
			7630 => x"0306b904",
			7631 => x"fe0e7819",
			7632 => x"00737819",
			7633 => x"0208b904",
			7634 => x"fdcf7819",
			7635 => x"fee57819",
			7636 => x"06016710",
			7637 => x"0c04ee08",
			7638 => x"0b052004",
			7639 => x"00207819",
			7640 => x"01b27819",
			7641 => x"0e064304",
			7642 => x"fe627819",
			7643 => x"00f77819",
			7644 => x"03068308",
			7645 => x"0004a004",
			7646 => x"fe7a7819",
			7647 => x"00907819",
			7648 => x"0306a504",
			7649 => x"01aa7819",
			7650 => x"ffe67819",
			7651 => x"02093044",
			7652 => x"0208f234",
			7653 => x"0c047518",
			7654 => x"0b048e10",
			7655 => x"09005d08",
			7656 => x"0303bd04",
			7657 => x"fef47819",
			7658 => x"01517819",
			7659 => x"0e03bd04",
			7660 => x"ff517819",
			7661 => x"fe477819",
			7662 => x"0d050f04",
			7663 => x"fefd7819",
			7664 => x"03107819",
			7665 => x"0704a810",
			7666 => x"040e6308",
			7667 => x"0d050004",
			7668 => x"ff397819",
			7669 => x"fe227819",
			7670 => x"06014604",
			7671 => x"00ee7819",
			7672 => x"ff477819",
			7673 => x"0704bd08",
			7674 => x"0803be04",
			7675 => x"00eb7819",
			7676 => x"ff597819",
			7677 => x"fe6c7819",
			7678 => x"0a02db04",
			7679 => x"fec27819",
			7680 => x"0e04bb08",
			7681 => x"02092804",
			7682 => x"ff0e7819",
			7683 => x"00f97819",
			7684 => x"024a7819",
			7685 => x"fe597819",
			7686 => x"0e053bc8",
			7687 => x"0c04935c",
			7688 => x"0c049240",
			7689 => x"040bbf20",
			7690 => x"00042e10",
			7691 => x"040b9108",
			7692 => x"02084604",
			7693 => x"00007aa5",
			7694 => x"fdfc7aa5",
			7695 => x"0e049604",
			7696 => x"02577aa5",
			7697 => x"003f7aa5",
			7698 => x"0e049d08",
			7699 => x"08033604",
			7700 => x"fe877aa5",
			7701 => x"ffc47aa5",
			7702 => x"0a029004",
			7703 => x"fdd87aa5",
			7704 => x"005c7aa5",
			7705 => x"0208ce10",
			7706 => x"00048a08",
			7707 => x"08038104",
			7708 => x"00447aa5",
			7709 => x"02a77aa5",
			7710 => x"0a02ac04",
			7711 => x"fe4f7aa5",
			7712 => x"000a7aa5",
			7713 => x"0c047208",
			7714 => x"040cf504",
			7715 => x"01187aa5",
			7716 => x"fe977aa5",
			7717 => x"05055804",
			7718 => x"fe517aa5",
			7719 => x"fff67aa5",
			7720 => x"0b049d08",
			7721 => x"00047804",
			7722 => x"fe5d7aa5",
			7723 => x"00ce7aa5",
			7724 => x"08031404",
			7725 => x"03c97aa5",
			7726 => x"06014108",
			7727 => x"05053a04",
			7728 => x"023b7aa5",
			7729 => x"ff887aa5",
			7730 => x"06014a04",
			7731 => x"036a7aa5",
			7732 => x"00637aa5",
			7733 => x"0c04962c",
			7734 => x"0a02c61c",
			7735 => x"02080e10",
			7736 => x"0e04a908",
			7737 => x"0a028004",
			7738 => x"fed87aa5",
			7739 => x"00627aa5",
			7740 => x"0802f904",
			7741 => x"ffc57aa5",
			7742 => x"01aa7aa5",
			7743 => x"0d051a04",
			7744 => x"00f17aa5",
			7745 => x"03057704",
			7746 => x"fef37aa5",
			7747 => x"ffed7aa5",
			7748 => x"0704c30c",
			7749 => x"0b04c008",
			7750 => x"0a02dd04",
			7751 => x"01077aa5",
			7752 => x"ff147aa5",
			7753 => x"fe587aa5",
			7754 => x"027b7aa5",
			7755 => x"0b04bf20",
			7756 => x"0b04b110",
			7757 => x"05053c08",
			7758 => x"01005304",
			7759 => x"fff17aa5",
			7760 => x"00fb7aa5",
			7761 => x"0e04b404",
			7762 => x"fe0e7aa5",
			7763 => x"00327aa5",
			7764 => x"0c049908",
			7765 => x"0704ac04",
			7766 => x"01f67aa5",
			7767 => x"038c7aa5",
			7768 => x"03051704",
			7769 => x"ff297aa5",
			7770 => x"01437aa5",
			7771 => x"0b04c110",
			7772 => x"05054908",
			7773 => x"06013904",
			7774 => x"01797aa5",
			7775 => x"fee47aa5",
			7776 => x"0c04b504",
			7777 => x"fe0f7aa5",
			7778 => x"00cb7aa5",
			7779 => x"02084608",
			7780 => x"0d05a904",
			7781 => x"008a7aa5",
			7782 => x"fee07aa5",
			7783 => x"08033304",
			7784 => x"fdef7aa5",
			7785 => x"ffd87aa5",
			7786 => x"0003ea48",
			7787 => x"040adc2c",
			7788 => x"0003d118",
			7789 => x"040abb10",
			7790 => x"06015708",
			7791 => x"0a024104",
			7792 => x"ff4f7aa5",
			7793 => x"00827aa5",
			7794 => x"040a4904",
			7795 => x"fd887aa5",
			7796 => x"00007aa5",
			7797 => x"00036804",
			7798 => x"007f7aa5",
			7799 => x"fd6e7aa5",
			7800 => x"0c04b408",
			7801 => x"0a026c04",
			7802 => x"01ae7aa5",
			7803 => x"fde07aa5",
			7804 => x"0b056308",
			7805 => x"0100a804",
			7806 => x"024e7aa5",
			7807 => x"00007aa5",
			7808 => x"ff237aa5",
			7809 => x"0208bb0c",
			7810 => x"02086204",
			7811 => x"ff267aa5",
			7812 => x"08030204",
			7813 => x"fe457aa5",
			7814 => x"fc657aa5",
			7815 => x"040b420c",
			7816 => x"08032008",
			7817 => x"0003d104",
			7818 => x"ffe77aa5",
			7819 => x"01607aa5",
			7820 => x"fee77aa5",
			7821 => x"fe717aa5",
			7822 => x"08031d14",
			7823 => x"040b560c",
			7824 => x"01006e08",
			7825 => x"0a026d04",
			7826 => x"00907aa5",
			7827 => x"01ef7aa5",
			7828 => x"02337aa5",
			7829 => x"00040804",
			7830 => x"fe1a7aa5",
			7831 => x"02a57aa5",
			7832 => x"03058004",
			7833 => x"fe277aa5",
			7834 => x"02088510",
			7835 => x"06015208",
			7836 => x"0d05a704",
			7837 => x"00a77aa5",
			7838 => x"01a57aa5",
			7839 => x"0c04cb04",
			7840 => x"00fb7aa5",
			7841 => x"fed47aa5",
			7842 => x"06014a08",
			7843 => x"05055904",
			7844 => x"00b57aa5",
			7845 => x"ff017aa5",
			7846 => x"0505a104",
			7847 => x"00a87aa5",
			7848 => x"00267aa5",
			7849 => x"0c059cb8",
			7850 => x"0f070558",
			7851 => x"0304d820",
			7852 => x"0704c11c",
			7853 => x"01005510",
			7854 => x"09007708",
			7855 => x"03048f04",
			7856 => x"ffd67c19",
			7857 => x"00c27c19",
			7858 => x"0207d704",
			7859 => x"00347c19",
			7860 => x"ff497c19",
			7861 => x"0304af04",
			7862 => x"05787c19",
			7863 => x"09008904",
			7864 => x"fe3e7c19",
			7865 => x"00f27c19",
			7866 => x"fe437c19",
			7867 => x"09008c1c",
			7868 => x"03051b10",
			7869 => x"0f06c108",
			7870 => x"0304f704",
			7871 => x"00ed7c19",
			7872 => x"02a37c19",
			7873 => x"02082a04",
			7874 => x"ff677c19",
			7875 => x"00ce7c19",
			7876 => x"01004b04",
			7877 => x"fcf57c19",
			7878 => x"09008b04",
			7879 => x"029a7c19",
			7880 => x"01587c19",
			7881 => x"0100550c",
			7882 => x"0f06e508",
			7883 => x"0f06bb04",
			7884 => x"fe8c7c19",
			7885 => x"fd0e7c19",
			7886 => x"ff3c7c19",
			7887 => x"06012b08",
			7888 => x"05056404",
			7889 => x"ffdf7c19",
			7890 => x"fe907c19",
			7891 => x"00049a04",
			7892 => x"008a7c19",
			7893 => x"fe957c19",
			7894 => x"03053320",
			7895 => x"03052f18",
			7896 => x"03052b10",
			7897 => x"0704a708",
			7898 => x"0a028704",
			7899 => x"fe1f7c19",
			7900 => x"00217c19",
			7901 => x"0c047a04",
			7902 => x"fe387c19",
			7903 => x"ff9c7c19",
			7904 => x"0c049104",
			7905 => x"02107c19",
			7906 => x"ffd07c19",
			7907 => x"0f071f04",
			7908 => x"fede7c19",
			7909 => x"fdb47c19",
			7910 => x"08039020",
			7911 => x"09008c10",
			7912 => x"0f074108",
			7913 => x"07049704",
			7914 => x"00a97c19",
			7915 => x"03327c19",
			7916 => x"06014104",
			7917 => x"fe817c19",
			7918 => x"01417c19",
			7919 => x"03055308",
			7920 => x"09009a04",
			7921 => x"00007c19",
			7922 => x"fec27c19",
			7923 => x"0900a804",
			7924 => x"005a7c19",
			7925 => x"00027c19",
			7926 => x"0a02cc10",
			7927 => x"0c04b008",
			7928 => x"0f076d04",
			7929 => x"06137c19",
			7930 => x"016a7c19",
			7931 => x"040cce04",
			7932 => x"016e7c19",
			7933 => x"fe7d7c19",
			7934 => x"0004a008",
			7935 => x"040cbf04",
			7936 => x"02717c19",
			7937 => x"fe627c19",
			7938 => x"0704aa04",
			7939 => x"01f37c19",
			7940 => x"ff817c19",
			7941 => x"fe747c19",
			7942 => x"0208bbb4",
			7943 => x"06016280",
			7944 => x"06014a40",
			7945 => x"02086c20",
			7946 => x"02086710",
			7947 => x"02086208",
			7948 => x"06013504",
			7949 => x"ffea7f07",
			7950 => x"003a7f07",
			7951 => x"0f06fb04",
			7952 => x"01c97f07",
			7953 => x"fe4a7f07",
			7954 => x"01005a08",
			7955 => x"0d052604",
			7956 => x"03017f07",
			7957 => x"fe807f07",
			7958 => x"01006604",
			7959 => x"02cb7f07",
			7960 => x"008c7f07",
			7961 => x"05058210",
			7962 => x"0208a608",
			7963 => x"0e04a504",
			7964 => x"ff377f07",
			7965 => x"00067f07",
			7966 => x"0a02b104",
			7967 => x"00557f07",
			7968 => x"02887f07",
			7969 => x"0e053b08",
			7970 => x"09009a04",
			7971 => x"017b7f07",
			7972 => x"fe177f07",
			7973 => x"02089f04",
			7974 => x"00147f07",
			7975 => x"fe567f07",
			7976 => x"06014d20",
			7977 => x"0e050710",
			7978 => x"08037c08",
			7979 => x"00048204",
			7980 => x"00657f07",
			7981 => x"fdff7f07",
			7982 => x"00049604",
			7983 => x"03a47f07",
			7984 => x"006f7f07",
			7985 => x"0900b908",
			7986 => x"0a029904",
			7987 => x"01257f07",
			7988 => x"02917f07",
			7989 => x"0f07a604",
			7990 => x"ff8e7f07",
			7991 => x"01f37f07",
			7992 => x"0c04cb10",
			7993 => x"0e056108",
			7994 => x"0900a804",
			7995 => x"008b7f07",
			7996 => x"ff3b7f07",
			7997 => x"06015a04",
			7998 => x"018c7f07",
			7999 => x"ffd67f07",
			8000 => x"0c050708",
			8001 => x"0f077904",
			8002 => x"feea7f07",
			8003 => x"fff07f07",
			8004 => x"0b055404",
			8005 => x"031b7f07",
			8006 => x"fff47f07",
			8007 => x"05060820",
			8008 => x"06016410",
			8009 => x"0208ab0c",
			8010 => x"02083804",
			8011 => x"ffb47f07",
			8012 => x"0e054b04",
			8013 => x"fe597f07",
			8014 => x"fd3a7f07",
			8015 => x"ff7d7f07",
			8016 => x"00041004",
			8017 => x"fd3e7f07",
			8018 => x"00046704",
			8019 => x"01b47f07",
			8020 => x"0b050104",
			8021 => x"00e07f07",
			8022 => x"fe057f07",
			8023 => x"0d064508",
			8024 => x"0c054c04",
			8025 => x"04697f07",
			8026 => x"00007f07",
			8027 => x"0d066a04",
			8028 => x"ffd77f07",
			8029 => x"05066a04",
			8030 => x"019d7f07",
			8031 => x"00007f07",
			8032 => x"06014f58",
			8033 => x"0c047624",
			8034 => x"0a02ac10",
			8035 => x"0208d608",
			8036 => x"08035e04",
			8037 => x"00007f07",
			8038 => x"02ac7f07",
			8039 => x"040c8c04",
			8040 => x"01917f07",
			8041 => x"fe6b7f07",
			8042 => x"0208f90c",
			8043 => x"0b048f08",
			8044 => x"0208c904",
			8045 => x"01d77f07",
			8046 => x"fe9f7f07",
			8047 => x"fda87f07",
			8048 => x"0c045904",
			8049 => x"ff657f07",
			8050 => x"01fb7f07",
			8051 => x"0505a018",
			8052 => x"0900b710",
			8053 => x"0900a408",
			8054 => x"05056804",
			8055 => x"ff147f07",
			8056 => x"01d37f07",
			8057 => x"0e056b04",
			8058 => x"fde97f07",
			8059 => x"ffdd7f07",
			8060 => x"06014d04",
			8061 => x"fe6d7f07",
			8062 => x"fc1f7f07",
			8063 => x"0601490c",
			8064 => x"0100a804",
			8065 => x"fdd17f07",
			8066 => x"0e089604",
			8067 => x"00b97f07",
			8068 => x"ff067f07",
			8069 => x"0f07fe08",
			8070 => x"040c4404",
			8071 => x"01887f07",
			8072 => x"fe3b7f07",
			8073 => x"0208f204",
			8074 => x"fd437f07",
			8075 => x"ffab7f07",
			8076 => x"0900c640",
			8077 => x"040c6620",
			8078 => x"0505af10",
			8079 => x"0900b508",
			8080 => x"05057604",
			8081 => x"ffe57f07",
			8082 => x"020a7f07",
			8083 => x"01006f04",
			8084 => x"fe3e7f07",
			8085 => x"ffe17f07",
			8086 => x"0f07ce08",
			8087 => x"0c04d004",
			8088 => x"01fb7f07",
			8089 => x"ff2f7f07",
			8090 => x"0e05c304",
			8091 => x"030f7f07",
			8092 => x"01ff7f07",
			8093 => x"0b04c010",
			8094 => x"0a02cc08",
			8095 => x"0e04f704",
			8096 => x"00527f07",
			8097 => x"03c47f07",
			8098 => x"0f079d04",
			8099 => x"01247f07",
			8100 => x"fe247f07",
			8101 => x"0b04e308",
			8102 => x"09009504",
			8103 => x"ffda7f07",
			8104 => x"fe1d7f07",
			8105 => x"06015f04",
			8106 => x"fefe7f07",
			8107 => x"00c57f07",
			8108 => x"0c04cc14",
			8109 => x"06015f04",
			8110 => x"fda57f07",
			8111 => x"040c1e08",
			8112 => x"0900cd04",
			8113 => x"01f67f07",
			8114 => x"feff7f07",
			8115 => x"0a02d704",
			8116 => x"fdbd7f07",
			8117 => x"00007f07",
			8118 => x"0c04ce08",
			8119 => x"06017c04",
			8120 => x"02817f07",
			8121 => x"fedd7f07",
			8122 => x"0f07ce08",
			8123 => x"06017404",
			8124 => x"fdbd7f07",
			8125 => x"01787f07",
			8126 => x"06016704",
			8127 => x"00987f07",
			8128 => x"ff6b7f07",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(2792, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(5598, initial_addr_3'length));
	end generate gen_rom_14;

	gen_rom_15: if SELECT_ROM = 15 generate
		bank <= (
			0 => x"00000005",
			1 => x"00000009",
			2 => x"0000000d",
			3 => x"00000011",
			4 => x"00000015",
			5 => x"00000019",
			6 => x"0000001d",
			7 => x"00000021",
			8 => x"00000025",
			9 => x"00000029",
			10 => x"0000002d",
			11 => x"00000031",
			12 => x"00000035",
			13 => x"00000039",
			14 => x"0000003d",
			15 => x"00000041",
			16 => x"00000045",
			17 => x"00000049",
			18 => x"0000004d",
			19 => x"0b05bf04",
			20 => x"00000059",
			21 => x"ffc80059",
			22 => x"07055d04",
			23 => x"00010065",
			24 => x"00000065",
			25 => x"0c046304",
			26 => x"00000071",
			27 => x"fffe0071",
			28 => x"0c046304",
			29 => x"00000085",
			30 => x"0a01e404",
			31 => x"00000085",
			32 => x"ffd40085",
			33 => x"07055d08",
			34 => x"0b043e04",
			35 => x"00000099",
			36 => x"000e0099",
			37 => x"00000099",
			38 => x"06010604",
			39 => x"000000ad",
			40 => x"06015b04",
			41 => x"ffef00ad",
			42 => x"000000ad",
			43 => x"06013608",
			44 => x"0600e104",
			45 => x"000000c1",
			46 => x"000400c1",
			47 => x"000000c1",
			48 => x"01004b08",
			49 => x"09002b04",
			50 => x"000000d5",
			51 => x"000000d5",
			52 => x"ffef00d5",
			53 => x"06011504",
			54 => x"000000e9",
			55 => x"06017c04",
			56 => x"fff300e9",
			57 => x"000000e9",
			58 => x"06012704",
			59 => x"00000105",
			60 => x"06015308",
			61 => x"04100804",
			62 => x"ff8b0105",
			63 => x"00000105",
			64 => x"00000105",
			65 => x"07055d0c",
			66 => x"0f062704",
			67 => x"00000121",
			68 => x"0c052a04",
			69 => x"00340121",
			70 => x"00000121",
			71 => x"00000121",
			72 => x"0601270c",
			73 => x"0600e104",
			74 => x"0000013d",
			75 => x"06011204",
			76 => x"0020013d",
			77 => x"0000013d",
			78 => x"ffd3013d",
			79 => x"07055d0c",
			80 => x"0f05f504",
			81 => x"00000159",
			82 => x"0100ba04",
			83 => x"00420159",
			84 => x"00000159",
			85 => x"00000159",
			86 => x"0601360c",
			87 => x"0a017904",
			88 => x"0000017d",
			89 => x"0a023604",
			90 => x"0042017d",
			91 => x"0000017d",
			92 => x"06017804",
			93 => x"ff95017d",
			94 => x"0000017d",
			95 => x"0100430c",
			96 => x"01001704",
			97 => x"000001a1",
			98 => x"02074b04",
			99 => x"000001a1",
			100 => x"001501a1",
			101 => x"0208b404",
			102 => x"ffec01a1",
			103 => x"000001a1",
			104 => x"0100360c",
			105 => x"0c047a08",
			106 => x"0f05b604",
			107 => x"000001cd",
			108 => x"005701cd",
			109 => x"000001cd",
			110 => x"00032c04",
			111 => x"000001cd",
			112 => x"06010e04",
			113 => x"000001cd",
			114 => x"ff3c01cd",
			115 => x"07055d10",
			116 => x"0a02570c",
			117 => x"0d04d904",
			118 => x"000001f1",
			119 => x"0801e404",
			120 => x"000001f1",
			121 => x"007a01f1",
			122 => x"000001f1",
			123 => x"ff9b01f1",
			124 => x"06010604",
			125 => x"00000215",
			126 => x"0c045404",
			127 => x"00000215",
			128 => x"0c056208",
			129 => x"06013604",
			130 => x"00000215",
			131 => x"ffbe0215",
			132 => x"00000215",
			133 => x"0b05d710",
			134 => x"0f05e604",
			135 => x"00000239",
			136 => x"0c052a08",
			137 => x"07055d04",
			138 => x"00440239",
			139 => x"00000239",
			140 => x"00000239",
			141 => x"00000239",
			142 => x"07055d10",
			143 => x"0f05b604",
			144 => x"0000025d",
			145 => x"0a017904",
			146 => x"0000025d",
			147 => x"0c052a04",
			148 => x"0041025d",
			149 => x"0000025d",
			150 => x"0000025d",
			151 => x"0f05b604",
			152 => x"00000281",
			153 => x"0c059e0c",
			154 => x"0f0a1908",
			155 => x"0705e604",
			156 => x"00210281",
			157 => x"00000281",
			158 => x"00000281",
			159 => x"00000281",
			160 => x"07054710",
			161 => x"0601360c",
			162 => x"0600e204",
			163 => x"000002ad",
			164 => x"0b043e04",
			165 => x"000002ad",
			166 => x"003a02ad",
			167 => x"000002ad",
			168 => x"0b063c04",
			169 => x"ffd702ad",
			170 => x"000002ad",
			171 => x"02088b0c",
			172 => x"01003604",
			173 => x"000002e1",
			174 => x"0c044304",
			175 => x"000002e1",
			176 => x"ffd102e1",
			177 => x"07055d0c",
			178 => x"0100ba08",
			179 => x"0c051104",
			180 => x"009d02e1",
			181 => x"000002e1",
			182 => x"000002e1",
			183 => x"000002e1",
			184 => x"01004b10",
			185 => x"09002b04",
			186 => x"00000315",
			187 => x"0504d404",
			188 => x"00000315",
			189 => x"0704aa04",
			190 => x"00370315",
			191 => x"00000315",
			192 => x"06015308",
			193 => x"01005304",
			194 => x"00000315",
			195 => x"ffa50315",
			196 => x"00000315",
			197 => x"07055d18",
			198 => x"0f06d60c",
			199 => x"06010604",
			200 => x"00000351",
			201 => x"01002304",
			202 => x"00000351",
			203 => x"ffcc0351",
			204 => x"0100ba08",
			205 => x"0a025704",
			206 => x"008f0351",
			207 => x"00000351",
			208 => x"00000351",
			209 => x"06017804",
			210 => x"ffd80351",
			211 => x"00000351",
			212 => x"07055d14",
			213 => x"0f05b604",
			214 => x"0000037d",
			215 => x"0a017904",
			216 => x"0000037d",
			217 => x"0c052a08",
			218 => x"0b043e04",
			219 => x"0000037d",
			220 => x"003c037d",
			221 => x"0000037d",
			222 => x"0000037d",
			223 => x"0c046304",
			224 => x"000003a9",
			225 => x"0600fd04",
			226 => x"000003a9",
			227 => x"0601780c",
			228 => x"07046204",
			229 => x"000003a9",
			230 => x"06010e04",
			231 => x"000003a9",
			232 => x"ffda03a9",
			233 => x"000003a9",
			234 => x"0c046314",
			235 => x"02076704",
			236 => x"000003e5",
			237 => x"01004b0c",
			238 => x"09002704",
			239 => x"000003e5",
			240 => x"0b043d04",
			241 => x"000003e5",
			242 => x"005d03e5",
			243 => x"000003e5",
			244 => x"06015308",
			245 => x"06012704",
			246 => x"000003e5",
			247 => x"ff7103e5",
			248 => x"000003e5",
			249 => x"0c046314",
			250 => x"01004b10",
			251 => x"0d04b104",
			252 => x"00000421",
			253 => x"09002604",
			254 => x"00000421",
			255 => x"07049704",
			256 => x"002f0421",
			257 => x"00000421",
			258 => x"00000421",
			259 => x"0705ce08",
			260 => x"01005304",
			261 => x"00000421",
			262 => x"ffc10421",
			263 => x"00000421",
			264 => x"01004310",
			265 => x"0c04d00c",
			266 => x"09002604",
			267 => x"00000465",
			268 => x"01001704",
			269 => x"00000465",
			270 => x"00170465",
			271 => x"00000465",
			272 => x"0c052810",
			273 => x"0601530c",
			274 => x"0c046304",
			275 => x"00000465",
			276 => x"0600e404",
			277 => x"00000465",
			278 => x"ffbc0465",
			279 => x"00000465",
			280 => x"00000465",
			281 => x"09006c0c",
			282 => x"03039404",
			283 => x"000004b1",
			284 => x"0704bb04",
			285 => x"008b04b1",
			286 => x"000004b1",
			287 => x"0e081610",
			288 => x"0a01ec04",
			289 => x"000004b1",
			290 => x"0c044304",
			291 => x"000004b1",
			292 => x"06010e04",
			293 => x"000004b1",
			294 => x"ff1c04b1",
			295 => x"0e082c04",
			296 => x"001804b1",
			297 => x"020a2004",
			298 => x"ffe104b1",
			299 => x"000004b1",
			300 => x"0c046314",
			301 => x"02074b04",
			302 => x"000004fd",
			303 => x"0b04a10c",
			304 => x"0b043e04",
			305 => x"000004fd",
			306 => x"07049704",
			307 => x"005404fd",
			308 => x"000004fd",
			309 => x"000004fd",
			310 => x"0208b408",
			311 => x"07046104",
			312 => x"000004fd",
			313 => x"ffcb04fd",
			314 => x"07055d08",
			315 => x"07053104",
			316 => x"000004fd",
			317 => x"002804fd",
			318 => x"000004fd",
			319 => x"0802d518",
			320 => x"0e040604",
			321 => x"00000549",
			322 => x"0e082c0c",
			323 => x"0a023608",
			324 => x"0002a704",
			325 => x"00000549",
			326 => x"00760549",
			327 => x"00000549",
			328 => x"0802a504",
			329 => x"fff60549",
			330 => x"00000549",
			331 => x"0e09870c",
			332 => x"0e03bd04",
			333 => x"00000549",
			334 => x"0a024c04",
			335 => x"00000549",
			336 => x"ff970549",
			337 => x"00000549",
			338 => x"01004b18",
			339 => x"02086210",
			340 => x"06010708",
			341 => x"03043504",
			342 => x"000005a5",
			343 => x"006505a5",
			344 => x"0e046b04",
			345 => x"ff9705a5",
			346 => x"000005a5",
			347 => x"0c049504",
			348 => x"00de05a5",
			349 => x"000005a5",
			350 => x"0d06fc08",
			351 => x"0a01d404",
			352 => x"000005a5",
			353 => x"fede05a5",
			354 => x"09016d0c",
			355 => x"0c059e08",
			356 => x"0d078804",
			357 => x"006305a5",
			358 => x"000005a5",
			359 => x"000005a5",
			360 => x"ffc805a5",
			361 => x"01003614",
			362 => x"0c047910",
			363 => x"09002704",
			364 => x"000005f1",
			365 => x"0b043d04",
			366 => x"000005f1",
			367 => x"01001704",
			368 => x"000005f1",
			369 => x"004505f1",
			370 => x"000005f1",
			371 => x"0209be10",
			372 => x"0c05280c",
			373 => x"08027904",
			374 => x"000005f1",
			375 => x"0c044304",
			376 => x"000005f1",
			377 => x"ff8905f1",
			378 => x"000005f1",
			379 => x"000005f1",
			380 => x"06013620",
			381 => x"0f070514",
			382 => x"0601060c",
			383 => x"01004508",
			384 => x"01001b04",
			385 => x"0000064d",
			386 => x"0037064d",
			387 => x"0000064d",
			388 => x"01002a04",
			389 => x"0000064d",
			390 => x"ff96064d",
			391 => x"0b05bf08",
			392 => x"0a023604",
			393 => x"009f064d",
			394 => x"0000064d",
			395 => x"0000064d",
			396 => x"0a03c10c",
			397 => x"0f09a308",
			398 => x"04095904",
			399 => x"0000064d",
			400 => x"ff2b064d",
			401 => x"0000064d",
			402 => x"0000064d",
			403 => x"0c059e18",
			404 => x"0f05e604",
			405 => x"00000681",
			406 => x"0a025710",
			407 => x"0308c70c",
			408 => x"0a017904",
			409 => x"00000681",
			410 => x"0d079604",
			411 => x"004b0681",
			412 => x"00000681",
			413 => x"00000681",
			414 => x"00000681",
			415 => x"00000681",
			416 => x"06011914",
			417 => x"09007b08",
			418 => x"02071704",
			419 => x"d39e06e5",
			420 => x"f8f806e5",
			421 => x"01005308",
			422 => x"0e045304",
			423 => x"c85806e5",
			424 => x"df7606e5",
			425 => x"c7f906e5",
			426 => x"06011f08",
			427 => x"02088b04",
			428 => x"c80706e5",
			429 => x"f57706e5",
			430 => x"0c045408",
			431 => x"0208ad04",
			432 => x"c7f906e5",
			433 => x"f34106e5",
			434 => x"0704680c",
			435 => x"0d04e604",
			436 => x"c7fd06e5",
			437 => x"0b047004",
			438 => x"d3e706e5",
			439 => x"c83b06e5",
			440 => x"c7fb06e5",
			441 => x"0208b414",
			442 => x"06012710",
			443 => x"02066104",
			444 => x"00000739",
			445 => x"06010e08",
			446 => x"01005504",
			447 => x"005c0739",
			448 => x"00000739",
			449 => x"00000739",
			450 => x"ff640739",
			451 => x"0100e014",
			452 => x"0c059e10",
			453 => x"09002b04",
			454 => x"00000739",
			455 => x"0416b608",
			456 => x"020a5b04",
			457 => x"00be0739",
			458 => x"00000739",
			459 => x"00000739",
			460 => x"00000739",
			461 => x"00000739",
			462 => x"01004510",
			463 => x"0f05e608",
			464 => x"07045104",
			465 => x"00000795",
			466 => x"ffdd0795",
			467 => x"0704bc04",
			468 => x"00fd0795",
			469 => x"00000795",
			470 => x"07051f08",
			471 => x"01004b04",
			472 => x"00000795",
			473 => x"fead0795",
			474 => x"0705d114",
			475 => x"0802f410",
			476 => x"0100e80c",
			477 => x"0f074904",
			478 => x"00000795",
			479 => x"08024104",
			480 => x"00000795",
			481 => x"00b30795",
			482 => x"00000795",
			483 => x"00000795",
			484 => x"ff7a0795",
			485 => x"0802d520",
			486 => x"0308c71c",
			487 => x"0208b414",
			488 => x"0100530c",
			489 => x"0e040604",
			490 => x"00000801",
			491 => x"0802be04",
			492 => x"009a0801",
			493 => x"00000801",
			494 => x"08024e04",
			495 => x"00000801",
			496 => x"ff9e0801",
			497 => x"01010b04",
			498 => x"00ec0801",
			499 => x"00000801",
			500 => x"ffe40801",
			501 => x"0900620c",
			502 => x"0c046308",
			503 => x"0d04b104",
			504 => x"00000801",
			505 => x"00240801",
			506 => x"00000801",
			507 => x"02092008",
			508 => x"0504e204",
			509 => x"00000801",
			510 => x"fede0801",
			511 => x"00000801",
			512 => x"01003c14",
			513 => x"0f061208",
			514 => x"0c045404",
			515 => x"0000086d",
			516 => x"ffed086d",
			517 => x"0d05a808",
			518 => x"09006204",
			519 => x"014a086d",
			520 => x"0000086d",
			521 => x"0000086d",
			522 => x"0003a21c",
			523 => x"0100e018",
			524 => x"0f089c0c",
			525 => x"01005308",
			526 => x"0e04b404",
			527 => x"0000086d",
			528 => x"00ce086d",
			529 => x"ff10086d",
			530 => x"09016d08",
			531 => x"05076404",
			532 => x"012c086d",
			533 => x"0000086d",
			534 => x"0000086d",
			535 => x"ff49086d",
			536 => x"06010e04",
			537 => x"0000086d",
			538 => x"fe99086d",
			539 => x"01004718",
			540 => x"0f05e604",
			541 => x"000008d9",
			542 => x"0d05a810",
			543 => x"0d04cb04",
			544 => x"000008d9",
			545 => x"0c049908",
			546 => x"0c041e04",
			547 => x"000008d9",
			548 => x"00b708d9",
			549 => x"000008d9",
			550 => x"000008d9",
			551 => x"09014b0c",
			552 => x"07048004",
			553 => x"000008d9",
			554 => x"0600e404",
			555 => x"000008d9",
			556 => x"fefb08d9",
			557 => x"0100e010",
			558 => x"0705e60c",
			559 => x"0c04ef04",
			560 => x"000008d9",
			561 => x"05075604",
			562 => x"005308d9",
			563 => x"000008d9",
			564 => x"000008d9",
			565 => x"000008d9",
			566 => x"01004318",
			567 => x"0f06120c",
			568 => x"0c045404",
			569 => x"00000955",
			570 => x"0e02bd04",
			571 => x"00000955",
			572 => x"ffac0955",
			573 => x"0d05a808",
			574 => x"01003604",
			575 => x"01520955",
			576 => x"000a0955",
			577 => x"00000955",
			578 => x"0003a21c",
			579 => x"0100e018",
			580 => x"0f089c0c",
			581 => x"01005308",
			582 => x"03053f04",
			583 => x"00000955",
			584 => x"006b0955",
			585 => x"ff1b0955",
			586 => x"09016d08",
			587 => x"05076404",
			588 => x"01190955",
			589 => x"00000955",
			590 => x"00000955",
			591 => x"ff540955",
			592 => x"09007104",
			593 => x"00000955",
			594 => x"0b046f04",
			595 => x"00000955",
			596 => x"fe9d0955",
			597 => x"0a025720",
			598 => x"09016d1c",
			599 => x"0f06d908",
			600 => x"01004304",
			601 => x"009f09c1",
			602 => x"ff5d09c1",
			603 => x"0c059e10",
			604 => x"08023004",
			605 => x"000009c1",
			606 => x"05074808",
			607 => x"0802dd04",
			608 => x"00fd09c1",
			609 => x"000009c1",
			610 => x"000009c1",
			611 => x"000009c1",
			612 => x"ff7209c1",
			613 => x"06012710",
			614 => x"040c9a04",
			615 => x"ffed09c1",
			616 => x"07049208",
			617 => x"03037b04",
			618 => x"000009c1",
			619 => x"00c409c1",
			620 => x"000009c1",
			621 => x"0c043e04",
			622 => x"000009c1",
			623 => x"fe9709c1",
			624 => x"06012724",
			625 => x"0208151c",
			626 => x"0a022b14",
			627 => x"0f05e604",
			628 => x"ff7e0a45",
			629 => x"0705450c",
			630 => x"00022e04",
			631 => x"00000a45",
			632 => x"0a021d04",
			633 => x"01530a45",
			634 => x"00000a45",
			635 => x"00000a45",
			636 => x"06010e04",
			637 => x"00000a45",
			638 => x"feb80a45",
			639 => x"0704a904",
			640 => x"01650a45",
			641 => x"ffeb0a45",
			642 => x"0003a214",
			643 => x"0506f108",
			644 => x"0f089c04",
			645 => x"ff360a45",
			646 => x"00f60a45",
			647 => x"0802f304",
			648 => x"fea60a45",
			649 => x"030a8a04",
			650 => x"00670a45",
			651 => x"00000a45",
			652 => x"0c043f04",
			653 => x"00000a45",
			654 => x"07046804",
			655 => x"00000a45",
			656 => x"fe750a45",
			657 => x"0c046310",
			658 => x"02086208",
			659 => x"06011504",
			660 => x"011e0ab9",
			661 => x"ff140ab9",
			662 => x"01004b04",
			663 => x"01b30ab9",
			664 => x"00000ab9",
			665 => x"0802f620",
			666 => x"0c05801c",
			667 => x"0a025314",
			668 => x"09008208",
			669 => x"0e041e04",
			670 => x"00000ab9",
			671 => x"00f30ab9",
			672 => x"00032c08",
			673 => x"02084d04",
			674 => x"00000ab9",
			675 => x"00c70ab9",
			676 => x"feb20ab9",
			677 => x"0e085e04",
			678 => x"00000ab9",
			679 => x"01670ab9",
			680 => x"fee40ab9",
			681 => x"06011204",
			682 => x"00000ab9",
			683 => x"07046104",
			684 => x"00000ab9",
			685 => x"fe7a0ab9",
			686 => x"06011f28",
			687 => x"01004714",
			688 => x"0f05b604",
			689 => x"fefd0b4d",
			690 => x"06011504",
			691 => x"01bb0b4d",
			692 => x"0c045704",
			693 => x"01950b4d",
			694 => x"06011c04",
			695 => x"ff6d0b4d",
			696 => x"01150b4d",
			697 => x"0f06e30c",
			698 => x"0600e408",
			699 => x"0f05e604",
			700 => x"ff420b4d",
			701 => x"01c30b4d",
			702 => x"fe680b4d",
			703 => x"01005a04",
			704 => x"02290b4d",
			705 => x"fef00b4d",
			706 => x"0c046310",
			707 => x"0208e40c",
			708 => x"02089304",
			709 => x"fe700b4d",
			710 => x"0f070504",
			711 => x"01520b4d",
			712 => x"fee40b4d",
			713 => x"028d0b4d",
			714 => x"0003a210",
			715 => x"0c05800c",
			716 => x"02090504",
			717 => x"fe960b4d",
			718 => x"0802cc04",
			719 => x"00f40b4d",
			720 => x"04400b4d",
			721 => x"fe690b4d",
			722 => x"fe650b4d",
			723 => x"06011510",
			724 => x"0f05d208",
			725 => x"00037804",
			726 => x"ff040bd1",
			727 => x"00000bd1",
			728 => x"09008a04",
			729 => x"01910bd1",
			730 => x"ff460bd1",
			731 => x"0003a218",
			732 => x"0705d114",
			733 => x"07053104",
			734 => x"ff080bd1",
			735 => x"07055d04",
			736 => x"025b0bd1",
			737 => x"0705ce04",
			738 => x"fe9a0bd1",
			739 => x"0100e804",
			740 => x"01db0bd1",
			741 => x"00000bd1",
			742 => x"fe850bd1",
			743 => x"0b04710c",
			744 => x"02088b04",
			745 => x"feb40bd1",
			746 => x"040e6304",
			747 => x"00000bd1",
			748 => x"01580bd1",
			749 => x"0802dd04",
			750 => x"00000bd1",
			751 => x"0504d504",
			752 => x"00000bd1",
			753 => x"0e02e204",
			754 => x"00000bd1",
			755 => x"fe690bd1",
			756 => x"06011514",
			757 => x"0f05d208",
			758 => x"0c045a04",
			759 => x"00000c5d",
			760 => x"ff070c5d",
			761 => x"09008a08",
			762 => x"01004e04",
			763 => x"01990c5d",
			764 => x"006f0c5d",
			765 => x"ff570c5d",
			766 => x"0003a218",
			767 => x"0c058514",
			768 => x"0c04ef04",
			769 => x"fee80c5d",
			770 => x"07055d04",
			771 => x"021f0c5d",
			772 => x"0705ce04",
			773 => x"feb60c5d",
			774 => x"0100f304",
			775 => x"01c00c5d",
			776 => x"00000c5d",
			777 => x"fe890c5d",
			778 => x"07046c10",
			779 => x"0208c20c",
			780 => x"06011f04",
			781 => x"00000c5d",
			782 => x"08049b04",
			783 => x"fed60c5d",
			784 => x"00000c5d",
			785 => x"010a0c5d",
			786 => x"0802dd04",
			787 => x"00000c5d",
			788 => x"0c043e04",
			789 => x"00000c5d",
			790 => x"fe6d0c5d",
			791 => x"06011f1c",
			792 => x"09008218",
			793 => x"00031a08",
			794 => x"0d052804",
			795 => x"03500cd9",
			796 => x"04f40cd9",
			797 => x"02076704",
			798 => x"fe3a0cd9",
			799 => x"0c047e08",
			800 => x"03037b04",
			801 => x"ff360cd9",
			802 => x"027c0cd9",
			803 => x"ff950cd9",
			804 => x"fe660cd9",
			805 => x"0c045408",
			806 => x"0208ad04",
			807 => x"fe660cd9",
			808 => x"02770cd9",
			809 => x"04085204",
			810 => x"03150cd9",
			811 => x"07045108",
			812 => x"0c045c04",
			813 => x"fe950cd9",
			814 => x"03a30cd9",
			815 => x"040ae80c",
			816 => x"0d07ca08",
			817 => x"0d06d404",
			818 => x"fe620cd9",
			819 => x"00f20cd9",
			820 => x"fe610cd9",
			821 => x"fe610cd9",
			822 => x"01003610",
			823 => x"0f05ee04",
			824 => x"00000d5d",
			825 => x"0704bc08",
			826 => x"0d04d804",
			827 => x"00000d5d",
			828 => x"01000d5d",
			829 => x"00000d5d",
			830 => x"0003c428",
			831 => x"040a951c",
			832 => x"04097210",
			833 => x"0f061204",
			834 => x"00000d5d",
			835 => x"07054708",
			836 => x"0801e404",
			837 => x"00000d5d",
			838 => x"00c50d5d",
			839 => x"00000d5d",
			840 => x"0b063c08",
			841 => x"01004e04",
			842 => x"00000d5d",
			843 => x"fef00d5d",
			844 => x"00000d5d",
			845 => x"0c056408",
			846 => x"0003ab04",
			847 => x"00d30d5d",
			848 => x"00000d5d",
			849 => x"00000d5d",
			850 => x"0a025604",
			851 => x"00000d5d",
			852 => x"0c043d04",
			853 => x"00000d5d",
			854 => x"fec00d5d",
			855 => x"06011f2c",
			856 => x"0100451c",
			857 => x"0601150c",
			858 => x"04138708",
			859 => x"0f05e604",
			860 => x"00bb0e11",
			861 => x"01aa0e11",
			862 => x"00270e11",
			863 => x"07046c08",
			864 => x"02088b04",
			865 => x"00000e11",
			866 => x"01ad0e11",
			867 => x"03043e04",
			868 => x"00570e11",
			869 => x"feb20e11",
			870 => x"0f070f08",
			871 => x"0f06e304",
			872 => x"fe6d0e11",
			873 => x"00000e11",
			874 => x"01005a04",
			875 => x"01ee0e11",
			876 => x"ffcc0e11",
			877 => x"0c045e10",
			878 => x"0a036e0c",
			879 => x"02089304",
			880 => x"fe7b0e11",
			881 => x"01003604",
			882 => x"01920e11",
			883 => x"fec20e11",
			884 => x"083c0e11",
			885 => x"0409c710",
			886 => x"08028704",
			887 => x"fe790e11",
			888 => x"0e07dc04",
			889 => x"ff320e11",
			890 => x"01011104",
			891 => x"02d60e11",
			892 => x"ffa30e11",
			893 => x"0003a20c",
			894 => x"09018308",
			895 => x"0f097d04",
			896 => x"feb40e11",
			897 => x"02580e11",
			898 => x"fe750e11",
			899 => x"fe670e11",
			900 => x"06011510",
			901 => x"0f05d208",
			902 => x"0b046d04",
			903 => x"00000e9d",
			904 => x"fef70e9d",
			905 => x"09008a04",
			906 => x"01980e9d",
			907 => x"ff360e9d",
			908 => x"0003a218",
			909 => x"0c058514",
			910 => x"0c04ef04",
			911 => x"fedc0e9d",
			912 => x"07055d04",
			913 => x"02ab0e9d",
			914 => x"0705ce04",
			915 => x"fea00e9d",
			916 => x"0100f304",
			917 => x"01fc0e9d",
			918 => x"00000e9d",
			919 => x"fe800e9d",
			920 => x"07046c10",
			921 => x"03037b04",
			922 => x"ff110e9d",
			923 => x"040e2308",
			924 => x"08033a04",
			925 => x"00000e9d",
			926 => x"ff030e9d",
			927 => x"014c0e9d",
			928 => x"0c043e04",
			929 => x"00000e9d",
			930 => x"0802dd04",
			931 => x"00000e9d",
			932 => x"0b044d04",
			933 => x"00000e9d",
			934 => x"fe6a0e9d",
			935 => x"06011f24",
			936 => x"01004b18",
			937 => x"0f05c308",
			938 => x"02078b04",
			939 => x"fe590f39",
			940 => x"00b40f39",
			941 => x"08026404",
			942 => x"05460f39",
			943 => x"02076704",
			944 => x"00b40f39",
			945 => x"0207aa04",
			946 => x"02a10f39",
			947 => x"03bf0f39",
			948 => x"01005308",
			949 => x"0c049504",
			950 => x"fe7b0f39",
			951 => x"054d0f39",
			952 => x"fe640f39",
			953 => x"0c045408",
			954 => x"0208ad04",
			955 => x"fe5f0f39",
			956 => x"04410f39",
			957 => x"0704680c",
			958 => x"0303b004",
			959 => x"fe640f39",
			960 => x"040d8804",
			961 => x"fe830f39",
			962 => x"0b670f39",
			963 => x"040aa114",
			964 => x"08028704",
			965 => x"fe5e0f39",
			966 => x"0409c708",
			967 => x"04098704",
			968 => x"01340f39",
			969 => x"ff9e0f39",
			970 => x"040a9504",
			971 => x"fe720f39",
			972 => x"ff520f39",
			973 => x"fe5d0f39",
			974 => x"01003618",
			975 => x"09002b08",
			976 => x"04129904",
			977 => x"00000fc5",
			978 => x"fffd0fc5",
			979 => x"0704bb0c",
			980 => x"0f05b604",
			981 => x"00000fc5",
			982 => x"0d04cb04",
			983 => x"00000fc5",
			984 => x"018c0fc5",
			985 => x"00000fc5",
			986 => x"0802f628",
			987 => x"0c059e24",
			988 => x"0f074614",
			989 => x"0601060c",
			990 => x"0f062704",
			991 => x"ffd30fc5",
			992 => x"01008004",
			993 => x"00bb0fc5",
			994 => x"00000fc5",
			995 => x"0a01f704",
			996 => x"00000fc5",
			997 => x"ff180fc5",
			998 => x"0100e00c",
			999 => x"05075608",
			1000 => x"0705b804",
			1001 => x"00650fc5",
			1002 => x"015c0fc5",
			1003 => x"00000fc5",
			1004 => x"00000fc5",
			1005 => x"ff240fc5",
			1006 => x"06011504",
			1007 => x"00000fc5",
			1008 => x"fe800fc5",
			1009 => x"06012728",
			1010 => x"02082420",
			1011 => x"0a022b18",
			1012 => x"0f05e604",
			1013 => x"ff441051",
			1014 => x"01009910",
			1015 => x"0a021008",
			1016 => x"0801e404",
			1017 => x"00001051",
			1018 => x"01a71051",
			1019 => x"07049404",
			1020 => x"00a21051",
			1021 => x"ffa61051",
			1022 => x"ffa91051",
			1023 => x"06010e04",
			1024 => x"009a1051",
			1025 => x"fe8c1051",
			1026 => x"0704a904",
			1027 => x"01931051",
			1028 => x"ff391051",
			1029 => x"02090004",
			1030 => x"fe6e1051",
			1031 => x"0c059e18",
			1032 => x"0003a210",
			1033 => x"0b063c08",
			1034 => x"0f090504",
			1035 => x"00961051",
			1036 => x"ff621051",
			1037 => x"0b065b04",
			1038 => x"015f1051",
			1039 => x"00001051",
			1040 => x"0b049f04",
			1041 => x"009e1051",
			1042 => x"fea81051",
			1043 => x"fe861051",
			1044 => x"06011f1c",
			1045 => x"09008a18",
			1046 => x"0601120c",
			1047 => x"0f05d204",
			1048 => x"002b10ed",
			1049 => x"08024704",
			1050 => x"02a310ed",
			1051 => x"01b810ed",
			1052 => x"02087b04",
			1053 => x"fe5e10ed",
			1054 => x"0504f204",
			1055 => x"01ab10ed",
			1056 => x"007210ed",
			1057 => x"fe8410ed",
			1058 => x"0c046310",
			1059 => x"02089304",
			1060 => x"fe6e10ed",
			1061 => x"01003608",
			1062 => x"0c043e04",
			1063 => x"019510ed",
			1064 => x"02f010ed",
			1065 => x"fec810ed",
			1066 => x"040ae820",
			1067 => x"040ae214",
			1068 => x"05075610",
			1069 => x"0b066308",
			1070 => x"0f08d404",
			1071 => x"fe6e10ed",
			1072 => x"ffdc10ed",
			1073 => x"02097804",
			1074 => x"000010ed",
			1075 => x"043110ed",
			1076 => x"fe6b10ed",
			1077 => x"0a027004",
			1078 => x"fefb10ed",
			1079 => x"0100a104",
			1080 => x"fff510ed",
			1081 => x"043510ed",
			1082 => x"fe6510ed",
			1083 => x"06011f20",
			1084 => x"0100531c",
			1085 => x"0207aa0c",
			1086 => x"06010e08",
			1087 => x"0d050d04",
			1088 => x"001c1189",
			1089 => x"01b51189",
			1090 => x"fe761189",
			1091 => x"06011908",
			1092 => x"0413e904",
			1093 => x"01ac1189",
			1094 => x"006b1189",
			1095 => x"01003604",
			1096 => x"014a1189",
			1097 => x"ff121189",
			1098 => x"fe9f1189",
			1099 => x"04085204",
			1100 => x"03241189",
			1101 => x"0003a210",
			1102 => x"0705e60c",
			1103 => x"0f089c04",
			1104 => x"feb61189",
			1105 => x"0100e304",
			1106 => x"028b1189",
			1107 => x"fef71189",
			1108 => x"fe6e1189",
			1109 => x"07046c0c",
			1110 => x"02089304",
			1111 => x"fe8e1189",
			1112 => x"06012804",
			1113 => x"01821189",
			1114 => x"006d1189",
			1115 => x"0c04540c",
			1116 => x"0e037908",
			1117 => x"0504d404",
			1118 => x"ff911189",
			1119 => x"008e1189",
			1120 => x"ff041189",
			1121 => x"fe671189",
			1122 => x"09006210",
			1123 => x"0f05b604",
			1124 => x"ffc2120d",
			1125 => x"05059208",
			1126 => x"09005d04",
			1127 => x"0167120d",
			1128 => x"0000120d",
			1129 => x"0000120d",
			1130 => x"0802f62c",
			1131 => x"0c059e28",
			1132 => x"0f074614",
			1133 => x"0601060c",
			1134 => x"0f062704",
			1135 => x"0000120d",
			1136 => x"02066104",
			1137 => x"0000120d",
			1138 => x"003e120d",
			1139 => x"0a01f704",
			1140 => x"0000120d",
			1141 => x"ff23120d",
			1142 => x"09018710",
			1143 => x"0705ce08",
			1144 => x"07054504",
			1145 => x"00ed120d",
			1146 => x"ff3c120d",
			1147 => x"05078104",
			1148 => x"014f120d",
			1149 => x"0000120d",
			1150 => x"0000120d",
			1151 => x"ff32120d",
			1152 => x"06011504",
			1153 => x"0000120d",
			1154 => x"fe83120d",
			1155 => x"06011910",
			1156 => x"0505bf0c",
			1157 => x"0207ca08",
			1158 => x"06010704",
			1159 => x"016e12a3",
			1160 => x"fe9a12a3",
			1161 => x"01a112a3",
			1162 => x"fec312a3",
			1163 => x"04085204",
			1164 => x"019d12a3",
			1165 => x"09004f1c",
			1166 => x"0f06ac10",
			1167 => x"06012308",
			1168 => x"02088b04",
			1169 => x"000012a3",
			1170 => x"00d812a3",
			1171 => x"0f068704",
			1172 => x"fe9912a3",
			1173 => x"000012a3",
			1174 => x"06015b08",
			1175 => x"0505df04",
			1176 => x"012312a3",
			1177 => x"000012a3",
			1178 => x"045c12a3",
			1179 => x"040a3a10",
			1180 => x"00033504",
			1181 => x"fe7712a3",
			1182 => x"0e07dc04",
			1183 => x"fee512a3",
			1184 => x"0308c704",
			1185 => x"020012a3",
			1186 => x"fef512a3",
			1187 => x"06011d08",
			1188 => x"0802e504",
			1189 => x"000c12a3",
			1190 => x"ff1412a3",
			1191 => x"fe7312a3",
			1192 => x"000012a5",
			1193 => x"000012a9",
			1194 => x"000012ad",
			1195 => x"000012b1",
			1196 => x"000012b5",
			1197 => x"000012b9",
			1198 => x"000012bd",
			1199 => x"000012c1",
			1200 => x"000012c5",
			1201 => x"000012c9",
			1202 => x"000012cd",
			1203 => x"000012d1",
			1204 => x"000012d5",
			1205 => x"000012d9",
			1206 => x"000012dd",
			1207 => x"000012e1",
			1208 => x"000012e5",
			1209 => x"000012e9",
			1210 => x"000012ed",
			1211 => x"07055d04",
			1212 => x"001412f9",
			1213 => x"000012f9",
			1214 => x"07049704",
			1215 => x"00001305",
			1216 => x"ffef1305",
			1217 => x"01004308",
			1218 => x"01001704",
			1219 => x"00001319",
			1220 => x"000d1319",
			1221 => x"00001319",
			1222 => x"06012708",
			1223 => x"0600e104",
			1224 => x"0000132d",
			1225 => x"0001132d",
			1226 => x"ffe3132d",
			1227 => x"01004308",
			1228 => x"01001904",
			1229 => x"00001341",
			1230 => x"000e1341",
			1231 => x"00001341",
			1232 => x"07048004",
			1233 => x"00001355",
			1234 => x"0705ce04",
			1235 => x"fff81355",
			1236 => x"00001355",
			1237 => x"07055d08",
			1238 => x"09002704",
			1239 => x"00001369",
			1240 => x"00191369",
			1241 => x"00001369",
			1242 => x"06011504",
			1243 => x"0000137d",
			1244 => x"06017c04",
			1245 => x"ffef137d",
			1246 => x"0000137d",
			1247 => x"01004b0c",
			1248 => x"01001704",
			1249 => x"00001399",
			1250 => x"01004304",
			1251 => x"000e1399",
			1252 => x"00001399",
			1253 => x"ffff1399",
			1254 => x"0f062704",
			1255 => x"000013b5",
			1256 => x"0b05d708",
			1257 => x"0c052a04",
			1258 => x"004013b5",
			1259 => x"000013b5",
			1260 => x"000013b5",
			1261 => x"0b05d70c",
			1262 => x"0f05e604",
			1263 => x"000013d1",
			1264 => x"07055d04",
			1265 => x"003813d1",
			1266 => x"000013d1",
			1267 => x"000013d1",
			1268 => x"0601270c",
			1269 => x"0600e104",
			1270 => x"000013ed",
			1271 => x"06011204",
			1272 => x"002013ed",
			1273 => x"000013ed",
			1274 => x"ffdd13ed",
			1275 => x"06011404",
			1276 => x"00001409",
			1277 => x"06015b08",
			1278 => x"06011504",
			1279 => x"00001409",
			1280 => x"ffcb1409",
			1281 => x"00001409",
			1282 => x"0601360c",
			1283 => x"0a017904",
			1284 => x"0000142d",
			1285 => x"0a035d04",
			1286 => x"0033142d",
			1287 => x"0000142d",
			1288 => x"06017804",
			1289 => x"ff9f142d",
			1290 => x"0000142d",
			1291 => x"06011208",
			1292 => x"0600e104",
			1293 => x"00001451",
			1294 => x"00031451",
			1295 => x"0c045404",
			1296 => x"00001451",
			1297 => x"0b044f04",
			1298 => x"00001451",
			1299 => x"ffb61451",
			1300 => x"0601360c",
			1301 => x"0801e404",
			1302 => x"0000147d",
			1303 => x"0a023604",
			1304 => x"004f147d",
			1305 => x"0000147d",
			1306 => x"06017808",
			1307 => x"0409c704",
			1308 => x"0000147d",
			1309 => x"ff6c147d",
			1310 => x"0000147d",
			1311 => x"0705d110",
			1312 => x"0f06d604",
			1313 => x"000014a1",
			1314 => x"08023004",
			1315 => x"000014a1",
			1316 => x"0100e004",
			1317 => x"004a14a1",
			1318 => x"000014a1",
			1319 => x"000014a1",
			1320 => x"07054710",
			1321 => x"0d04cb04",
			1322 => x"000014c5",
			1323 => x"06013d08",
			1324 => x"0600e204",
			1325 => x"000014c5",
			1326 => x"001014c5",
			1327 => x"000014c5",
			1328 => x"ffa114c5",
			1329 => x"07055d10",
			1330 => x"0f05f504",
			1331 => x"000014e9",
			1332 => x"0100ba08",
			1333 => x"0c052a04",
			1334 => x"004d14e9",
			1335 => x"000014e9",
			1336 => x"000014e9",
			1337 => x"000014e9",
			1338 => x"07055d10",
			1339 => x"0f05b604",
			1340 => x"0000150d",
			1341 => x"0c052a08",
			1342 => x"0b043e04",
			1343 => x"0000150d",
			1344 => x"0034150d",
			1345 => x"0000150d",
			1346 => x"0000150d",
			1347 => x"01004710",
			1348 => x"0f05e604",
			1349 => x"00001539",
			1350 => x"05059208",
			1351 => x"0c049904",
			1352 => x"00651539",
			1353 => x"00001539",
			1354 => x"00001539",
			1355 => x"00032404",
			1356 => x"00001539",
			1357 => x"ff341539",
			1358 => x"07055d14",
			1359 => x"0b05970c",
			1360 => x"06011408",
			1361 => x"0600e104",
			1362 => x"00001565",
			1363 => x"001f1565",
			1364 => x"ffc71565",
			1365 => x"06012504",
			1366 => x"00001565",
			1367 => x"00771565",
			1368 => x"ff941565",
			1369 => x"06013610",
			1370 => x"0f062704",
			1371 => x"00001599",
			1372 => x"07054708",
			1373 => x"0a024904",
			1374 => x"004b1599",
			1375 => x"00001599",
			1376 => x"00001599",
			1377 => x"04095904",
			1378 => x"00001599",
			1379 => x"06017804",
			1380 => x"ff5c1599",
			1381 => x"00001599",
			1382 => x"01004b10",
			1383 => x"0505df0c",
			1384 => x"0d050d04",
			1385 => x"000015d5",
			1386 => x"0504f304",
			1387 => x"000015d5",
			1388 => x"006c15d5",
			1389 => x"000015d5",
			1390 => x"0d06fc08",
			1391 => x"0600e404",
			1392 => x"000015d5",
			1393 => x"ff9f15d5",
			1394 => x"09016d04",
			1395 => x"000715d5",
			1396 => x"000015d5",
			1397 => x"0c046310",
			1398 => x"0b049d0c",
			1399 => x"09002b04",
			1400 => x"00001611",
			1401 => x"01004b04",
			1402 => x"00371611",
			1403 => x"00001611",
			1404 => x"00001611",
			1405 => x"0601530c",
			1406 => x"06011204",
			1407 => x"00001611",
			1408 => x"07046204",
			1409 => x"00001611",
			1410 => x"ff821611",
			1411 => x"00001611",
			1412 => x"0705e614",
			1413 => x"0f05e604",
			1414 => x"0000163d",
			1415 => x"01001504",
			1416 => x"0000163d",
			1417 => x"0100e008",
			1418 => x"05075604",
			1419 => x"0025163d",
			1420 => x"0000163d",
			1421 => x"0000163d",
			1422 => x"0000163d",
			1423 => x"0208b418",
			1424 => x"0601120c",
			1425 => x"09008a08",
			1426 => x"0600e804",
			1427 => x"00001681",
			1428 => x"00161681",
			1429 => x"00001681",
			1430 => x"0a01db04",
			1431 => x"00001681",
			1432 => x"09003404",
			1433 => x"00001681",
			1434 => x"ff5e1681",
			1435 => x"07055d08",
			1436 => x"0100ba04",
			1437 => x"009d1681",
			1438 => x"00001681",
			1439 => x"00001681",
			1440 => x"0208b40c",
			1441 => x"06010a04",
			1442 => x"000016bd",
			1443 => x"0a01db04",
			1444 => x"000016bd",
			1445 => x"ff8816bd",
			1446 => x"0705e610",
			1447 => x"0100e00c",
			1448 => x"0416b608",
			1449 => x"020a5b04",
			1450 => x"009a16bd",
			1451 => x"000016bd",
			1452 => x"000016bd",
			1453 => x"000016bd",
			1454 => x"000016bd",
			1455 => x"0c046314",
			1456 => x"02074b04",
			1457 => x"00001701",
			1458 => x"01004b0c",
			1459 => x"01001704",
			1460 => x"00001701",
			1461 => x"07049704",
			1462 => x"005b1701",
			1463 => x"00001701",
			1464 => x"00001701",
			1465 => x"0209810c",
			1466 => x"0b063c08",
			1467 => x"07046104",
			1468 => x"00001701",
			1469 => x"ffcf1701",
			1470 => x"00001701",
			1471 => x"00001701",
			1472 => x"01004b10",
			1473 => x"0f061204",
			1474 => x"0000174d",
			1475 => x"0c049808",
			1476 => x"06011904",
			1477 => x"00e5174d",
			1478 => x"0000174d",
			1479 => x"0000174d",
			1480 => x"0f091f08",
			1481 => x"0a01cf04",
			1482 => x"0000174d",
			1483 => x"ff10174d",
			1484 => x"0901800c",
			1485 => x"0b065b08",
			1486 => x"09014f04",
			1487 => x"0000174d",
			1488 => x"0030174d",
			1489 => x"0000174d",
			1490 => x"0000174d",
			1491 => x"09006c0c",
			1492 => x"03039404",
			1493 => x"00001799",
			1494 => x"0704bb04",
			1495 => x"00821799",
			1496 => x"00001799",
			1497 => x"06016310",
			1498 => x"00032404",
			1499 => x"00001799",
			1500 => x"06010e04",
			1501 => x"00001799",
			1502 => x"0c044304",
			1503 => x"00001799",
			1504 => x"ff0f1799",
			1505 => x"0100e008",
			1506 => x"0100d604",
			1507 => x"00001799",
			1508 => x"00571799",
			1509 => x"00001799",
			1510 => x"0601361c",
			1511 => x"0f070514",
			1512 => x"0601060c",
			1513 => x"01004508",
			1514 => x"01001b04",
			1515 => x"000017ed",
			1516 => x"003b17ed",
			1517 => x"000017ed",
			1518 => x"01002a04",
			1519 => x"000017ed",
			1520 => x"ff8817ed",
			1521 => x"0b05bf04",
			1522 => x"00a817ed",
			1523 => x"000017ed",
			1524 => x"0209be08",
			1525 => x"0b063c04",
			1526 => x"ff1117ed",
			1527 => x"000017ed",
			1528 => x"0c051104",
			1529 => x"007117ed",
			1530 => x"000017ed",
			1531 => x"07055d20",
			1532 => x"02088b14",
			1533 => x"0a01f70c",
			1534 => x"0e04db04",
			1535 => x"00001839",
			1536 => x"0600e204",
			1537 => x"00001839",
			1538 => x"001b1839",
			1539 => x"06010604",
			1540 => x"00001839",
			1541 => x"ff711839",
			1542 => x"0100ba08",
			1543 => x"0c051104",
			1544 => x"00911839",
			1545 => x"00001839",
			1546 => x"00001839",
			1547 => x"06017804",
			1548 => x"ffdc1839",
			1549 => x"00001839",
			1550 => x"0802f618",
			1551 => x"0705e614",
			1552 => x"0f05e604",
			1553 => x"0000187d",
			1554 => x"0100e30c",
			1555 => x"0801e404",
			1556 => x"0000187d",
			1557 => x"05075604",
			1558 => x"008d187d",
			1559 => x"0000187d",
			1560 => x"0000187d",
			1561 => x"0000187d",
			1562 => x"06011504",
			1563 => x"0000187d",
			1564 => x"09004204",
			1565 => x"0000187d",
			1566 => x"ff1b187d",
			1567 => x"0b049d18",
			1568 => x"0d04b304",
			1569 => x"000018c9",
			1570 => x"0c046310",
			1571 => x"0900820c",
			1572 => x"07049708",
			1573 => x"09002704",
			1574 => x"000018c9",
			1575 => x"004518c9",
			1576 => x"000018c9",
			1577 => x"000018c9",
			1578 => x"000018c9",
			1579 => x"0d06fc08",
			1580 => x"09007104",
			1581 => x"000018c9",
			1582 => x"ffa318c9",
			1583 => x"09016d04",
			1584 => x"000a18c9",
			1585 => x"000018c9",
			1586 => x"06013620",
			1587 => x"0f074914",
			1588 => x"06010e0c",
			1589 => x"0f05d204",
			1590 => x"0000192d",
			1591 => x"0505f904",
			1592 => x"00dc192d",
			1593 => x"0000192d",
			1594 => x"09004604",
			1595 => x"0000192d",
			1596 => x"ff10192d",
			1597 => x"07054708",
			1598 => x"0a029904",
			1599 => x"00f5192d",
			1600 => x"0000192d",
			1601 => x"0000192d",
			1602 => x"020a2008",
			1603 => x"0705d004",
			1604 => x"feb4192d",
			1605 => x"0000192d",
			1606 => x"0705cf08",
			1607 => x"020a5b04",
			1608 => x"00b8192d",
			1609 => x"0000192d",
			1610 => x"0000192d",
			1611 => x"0802d518",
			1612 => x"0c059e14",
			1613 => x"0e040604",
			1614 => x"00001979",
			1615 => x"0e08a10c",
			1616 => x"0a023608",
			1617 => x"0801e404",
			1618 => x"00001979",
			1619 => x"007c1979",
			1620 => x"00001979",
			1621 => x"00001979",
			1622 => x"00001979",
			1623 => x"0c045404",
			1624 => x"00001979",
			1625 => x"0e098708",
			1626 => x"0e02ea04",
			1627 => x"00001979",
			1628 => x"ff7f1979",
			1629 => x"00001979",
			1630 => x"06013624",
			1631 => x"0f074918",
			1632 => x"0601060c",
			1633 => x"0f05b604",
			1634 => x"000019ed",
			1635 => x"0505f604",
			1636 => x"00cd19ed",
			1637 => x"000019ed",
			1638 => x"01003604",
			1639 => x"000019ed",
			1640 => x"0a01f704",
			1641 => x"000019ed",
			1642 => x"ff0619ed",
			1643 => x"07054708",
			1644 => x"0a029904",
			1645 => x"00e819ed",
			1646 => x"000019ed",
			1647 => x"000019ed",
			1648 => x"020a200c",
			1649 => x"0705d008",
			1650 => x"01002504",
			1651 => x"000019ed",
			1652 => x"feb819ed",
			1653 => x"000019ed",
			1654 => x"0705cf08",
			1655 => x"020a5b04",
			1656 => x"00a819ed",
			1657 => x"000019ed",
			1658 => x"000019ed",
			1659 => x"0208b414",
			1660 => x"06012710",
			1661 => x"02066104",
			1662 => x"00001a41",
			1663 => x"06010e08",
			1664 => x"01005504",
			1665 => x"00561a41",
			1666 => x"00001a41",
			1667 => x"00001a41",
			1668 => x"ff6c1a41",
			1669 => x"0100e014",
			1670 => x"0c059e10",
			1671 => x"09002b04",
			1672 => x"00001a41",
			1673 => x"0006f108",
			1674 => x"020a5b04",
			1675 => x"00ad1a41",
			1676 => x"00001a41",
			1677 => x"00001a41",
			1678 => x"00001a41",
			1679 => x"00001a41",
			1680 => x"01004518",
			1681 => x"02086210",
			1682 => x"06010e08",
			1683 => x"03043504",
			1684 => x"00001abd",
			1685 => x"00211abd",
			1686 => x"0e045304",
			1687 => x"ffc61abd",
			1688 => x"00001abd",
			1689 => x"0704aa04",
			1690 => x"00d31abd",
			1691 => x"00001abd",
			1692 => x"07053410",
			1693 => x"0002dd04",
			1694 => x"00001abd",
			1695 => x"02092008",
			1696 => x"0c043e04",
			1697 => x"00001abd",
			1698 => x"fefb1abd",
			1699 => x"00001abd",
			1700 => x"07055d0c",
			1701 => x"06015608",
			1702 => x"02078004",
			1703 => x"00001abd",
			1704 => x"00bf1abd",
			1705 => x"00001abd",
			1706 => x"06017808",
			1707 => x"04095904",
			1708 => x"00001abd",
			1709 => x"ff701abd",
			1710 => x"00001abd",
			1711 => x"0a027224",
			1712 => x"0705e620",
			1713 => x"0e07dc14",
			1714 => x"01004b0c",
			1715 => x"0d04d804",
			1716 => x"00001b19",
			1717 => x"06011504",
			1718 => x"00bb1b19",
			1719 => x"00001b19",
			1720 => x"04089204",
			1721 => x"00001b19",
			1722 => x"ff781b19",
			1723 => x"09016d08",
			1724 => x"00031a04",
			1725 => x"00001b19",
			1726 => x"00e31b19",
			1727 => x"00001b19",
			1728 => x"00001b19",
			1729 => x"06012704",
			1730 => x"00001b19",
			1731 => x"01002304",
			1732 => x"00001b19",
			1733 => x"ff2a1b19",
			1734 => x"01004518",
			1735 => x"02086210",
			1736 => x"06010e08",
			1737 => x"0303b004",
			1738 => x"00001b85",
			1739 => x"00b01b85",
			1740 => x"0e044b04",
			1741 => x"ff6e1b85",
			1742 => x"00001b85",
			1743 => x"0704aa04",
			1744 => x"013f1b85",
			1745 => x"00001b85",
			1746 => x"0c050d08",
			1747 => x"06011504",
			1748 => x"00001b85",
			1749 => x"fead1b85",
			1750 => x"0c058514",
			1751 => x"0e06e204",
			1752 => x"00001b85",
			1753 => x"0003a20c",
			1754 => x"0002cc04",
			1755 => x"00001b85",
			1756 => x"0705d104",
			1757 => x"01291b85",
			1758 => x"00001b85",
			1759 => x"00001b85",
			1760 => x"ff511b85",
			1761 => x"01004718",
			1762 => x"0f05e604",
			1763 => x"00001bf1",
			1764 => x"0d05a810",
			1765 => x"0d04cb04",
			1766 => x"00001bf1",
			1767 => x"0c049908",
			1768 => x"0c041e04",
			1769 => x"00001bf1",
			1770 => x"00a91bf1",
			1771 => x"00001bf1",
			1772 => x"00001bf1",
			1773 => x"0100b70c",
			1774 => x"07046c04",
			1775 => x"00001bf1",
			1776 => x"0600e404",
			1777 => x"00001bf1",
			1778 => x"ff0d1bf1",
			1779 => x"0100e010",
			1780 => x"0c059e0c",
			1781 => x"0c04ef04",
			1782 => x"00001bf1",
			1783 => x"0705e604",
			1784 => x"00351bf1",
			1785 => x"00001bf1",
			1786 => x"00001bf1",
			1787 => x"00001bf1",
			1788 => x"01004318",
			1789 => x"0f06120c",
			1790 => x"0c045404",
			1791 => x"00001c6d",
			1792 => x"07045104",
			1793 => x"00001c6d",
			1794 => x"ffaa1c6d",
			1795 => x"0d05a808",
			1796 => x"01003c04",
			1797 => x"01271c6d",
			1798 => x"00001c6d",
			1799 => x"00001c6d",
			1800 => x"0003a21c",
			1801 => x"0100e018",
			1802 => x"0f089c0c",
			1803 => x"01005308",
			1804 => x"03053f04",
			1805 => x"00001c6d",
			1806 => x"00621c6d",
			1807 => x"ff271c6d",
			1808 => x"09016d08",
			1809 => x"0d07a304",
			1810 => x"01071c6d",
			1811 => x"00001c6d",
			1812 => x"00001c6d",
			1813 => x"ff5f1c6d",
			1814 => x"09007104",
			1815 => x"00001c6d",
			1816 => x"0802e004",
			1817 => x"00001c6d",
			1818 => x"fe961c6d",
			1819 => x"0802dd24",
			1820 => x"0308c720",
			1821 => x"0208b418",
			1822 => x"0a01fa0c",
			1823 => x"0d067708",
			1824 => x"02066104",
			1825 => x"00001ce1",
			1826 => x"00b01ce1",
			1827 => x"00001ce1",
			1828 => x"01004104",
			1829 => x"00001ce1",
			1830 => x"0b049e04",
			1831 => x"00001ce1",
			1832 => x"ff771ce1",
			1833 => x"01010b04",
			1834 => x"01041ce1",
			1835 => x"00001ce1",
			1836 => x"ffce1ce1",
			1837 => x"06011508",
			1838 => x"0d052704",
			1839 => x"00611ce1",
			1840 => x"00001ce1",
			1841 => x"09004204",
			1842 => x"00001ce1",
			1843 => x"0003a204",
			1844 => x"00001ce1",
			1845 => x"0c043d04",
			1846 => x"00001ce1",
			1847 => x"fec21ce1",
			1848 => x"0c046318",
			1849 => x"01003608",
			1850 => x"0f05b604",
			1851 => x"00001d65",
			1852 => x"01451d65",
			1853 => x"0e04a008",
			1854 => x"0f073904",
			1855 => x"ff951d65",
			1856 => x"00001d65",
			1857 => x"0a027004",
			1858 => x"00ad1d65",
			1859 => x"00001d65",
			1860 => x"0003a21c",
			1861 => x"0c058518",
			1862 => x"0c050d0c",
			1863 => x"01005308",
			1864 => x"0e047104",
			1865 => x"00001d65",
			1866 => x"00261d65",
			1867 => x"ff3d1d65",
			1868 => x"08024704",
			1869 => x"00001d65",
			1870 => x"0100ff04",
			1871 => x"01321d65",
			1872 => x"00001d65",
			1873 => x"ff771d65",
			1874 => x"0802d204",
			1875 => x"00001d65",
			1876 => x"07046104",
			1877 => x"00001d65",
			1878 => x"0b044d04",
			1879 => x"00001d65",
			1880 => x"feae1d65",
			1881 => x"06012724",
			1882 => x"02081b1c",
			1883 => x"0a022b14",
			1884 => x"0f05e604",
			1885 => x"ff851df1",
			1886 => x"0705450c",
			1887 => x"00022e04",
			1888 => x"00001df1",
			1889 => x"0a021d04",
			1890 => x"01421df1",
			1891 => x"00001df1",
			1892 => x"00001df1",
			1893 => x"06010e04",
			1894 => x"00001df1",
			1895 => x"febe1df1",
			1896 => x"0704a904",
			1897 => x"015f1df1",
			1898 => x"00001df1",
			1899 => x"0003a218",
			1900 => x"00038c0c",
			1901 => x"0e082c08",
			1902 => x"0f08b104",
			1903 => x"ff531df1",
			1904 => x"00d91df1",
			1905 => x"feb91df1",
			1906 => x"0c056408",
			1907 => x"0a024704",
			1908 => x"00001df1",
			1909 => x"01091df1",
			1910 => x"ffce1df1",
			1911 => x"0c043f04",
			1912 => x"00001df1",
			1913 => x"07046804",
			1914 => x"00001df1",
			1915 => x"fe771df1",
			1916 => x"0c04631c",
			1917 => x"09005d0c",
			1918 => x"0f05b604",
			1919 => x"00001e75",
			1920 => x"0d04cb04",
			1921 => x"00001e75",
			1922 => x"01ab1e75",
			1923 => x"0e04e208",
			1924 => x"0e04a004",
			1925 => x"ff641e75",
			1926 => x"00001e75",
			1927 => x"0a027004",
			1928 => x"00f21e75",
			1929 => x"00001e75",
			1930 => x"0802f620",
			1931 => x"0c05801c",
			1932 => x"0a025314",
			1933 => x"09008208",
			1934 => x"0e041e04",
			1935 => x"00001e75",
			1936 => x"00e31e75",
			1937 => x"00032c08",
			1938 => x"0f087204",
			1939 => x"00001e75",
			1940 => x"00bd1e75",
			1941 => x"febc1e75",
			1942 => x"0e085e04",
			1943 => x"00001e75",
			1944 => x"01561e75",
			1945 => x"fef01e75",
			1946 => x"07046104",
			1947 => x"00001e75",
			1948 => x"fe871e75",
			1949 => x"06011f20",
			1950 => x"01004b14",
			1951 => x"0f05b604",
			1952 => x"fec21f01",
			1953 => x"08026404",
			1954 => x"03a31f01",
			1955 => x"0c048f08",
			1956 => x"03058004",
			1957 => x"02411f01",
			1958 => x"02dd1f01",
			1959 => x"ffb71f01",
			1960 => x"01005108",
			1961 => x"0d054004",
			1962 => x"feaa1f01",
			1963 => x"01a81f01",
			1964 => x"fe6b1f01",
			1965 => x"0c04540c",
			1966 => x"0f05ee04",
			1967 => x"fe691f01",
			1968 => x"01003204",
			1969 => x"02781f01",
			1970 => x"fe621f01",
			1971 => x"04085204",
			1972 => x"02981f01",
			1973 => x"07045108",
			1974 => x"0c045c04",
			1975 => x"fe9f1f01",
			1976 => x"02c71f01",
			1977 => x"040ae80c",
			1978 => x"05075608",
			1979 => x"0e089604",
			1980 => x"febb1f01",
			1981 => x"05d01f01",
			1982 => x"fe621f01",
			1983 => x"fe621f01",
			1984 => x"06011510",
			1985 => x"09008a0c",
			1986 => x"0f05d204",
			1987 => x"00001f95",
			1988 => x"04138704",
			1989 => x"01a11f95",
			1990 => x"00041f95",
			1991 => x"fee11f95",
			1992 => x"0c046318",
			1993 => x"02088b08",
			1994 => x"02087b04",
			1995 => x"fe7b1f95",
			1996 => x"00001f95",
			1997 => x"01004508",
			1998 => x"06013d04",
			1999 => x"01921f95",
			2000 => x"03f61f95",
			2001 => x"040c3e04",
			2002 => x"00011f95",
			2003 => x"fef71f95",
			2004 => x"0409c710",
			2005 => x"08028704",
			2006 => x"fe851f95",
			2007 => x"0f089c04",
			2008 => x"ff391f95",
			2009 => x"0c059f04",
			2010 => x"025c1f95",
			2011 => x"ffab1f95",
			2012 => x"0003a20c",
			2013 => x"0705cf08",
			2014 => x"02099d04",
			2015 => x"febd1f95",
			2016 => x"027b1f95",
			2017 => x"fe7b1f95",
			2018 => x"07046204",
			2019 => x"00001f95",
			2020 => x"fe661f95",
			2021 => x"06011914",
			2022 => x"01004708",
			2023 => x"02076704",
			2024 => x"005d2011",
			2025 => x"01962011",
			2026 => x"0f067a04",
			2027 => x"febf2011",
			2028 => x"09008904",
			2029 => x"00bf2011",
			2030 => x"ff3f2011",
			2031 => x"04085204",
			2032 => x"022c2011",
			2033 => x"0c046314",
			2034 => x"0208bb08",
			2035 => x"08048f04",
			2036 => x"fe872011",
			2037 => x"00002011",
			2038 => x"0b049d08",
			2039 => x"00067e04",
			2040 => x"01562011",
			2041 => x"03962011",
			2042 => x"ff932011",
			2043 => x"040a3a10",
			2044 => x"00033504",
			2045 => x"fe732011",
			2046 => x"0c050d04",
			2047 => x"fec62011",
			2048 => x"0705e704",
			2049 => x"02392011",
			2050 => x"ff0f2011",
			2051 => x"fe712011",
			2052 => x"0601151c",
			2053 => x"0207aa14",
			2054 => x"01004308",
			2055 => x"05051004",
			2056 => x"000020b5",
			2057 => x"010520b5",
			2058 => x"0e04f004",
			2059 => x"fef520b5",
			2060 => x"0b053104",
			2061 => x"005a20b5",
			2062 => x"000020b5",
			2063 => x"01005504",
			2064 => x"018120b5",
			2065 => x"000020b5",
			2066 => x"02098124",
			2067 => x"0f089c14",
			2068 => x"01002d0c",
			2069 => x"02087b04",
			2070 => x"ff3320b5",
			2071 => x"0505f604",
			2072 => x"00f520b5",
			2073 => x"000020b5",
			2074 => x"0504d404",
			2075 => x"000020b5",
			2076 => x"fe7720b5",
			2077 => x"07054708",
			2078 => x"0003c404",
			2079 => x"017320b5",
			2080 => x"000020b5",
			2081 => x"0802a504",
			2082 => x"feca20b5",
			2083 => x"000020b5",
			2084 => x"0c058010",
			2085 => x"0601940c",
			2086 => x"0100e008",
			2087 => x"020a5b04",
			2088 => x"020d20b5",
			2089 => x"000020b5",
			2090 => x"000020b5",
			2091 => x"000020b5",
			2092 => x"feab20b5",
			2093 => x"06012734",
			2094 => x"01004718",
			2095 => x"0601150c",
			2096 => x"01001804",
			2097 => x"00002169",
			2098 => x"0d04bf04",
			2099 => x"00002169",
			2100 => x"01972169",
			2101 => x"02087b04",
			2102 => x"feb42169",
			2103 => x"07046804",
			2104 => x"01732169",
			2105 => x"00002169",
			2106 => x"06012514",
			2107 => x"07048008",
			2108 => x"0207da04",
			2109 => x"00002169",
			2110 => x"00c32169",
			2111 => x"0600fb08",
			2112 => x"0d05e904",
			2113 => x"00b22169",
			2114 => x"ff8d2169",
			2115 => x"fe8e2169",
			2116 => x"04089204",
			2117 => x"03962169",
			2118 => x"00002169",
			2119 => x"040a3a10",
			2120 => x"00033504",
			2121 => x"fe762169",
			2122 => x"09016d08",
			2123 => x"0307f404",
			2124 => x"ff0b2169",
			2125 => x"01d62169",
			2126 => x"feff2169",
			2127 => x"0e032608",
			2128 => x"02096004",
			2129 => x"feb82169",
			2130 => x"03282169",
			2131 => x"0704680c",
			2132 => x"07046608",
			2133 => x"0504e404",
			2134 => x"00002169",
			2135 => x"ff652169",
			2136 => x"00002169",
			2137 => x"fe762169",
			2138 => x"06011f1c",
			2139 => x"01004b18",
			2140 => x"0a01cf04",
			2141 => x"045521ed",
			2142 => x"0c048f10",
			2143 => x"03037b04",
			2144 => x"ff2d21ed",
			2145 => x"02076704",
			2146 => x"00d321ed",
			2147 => x"03058704",
			2148 => x"022021ed",
			2149 => x"02d821ed",
			2150 => x"fe7c21ed",
			2151 => x"fe6921ed",
			2152 => x"07046c0c",
			2153 => x"02089304",
			2154 => x"fe6721ed",
			2155 => x"0208f004",
			2156 => x"01c221ed",
			2157 => x"030821ed",
			2158 => x"0c043a08",
			2159 => x"08046904",
			2160 => x"ff7721ed",
			2161 => x"00a121ed",
			2162 => x"040ae810",
			2163 => x"040ae204",
			2164 => x"fe8021ed",
			2165 => x"0802f304",
			2166 => x"fea721ed",
			2167 => x"0003c804",
			2168 => x"07e621ed",
			2169 => x"fef121ed",
			2170 => x"fe6421ed",
			2171 => x"01003c14",
			2172 => x"0c049910",
			2173 => x"0f05b604",
			2174 => x"ff672261",
			2175 => x"01003604",
			2176 => x"01ba2261",
			2177 => x"0a027704",
			2178 => x"00d12261",
			2179 => x"00002261",
			2180 => x"ff152261",
			2181 => x"0802f424",
			2182 => x"0c059e20",
			2183 => x"0f074610",
			2184 => x"09007508",
			2185 => x"0d050d04",
			2186 => x"ffbb2261",
			2187 => x"00a72261",
			2188 => x"0a018404",
			2189 => x"00002261",
			2190 => x"fecc2261",
			2191 => x"0100e00c",
			2192 => x"02092408",
			2193 => x"04097204",
			2194 => x"018f2261",
			2195 => x"00002261",
			2196 => x"01ba2261",
			2197 => x"00002261",
			2198 => x"feb12261",
			2199 => x"fe7b2261",
			2200 => x"06011f1c",
			2201 => x"01005318",
			2202 => x"06011510",
			2203 => x"08024704",
			2204 => x"034122fd",
			2205 => x"09007104",
			2206 => x"01d322fd",
			2207 => x"0b049104",
			2208 => x"01f722fd",
			2209 => x"fff122fd",
			2210 => x"02088b04",
			2211 => x"fe3922fd",
			2212 => x"01a822fd",
			2213 => x"fe7922fd",
			2214 => x"07046c0c",
			2215 => x"02089304",
			2216 => x"fe7022fd",
			2217 => x"0d04f304",
			2218 => x"024222fd",
			2219 => x"010c22fd",
			2220 => x"0a023310",
			2221 => x"0507390c",
			2222 => x"0c04ef04",
			2223 => x"fec522fd",
			2224 => x"09016d04",
			2225 => x"068e22fd",
			2226 => x"ff6b22fd",
			2227 => x"fe6a22fd",
			2228 => x"0c045e14",
			2229 => x"0c045c0c",
			2230 => x"0c045408",
			2231 => x"09003d04",
			2232 => x"000022fd",
			2233 => x"fe8122fd",
			2234 => x"fe7222fd",
			2235 => x"03045e04",
			2236 => x"079122fd",
			2237 => x"ffad22fd",
			2238 => x"fe6722fd",
			2239 => x"06011f1c",
			2240 => x"09008a18",
			2241 => x"06011510",
			2242 => x"0f05c304",
			2243 => x"ffd72391",
			2244 => x"08024704",
			2245 => x"03182391",
			2246 => x"09007704",
			2247 => x"01cb2391",
			2248 => x"00fa2391",
			2249 => x"02088b04",
			2250 => x"fe462391",
			2251 => x"01932391",
			2252 => x"fe7c2391",
			2253 => x"07046c0c",
			2254 => x"02089304",
			2255 => x"fe732391",
			2256 => x"0f06ed04",
			2257 => x"02232391",
			2258 => x"00bd2391",
			2259 => x"04085204",
			2260 => x"020f2391",
			2261 => x"0409c70c",
			2262 => x"0c059e08",
			2263 => x"0208b404",
			2264 => x"feb82391",
			2265 => x"05452391",
			2266 => x"fe6d2391",
			2267 => x"0c045e10",
			2268 => x"0c045c08",
			2269 => x"0c045404",
			2270 => x"ff692391",
			2271 => x"fe752391",
			2272 => x"03045e04",
			2273 => x"05292391",
			2274 => x"ffbc2391",
			2275 => x"fe682391",
			2276 => x"0601151c",
			2277 => x"0207aa14",
			2278 => x"01004308",
			2279 => x"05051004",
			2280 => x"0000244d",
			2281 => x"00ed244d",
			2282 => x"0e04f004",
			2283 => x"ff0e244d",
			2284 => x"0d05ed04",
			2285 => x"003a244d",
			2286 => x"0000244d",
			2287 => x"01005504",
			2288 => x"0171244d",
			2289 => x"0000244d",
			2290 => x"02098130",
			2291 => x"0f089c1c",
			2292 => x"01002d0c",
			2293 => x"02087b04",
			2294 => x"ff5f244d",
			2295 => x"0505f604",
			2296 => x"00d3244d",
			2297 => x"0000244d",
			2298 => x"0504d404",
			2299 => x"0000244d",
			2300 => x"02092004",
			2301 => x"fe72244d",
			2302 => x"02092404",
			2303 => x"0000244d",
			2304 => x"ff97244d",
			2305 => x"06013608",
			2306 => x"0e086804",
			2307 => x"013b244d",
			2308 => x"0000244d",
			2309 => x"0f091f04",
			2310 => x"fee0244d",
			2311 => x"0f092a04",
			2312 => x"0000244d",
			2313 => x"ffdf244d",
			2314 => x"0c058010",
			2315 => x"0601940c",
			2316 => x"0100e008",
			2317 => x"020a5b04",
			2318 => x"01bb244d",
			2319 => x"0000244d",
			2320 => x"0000244d",
			2321 => x"0000244d",
			2322 => x"febe244d",
			2323 => x"06011f20",
			2324 => x"09008a1c",
			2325 => x"0207aa0c",
			2326 => x"06010e08",
			2327 => x"0304d604",
			2328 => x"004524e1",
			2329 => x"01de24e1",
			2330 => x"fe6524e1",
			2331 => x"06011908",
			2332 => x"03058704",
			2333 => x"01a524e1",
			2334 => x"026f24e1",
			2335 => x"01003604",
			2336 => x"016824e1",
			2337 => x"ff0924e1",
			2338 => x"fe9024e1",
			2339 => x"04085204",
			2340 => x"063724e1",
			2341 => x"07046c08",
			2342 => x"02089304",
			2343 => x"fe8224e1",
			2344 => x"016624e1",
			2345 => x"0003a210",
			2346 => x"0c059e0c",
			2347 => x"0f089c04",
			2348 => x"feae24e1",
			2349 => x"0100e304",
			2350 => x"038024e1",
			2351 => x"fed624e1",
			2352 => x"fe6b24e1",
			2353 => x"0c04540c",
			2354 => x"0b048108",
			2355 => x"0b046d04",
			2356 => x"000024e1",
			2357 => x"fef824e1",
			2358 => x"000024e1",
			2359 => x"fe6624e1",
			2360 => x"0601151c",
			2361 => x"0207aa14",
			2362 => x"01004308",
			2363 => x"05051004",
			2364 => x"000025a5",
			2365 => x"00f925a5",
			2366 => x"03052f04",
			2367 => x"ff0725a5",
			2368 => x"0b053104",
			2369 => x"003325a5",
			2370 => x"000025a5",
			2371 => x"01005504",
			2372 => x"017925a5",
			2373 => x"000025a5",
			2374 => x"02098130",
			2375 => x"0f089c1c",
			2376 => x"01002d0c",
			2377 => x"02087b04",
			2378 => x"ff4825a5",
			2379 => x"0505f604",
			2380 => x"00e525a5",
			2381 => x"000025a5",
			2382 => x"02092008",
			2383 => x"0504d404",
			2384 => x"000025a5",
			2385 => x"fe7025a5",
			2386 => x"05053c04",
			2387 => x"000025a5",
			2388 => x"ff8125a5",
			2389 => x"06013608",
			2390 => x"09015a04",
			2391 => x"015e25a5",
			2392 => x"000025a5",
			2393 => x"0f091f04",
			2394 => x"fed625a5",
			2395 => x"0f092a04",
			2396 => x"000025a5",
			2397 => x"ffd425a5",
			2398 => x"0705cf14",
			2399 => x"06019410",
			2400 => x"0100e00c",
			2401 => x"020a5b08",
			2402 => x"04173404",
			2403 => x"01e125a5",
			2404 => x"000025a5",
			2405 => x"000025a5",
			2406 => x"000025a5",
			2407 => x"000025a5",
			2408 => x"feb425a5",
			2409 => x"06011f20",
			2410 => x"09008a1c",
			2411 => x"06011208",
			2412 => x"0002dd04",
			2413 => x"02b2265b",
			2414 => x"01bb265b",
			2415 => x"0b04810c",
			2416 => x"03037b04",
			2417 => x"0000265b",
			2418 => x"040da904",
			2419 => x"0000265b",
			2420 => x"01b6265b",
			2421 => x"05051d04",
			2422 => x"ffc1265b",
			2423 => x"fe1c265b",
			2424 => x"fe7f265b",
			2425 => x"0c046318",
			2426 => x"0804ac14",
			2427 => x"03039404",
			2428 => x"fe73265b",
			2429 => x"09004f0c",
			2430 => x"07048008",
			2431 => x"0d04d804",
			2432 => x"0075265b",
			2433 => x"0204265b",
			2434 => x"0000265b",
			2435 => x"fe72265b",
			2436 => x"0388265b",
			2437 => x"040ae820",
			2438 => x"040ae214",
			2439 => x"0d079610",
			2440 => x"05074808",
			2441 => x"0307f404",
			2442 => x"fe6c265b",
			2443 => x"fffa265b",
			2444 => x"05075604",
			2445 => x"04a3265b",
			2446 => x"0000265b",
			2447 => x"fe69265b",
			2448 => x"0a027004",
			2449 => x"feea265b",
			2450 => x"08032004",
			2451 => x"05a0265b",
			2452 => x"fff4265b",
			2453 => x"fe65265b",
			2454 => x"0000265d",
			2455 => x"00002661",
			2456 => x"00002665",
			2457 => x"00002669",
			2458 => x"0000266d",
			2459 => x"00002671",
			2460 => x"00002675",
			2461 => x"00002679",
			2462 => x"0000267d",
			2463 => x"00002681",
			2464 => x"00002685",
			2465 => x"00002689",
			2466 => x"0000268d",
			2467 => x"00002691",
			2468 => x"00002695",
			2469 => x"00002699",
			2470 => x"0000269d",
			2471 => x"000026a1",
			2472 => x"0c046304",
			2473 => x"000026ad",
			2474 => x"fffa26ad",
			2475 => x"07055d04",
			2476 => x"001326b9",
			2477 => x"000026b9",
			2478 => x"07049704",
			2479 => x"000026c5",
			2480 => x"fff126c5",
			2481 => x"06012704",
			2482 => x"000026d9",
			2483 => x"0c050d04",
			2484 => x"ffc326d9",
			2485 => x"000026d9",
			2486 => x"07055d08",
			2487 => x"0b043e04",
			2488 => x"000026ed",
			2489 => x"000f26ed",
			2490 => x"000026ed",
			2491 => x"06012704",
			2492 => x"00002701",
			2493 => x"06015304",
			2494 => x"ff9f2701",
			2495 => x"00002701",
			2496 => x"06013608",
			2497 => x"0600e104",
			2498 => x"00002715",
			2499 => x"00032715",
			2500 => x"00002715",
			2501 => x"06011404",
			2502 => x"00002729",
			2503 => x"06015b04",
			2504 => x"ffc82729",
			2505 => x"00002729",
			2506 => x"06011504",
			2507 => x"0000273d",
			2508 => x"06017c04",
			2509 => x"fff1273d",
			2510 => x"0000273d",
			2511 => x"07055d0c",
			2512 => x"0c052a08",
			2513 => x"0b043e04",
			2514 => x"00002759",
			2515 => x"00132759",
			2516 => x"00002759",
			2517 => x"00002759",
			2518 => x"07055d0c",
			2519 => x"0f062704",
			2520 => x"00002775",
			2521 => x"0c052a04",
			2522 => x"00392775",
			2523 => x"00002775",
			2524 => x"00002775",
			2525 => x"0601270c",
			2526 => x"0600e104",
			2527 => x"00002791",
			2528 => x"06011204",
			2529 => x"001f2791",
			2530 => x"00002791",
			2531 => x"ffd02791",
			2532 => x"0705470c",
			2533 => x"0f05f504",
			2534 => x"000027ad",
			2535 => x"06013604",
			2536 => x"005827ad",
			2537 => x"000027ad",
			2538 => x"000027ad",
			2539 => x"06011404",
			2540 => x"000027c9",
			2541 => x"06015b08",
			2542 => x"06011504",
			2543 => x"000027c9",
			2544 => x"ffd027c9",
			2545 => x"000027c9",
			2546 => x"0705470c",
			2547 => x"06013608",
			2548 => x"0600e204",
			2549 => x"000027ed",
			2550 => x"003427ed",
			2551 => x"000027ed",
			2552 => x"0705ce04",
			2553 => x"fff927ed",
			2554 => x"000027ed",
			2555 => x"06011208",
			2556 => x"0600e104",
			2557 => x"00002811",
			2558 => x"00032811",
			2559 => x"0c045404",
			2560 => x"00002811",
			2561 => x"0b044f04",
			2562 => x"00002811",
			2563 => x"ffbf2811",
			2564 => x"0601360c",
			2565 => x"0f062704",
			2566 => x"0000283d",
			2567 => x"07054704",
			2568 => x"002b283d",
			2569 => x"0000283d",
			2570 => x"04095904",
			2571 => x"0000283d",
			2572 => x"06017804",
			2573 => x"ff6d283d",
			2574 => x"0000283d",
			2575 => x"0c046304",
			2576 => x"00002861",
			2577 => x"0a01df04",
			2578 => x"00002861",
			2579 => x"0f091f08",
			2580 => x"0b063c04",
			2581 => x"ff8a2861",
			2582 => x"00002861",
			2583 => x"00002861",
			2584 => x"07054710",
			2585 => x"0d04cb04",
			2586 => x"00002885",
			2587 => x"06013d08",
			2588 => x"0600e204",
			2589 => x"00002885",
			2590 => x"00102885",
			2591 => x"00002885",
			2592 => x"ffa72885",
			2593 => x"06011204",
			2594 => x"000028a9",
			2595 => x"04097204",
			2596 => x"000028a9",
			2597 => x"0c045404",
			2598 => x"000028a9",
			2599 => x"0b044f04",
			2600 => x"000028a9",
			2601 => x"ff8728a9",
			2602 => x"0f05b604",
			2603 => x"000028cd",
			2604 => x"0c059e0c",
			2605 => x"0f0a1908",
			2606 => x"0705e604",
			2607 => x"002128cd",
			2608 => x"000028cd",
			2609 => x"000028cd",
			2610 => x"000028cd",
			2611 => x"07054710",
			2612 => x"0601360c",
			2613 => x"0600e204",
			2614 => x"000028f9",
			2615 => x"0b043e04",
			2616 => x"000028f9",
			2617 => x"004128f9",
			2618 => x"000028f9",
			2619 => x"0b063c04",
			2620 => x"ffd528f9",
			2621 => x"000028f9",
			2622 => x"0705d114",
			2623 => x"0208ab08",
			2624 => x"06010e04",
			2625 => x"00002925",
			2626 => x"00002925",
			2627 => x"0100e008",
			2628 => x"0006f104",
			2629 => x"00612925",
			2630 => x"00002925",
			2631 => x"00002925",
			2632 => x"00002925",
			2633 => x"06013610",
			2634 => x"0f062704",
			2635 => x"00002959",
			2636 => x"07054708",
			2637 => x"0a024904",
			2638 => x"00472959",
			2639 => x"00002959",
			2640 => x"00002959",
			2641 => x"0b063c08",
			2642 => x"0c043d04",
			2643 => x"00002959",
			2644 => x"ff722959",
			2645 => x"00002959",
			2646 => x"01004b10",
			2647 => x"0c04d10c",
			2648 => x"0d050d04",
			2649 => x"00002995",
			2650 => x"0504f304",
			2651 => x"00002995",
			2652 => x"00642995",
			2653 => x"00002995",
			2654 => x"0d06fc08",
			2655 => x"0600e404",
			2656 => x"00002995",
			2657 => x"ffa62995",
			2658 => x"09016d04",
			2659 => x"00072995",
			2660 => x"00002995",
			2661 => x"06013614",
			2662 => x"0f05e604",
			2663 => x"000029c9",
			2664 => x"0a024c0c",
			2665 => x"07054708",
			2666 => x"0a018404",
			2667 => x"000029c9",
			2668 => x"007a29c9",
			2669 => x"000029c9",
			2670 => x"000029c9",
			2671 => x"06016304",
			2672 => x"fff829c9",
			2673 => x"000029c9",
			2674 => x"0c046304",
			2675 => x"000029f5",
			2676 => x"0600fd04",
			2677 => x"000029f5",
			2678 => x"0601780c",
			2679 => x"06010e04",
			2680 => x"000029f5",
			2681 => x"07046204",
			2682 => x"000029f5",
			2683 => x"ffd429f5",
			2684 => x"000029f5",
			2685 => x"01003614",
			2686 => x"0c047910",
			2687 => x"09002704",
			2688 => x"00002a31",
			2689 => x"0b043d04",
			2690 => x"00002a31",
			2691 => x"01001704",
			2692 => x"00002a31",
			2693 => x"00482a31",
			2694 => x"00002a31",
			2695 => x"06015308",
			2696 => x"06012704",
			2697 => x"00002a31",
			2698 => x"ff5b2a31",
			2699 => x"00002a31",
			2700 => x"0208b40c",
			2701 => x"06010a04",
			2702 => x"00002a6d",
			2703 => x"0a01db04",
			2704 => x"00002a6d",
			2705 => x"ff902a6d",
			2706 => x"0c059e10",
			2707 => x"0100e00c",
			2708 => x"0416b608",
			2709 => x"020a5b04",
			2710 => x"00882a6d",
			2711 => x"00002a6d",
			2712 => x"00002a6d",
			2713 => x"00002a6d",
			2714 => x"00002a6d",
			2715 => x"0208b410",
			2716 => x"06010604",
			2717 => x"00002ab1",
			2718 => x"0a01db04",
			2719 => x"00002ab1",
			2720 => x"01002304",
			2721 => x"00002ab1",
			2722 => x"ff7c2ab1",
			2723 => x"0705e610",
			2724 => x"0100e00c",
			2725 => x"0416b608",
			2726 => x"020a5b04",
			2727 => x"00a82ab1",
			2728 => x"00002ab1",
			2729 => x"00002ab1",
			2730 => x"00002ab1",
			2731 => x"00002ab1",
			2732 => x"0c046314",
			2733 => x"0f05ee04",
			2734 => x"00002afd",
			2735 => x"0900820c",
			2736 => x"07049708",
			2737 => x"0d04cb04",
			2738 => x"00002afd",
			2739 => x"008e2afd",
			2740 => x"00002afd",
			2741 => x"00002afd",
			2742 => x"09014b0c",
			2743 => x"06011204",
			2744 => x"00002afd",
			2745 => x"07046104",
			2746 => x"00002afd",
			2747 => x"ff052afd",
			2748 => x"09016d04",
			2749 => x"00332afd",
			2750 => x"00002afd",
			2751 => x"09006c0c",
			2752 => x"03039404",
			2753 => x"00002b49",
			2754 => x"0704bb04",
			2755 => x"00782b49",
			2756 => x"00002b49",
			2757 => x"06016310",
			2758 => x"00032404",
			2759 => x"00002b49",
			2760 => x"0c044304",
			2761 => x"00002b49",
			2762 => x"06010e04",
			2763 => x"00002b49",
			2764 => x"ff172b49",
			2765 => x"0100e008",
			2766 => x"0100d604",
			2767 => x"00002b49",
			2768 => x"00542b49",
			2769 => x"00002b49",
			2770 => x"0601361c",
			2771 => x"0f070514",
			2772 => x"0601060c",
			2773 => x"01004508",
			2774 => x"01001b04",
			2775 => x"00002b9d",
			2776 => x"00392b9d",
			2777 => x"00002b9d",
			2778 => x"01002a04",
			2779 => x"00002b9d",
			2780 => x"ff902b9d",
			2781 => x"0b05bf04",
			2782 => x"009f2b9d",
			2783 => x"00002b9d",
			2784 => x"0209be08",
			2785 => x"0b063c04",
			2786 => x"ff1b2b9d",
			2787 => x"00002b9d",
			2788 => x"0c051104",
			2789 => x"006a2b9d",
			2790 => x"00002b9d",
			2791 => x"01004718",
			2792 => x"0b047004",
			2793 => x"00002bd9",
			2794 => x"0704aa10",
			2795 => x"03040504",
			2796 => x"00002bd9",
			2797 => x"0c045904",
			2798 => x"00002bd9",
			2799 => x"0504e504",
			2800 => x"00002bd9",
			2801 => x"004a2bd9",
			2802 => x"00002bd9",
			2803 => x"00032404",
			2804 => x"00002bd9",
			2805 => x"ff4f2bd9",
			2806 => x"0601150c",
			2807 => x"0600e604",
			2808 => x"00002c25",
			2809 => x"0c04ee04",
			2810 => x"00772c25",
			2811 => x"00002c25",
			2812 => x"0c050d08",
			2813 => x"00066504",
			2814 => x"ff402c25",
			2815 => x"00002c25",
			2816 => x"0c059e10",
			2817 => x"0e09a20c",
			2818 => x"0003a208",
			2819 => x"00033504",
			2820 => x"00002c25",
			2821 => x"008c2c25",
			2822 => x"00002c25",
			2823 => x"00002c25",
			2824 => x"00002c25",
			2825 => x"01004b14",
			2826 => x"0f061204",
			2827 => x"00002c79",
			2828 => x"0c04980c",
			2829 => x"06012304",
			2830 => x"00e52c79",
			2831 => x"06015704",
			2832 => x"00002c79",
			2833 => x"00042c79",
			2834 => x"00002c79",
			2835 => x"0506b908",
			2836 => x"08024e04",
			2837 => x"00002c79",
			2838 => x"fee72c79",
			2839 => x"09016d0c",
			2840 => x"0c059e08",
			2841 => x"05073904",
			2842 => x"005c2c79",
			2843 => x"00002c79",
			2844 => x"00002c79",
			2845 => x"ffce2c79",
			2846 => x"0b05d718",
			2847 => x"0c052a14",
			2848 => x"0504d504",
			2849 => x"00002cad",
			2850 => x"07055d0c",
			2851 => x"07044e04",
			2852 => x"00002cad",
			2853 => x"09002b04",
			2854 => x"00002cad",
			2855 => x"00232cad",
			2856 => x"00002cad",
			2857 => x"00002cad",
			2858 => x"00002cad",
			2859 => x"0a025718",
			2860 => x"09016d14",
			2861 => x"0f06d908",
			2862 => x"01004304",
			2863 => x"00a62d01",
			2864 => x"ff512d01",
			2865 => x"0002b704",
			2866 => x"00002d01",
			2867 => x"05074804",
			2868 => x"01022d01",
			2869 => x"00002d01",
			2870 => x"ff682d01",
			2871 => x"06012710",
			2872 => x"040c9a04",
			2873 => x"ffec2d01",
			2874 => x"0c049108",
			2875 => x"03037b04",
			2876 => x"00002d01",
			2877 => x"00cb2d01",
			2878 => x"00002d01",
			2879 => x"fe982d01",
			2880 => x"0802dd18",
			2881 => x"07055d10",
			2882 => x"0f05e604",
			2883 => x"00002d65",
			2884 => x"0801e404",
			2885 => x"00002d65",
			2886 => x"0802d504",
			2887 => x"00b92d65",
			2888 => x"00002d65",
			2889 => x"06017804",
			2890 => x"ffc12d65",
			2891 => x"00002d65",
			2892 => x"06011508",
			2893 => x"05051e04",
			2894 => x"005d2d65",
			2895 => x"00002d65",
			2896 => x"0003a204",
			2897 => x"00002d65",
			2898 => x"09004204",
			2899 => x"00002d65",
			2900 => x"0504c904",
			2901 => x"00002d65",
			2902 => x"07046204",
			2903 => x"00002d65",
			2904 => x"fed02d65",
			2905 => x"0208b414",
			2906 => x"06012710",
			2907 => x"02069d04",
			2908 => x"00002db9",
			2909 => x"06010e08",
			2910 => x"01005504",
			2911 => x"00532db9",
			2912 => x"00002db9",
			2913 => x"00002db9",
			2914 => x"ff752db9",
			2915 => x"0100e014",
			2916 => x"0c059e10",
			2917 => x"09002804",
			2918 => x"00002db9",
			2919 => x"0416b608",
			2920 => x"020a5b04",
			2921 => x"00a32db9",
			2922 => x"00002db9",
			2923 => x"00002db9",
			2924 => x"00002db9",
			2925 => x"00002db9",
			2926 => x"06011510",
			2927 => x"0f05e604",
			2928 => x"00002e25",
			2929 => x"01004e08",
			2930 => x"04134d04",
			2931 => x"011f2e25",
			2932 => x"00002e25",
			2933 => x"00002e25",
			2934 => x"0409b30c",
			2935 => x"07053104",
			2936 => x"00002e25",
			2937 => x"0c056104",
			2938 => x"00db2e25",
			2939 => x"00002e25",
			2940 => x"09004210",
			2941 => x"09002b04",
			2942 => x"00002e25",
			2943 => x"0c047508",
			2944 => x"03037b04",
			2945 => x"00002e25",
			2946 => x"00a62e25",
			2947 => x"00002e25",
			2948 => x"0b063c04",
			2949 => x"fead2e25",
			2950 => x"0b065b04",
			2951 => x"00002e25",
			2952 => x"ffd12e25",
			2953 => x"0802f61c",
			2954 => x"0c059e18",
			2955 => x"0f05e604",
			2956 => x"00002e79",
			2957 => x"0100e310",
			2958 => x"0801e404",
			2959 => x"00002e79",
			2960 => x"05075608",
			2961 => x"0003a204",
			2962 => x"008d2e79",
			2963 => x"00002e79",
			2964 => x"00002e79",
			2965 => x"00002e79",
			2966 => x"00002e79",
			2967 => x"06011504",
			2968 => x"00002e79",
			2969 => x"0c045404",
			2970 => x"00002e79",
			2971 => x"09004204",
			2972 => x"00002e79",
			2973 => x"ff172e79",
			2974 => x"09006210",
			2975 => x"0f05b604",
			2976 => x"00002ee5",
			2977 => x"0b04e308",
			2978 => x"0b044004",
			2979 => x"00002ee5",
			2980 => x"00cb2ee5",
			2981 => x"00002ee5",
			2982 => x"08030220",
			2983 => x"0f074610",
			2984 => x"09006c04",
			2985 => x"00002ee5",
			2986 => x"040b3008",
			2987 => x"0600e404",
			2988 => x"00002ee5",
			2989 => x"ff832ee5",
			2990 => x"00002ee5",
			2991 => x"07055d04",
			2992 => x"009d2ee5",
			2993 => x"06017808",
			2994 => x"0f08b804",
			2995 => x"00002ee5",
			2996 => x"ff5c2ee5",
			2997 => x"00002ee5",
			2998 => x"0a025604",
			2999 => x"00002ee5",
			3000 => x"fefb2ee5",
			3001 => x"0601361c",
			3002 => x"07054718",
			3003 => x"0600e104",
			3004 => x"00002f21",
			3005 => x"0a024910",
			3006 => x"0504e404",
			3007 => x"00002f21",
			3008 => x"0a023608",
			3009 => x"0406ea04",
			3010 => x"00002f21",
			3011 => x"006e2f21",
			3012 => x"00002f21",
			3013 => x"00002f21",
			3014 => x"00002f21",
			3015 => x"ffb32f21",
			3016 => x"06012728",
			3017 => x"01003f0c",
			3018 => x"0f05b604",
			3019 => x"00002fad",
			3020 => x"0c047b04",
			3021 => x"01572fad",
			3022 => x"00002fad",
			3023 => x"0e04f00c",
			3024 => x"06010604",
			3025 => x"00002fad",
			3026 => x"040bff04",
			3027 => x"febc2fad",
			3028 => x"00002fad",
			3029 => x"0002b304",
			3030 => x"00002fad",
			3031 => x"0e050704",
			3032 => x"00002fad",
			3033 => x"0100a104",
			3034 => x"01292fad",
			3035 => x"00002fad",
			3036 => x"0003a214",
			3037 => x"040a950c",
			3038 => x"0e082c08",
			3039 => x"0307f404",
			3040 => x"ff502fad",
			3041 => x"00bb2fad",
			3042 => x"fec02fad",
			3043 => x"0c057e04",
			3044 => x"013e2fad",
			3045 => x"ffa62fad",
			3046 => x"01002308",
			3047 => x"09002f04",
			3048 => x"ffc02fad",
			3049 => x"00002fad",
			3050 => x"fe792fad",
			3051 => x"09006210",
			3052 => x"0f05b604",
			3053 => x"00003021",
			3054 => x"0b04e308",
			3055 => x"0b044004",
			3056 => x"00003021",
			3057 => x"00bd3021",
			3058 => x"00003021",
			3059 => x"08030224",
			3060 => x"040a9518",
			3061 => x"0409720c",
			3062 => x"0f074904",
			3063 => x"00003021",
			3064 => x"0506f104",
			3065 => x"00943021",
			3066 => x"00003021",
			3067 => x"09007b04",
			3068 => x"00003021",
			3069 => x"0f097d04",
			3070 => x"ff253021",
			3071 => x"00003021",
			3072 => x"0c056308",
			3073 => x"0f076d04",
			3074 => x"00003021",
			3075 => x"00993021",
			3076 => x"00003021",
			3077 => x"0a025604",
			3078 => x"00003021",
			3079 => x"ff053021",
			3080 => x"0c046320",
			3081 => x"09005d10",
			3082 => x"0f05b604",
			3083 => x"ff6930ad",
			3084 => x"04143608",
			3085 => x"06013504",
			3086 => x"018330ad",
			3087 => x"000030ad",
			3088 => x"040a30ad",
			3089 => x"0e04a008",
			3090 => x"01003c04",
			3091 => x"000030ad",
			3092 => x"fead30ad",
			3093 => x"06012004",
			3094 => x"015a30ad",
			3095 => x"ffbe30ad",
			3096 => x"0003a21c",
			3097 => x"0c059e18",
			3098 => x"0c04ed0c",
			3099 => x"09008408",
			3100 => x"0d052604",
			3101 => x"000030ad",
			3102 => x"00ef30ad",
			3103 => x"fefd30ad",
			3104 => x"08024104",
			3105 => x"000030ad",
			3106 => x"0100e304",
			3107 => x"01a430ad",
			3108 => x"000030ad",
			3109 => x"fea330ad",
			3110 => x"06010e04",
			3111 => x"000030ad",
			3112 => x"0b045e04",
			3113 => x"000030ad",
			3114 => x"fe6e30ad",
			3115 => x"0100451c",
			3116 => x"0f05e608",
			3117 => x"0600fd04",
			3118 => x"00003139",
			3119 => x"ff8a3139",
			3120 => x"0c049910",
			3121 => x"01003608",
			3122 => x"0d04cb04",
			3123 => x"00003139",
			3124 => x"019f3139",
			3125 => x"0d050f04",
			3126 => x"ffeb3139",
			3127 => x"00c73139",
			3128 => x"00003139",
			3129 => x"0003a21c",
			3130 => x"0a025314",
			3131 => x"0c04f110",
			3132 => x"00032c08",
			3133 => x"0f064a04",
			3134 => x"00003139",
			3135 => x"00d73139",
			3136 => x"0d055904",
			3137 => x"00003139",
			3138 => x"ff683139",
			3139 => x"fed53139",
			3140 => x"0c058104",
			3141 => x"013e3139",
			3142 => x"ffcf3139",
			3143 => x"05050304",
			3144 => x"00003139",
			3145 => x"09007104",
			3146 => x"00003139",
			3147 => x"0a023004",
			3148 => x"00003139",
			3149 => x"fe823139",
			3150 => x"0a025720",
			3151 => x"09016d1c",
			3152 => x"0f06d908",
			3153 => x"01004304",
			3154 => x"009631b5",
			3155 => x"ff6531b5",
			3156 => x"0002b704",
			3157 => x"000031b5",
			3158 => x"0507480c",
			3159 => x"0a023604",
			3160 => x"010231b5",
			3161 => x"0802d404",
			3162 => x"000031b5",
			3163 => x"003931b5",
			3164 => x"000031b5",
			3165 => x"ff7931b5",
			3166 => x"09005d18",
			3167 => x"06012710",
			3168 => x"0704920c",
			3169 => x"0f05c304",
			3170 => x"000031b5",
			3171 => x"040d8804",
			3172 => x"000031b5",
			3173 => x"00a931b5",
			3174 => x"000031b5",
			3175 => x"0f068704",
			3176 => x"fffd31b5",
			3177 => x"000031b5",
			3178 => x"0504d704",
			3179 => x"000031b5",
			3180 => x"fe9a31b5",
			3181 => x"06011f1c",
			3182 => x"01005318",
			3183 => x"06011510",
			3184 => x"0c04930c",
			3185 => x"0f05d204",
			3186 => x"00673241",
			3187 => x"09007b04",
			3188 => x"01e73241",
			3189 => x"00003241",
			3190 => x"03b53241",
			3191 => x"02088b04",
			3192 => x"fe2d3241",
			3193 => x"01be3241",
			3194 => x"fe763241",
			3195 => x"07046c0c",
			3196 => x"02089304",
			3197 => x"fe6d3241",
			3198 => x"0f06ed04",
			3199 => x"026c3241",
			3200 => x"01273241",
			3201 => x"0a023310",
			3202 => x"0b064b0c",
			3203 => x"0b059704",
			3204 => x"fec73241",
			3205 => x"02092e04",
			3206 => x"09b43241",
			3207 => x"ff983241",
			3208 => x"fe693241",
			3209 => x"0c04540c",
			3210 => x"03042608",
			3211 => x"03037b04",
			3212 => x"feb83241",
			3213 => x"01753241",
			3214 => x"fe753241",
			3215 => x"fe693241",
			3216 => x"06012724",
			3217 => x"01004510",
			3218 => x"0f05b604",
			3219 => x"ff2432d5",
			3220 => x"0704a908",
			3221 => x"06011504",
			3222 => x"019532d5",
			3223 => x"00ad32d5",
			3224 => x"000032d5",
			3225 => x"0f070f08",
			3226 => x"09007304",
			3227 => x"000032d5",
			3228 => x"fe9132d5",
			3229 => x"03071b08",
			3230 => x"0f074904",
			3231 => x"000032d5",
			3232 => x"01ec32d5",
			3233 => x"ff7e32d5",
			3234 => x"0409c70c",
			3235 => x"00033504",
			3236 => x"feb732d5",
			3237 => x"0e07dc04",
			3238 => x"000032d5",
			3239 => x"012032d5",
			3240 => x"07046c18",
			3241 => x"09004f14",
			3242 => x"0d04e60c",
			3243 => x"07046808",
			3244 => x"0d04d804",
			3245 => x"ffce32d5",
			3246 => x"000032d5",
			3247 => x"000032d5",
			3248 => x"01001c04",
			3249 => x"000032d5",
			3250 => x"008232d5",
			3251 => x"ff2732d5",
			3252 => x"fe7e32d5",
			3253 => x"01003610",
			3254 => x"0f05ee04",
			3255 => x"00003359",
			3256 => x"05059508",
			3257 => x"0d04d804",
			3258 => x"00003359",
			3259 => x"010d3359",
			3260 => x"00003359",
			3261 => x"0003c428",
			3262 => x"040a951c",
			3263 => x"04097210",
			3264 => x"0f061204",
			3265 => x"00003359",
			3266 => x"07054708",
			3267 => x"0801e404",
			3268 => x"00003359",
			3269 => x"00d53359",
			3270 => x"00003359",
			3271 => x"0705ce08",
			3272 => x"01004e04",
			3273 => x"00003359",
			3274 => x"fee83359",
			3275 => x"00003359",
			3276 => x"0c056408",
			3277 => x"0003ab04",
			3278 => x"00de3359",
			3279 => x"00003359",
			3280 => x"00003359",
			3281 => x"06011204",
			3282 => x"00003359",
			3283 => x"0504d504",
			3284 => x"00003359",
			3285 => x"feb63359",
			3286 => x"01003614",
			3287 => x"01001b04",
			3288 => x"000033cd",
			3289 => x"0c04790c",
			3290 => x"0f05b604",
			3291 => x"000033cd",
			3292 => x"0d04cb04",
			3293 => x"000033cd",
			3294 => x"017133cd",
			3295 => x"000033cd",
			3296 => x"0802f620",
			3297 => x"0c059e1c",
			3298 => x"0e04c908",
			3299 => x"040af504",
			3300 => x"ff3c33cd",
			3301 => x"000033cd",
			3302 => x"0100e010",
			3303 => x"0705ce08",
			3304 => x"06012804",
			3305 => x"00f533cd",
			3306 => x"ff7b33cd",
			3307 => x"0100d604",
			3308 => x"000033cd",
			3309 => x"014233cd",
			3310 => x"000033cd",
			3311 => x"ff4133cd",
			3312 => x"06011504",
			3313 => x"000033cd",
			3314 => x"fe8533cd",
			3315 => x"01003610",
			3316 => x"0f061204",
			3317 => x"00003451",
			3318 => x"05059508",
			3319 => x"0d04d804",
			3320 => x"00003451",
			3321 => x"01243451",
			3322 => x"00003451",
			3323 => x"0003c428",
			3324 => x"09016d1c",
			3325 => x"09014b14",
			3326 => x"06012810",
			3327 => x"0e04a008",
			3328 => x"0d054104",
			3329 => x"ffd23451",
			3330 => x"00003451",
			3331 => x"05064204",
			3332 => x"00b93451",
			3333 => x"00003451",
			3334 => x"ff353451",
			3335 => x"0d079604",
			3336 => x"00e03451",
			3337 => x"00003451",
			3338 => x"0a027004",
			3339 => x"ff303451",
			3340 => x"0901b204",
			3341 => x"00333451",
			3342 => x"00003451",
			3343 => x"06011204",
			3344 => x"00003451",
			3345 => x"0504d504",
			3346 => x"00003451",
			3347 => x"feaf3451",
			3348 => x"06011f20",
			3349 => x"0900821c",
			3350 => x"0f05c308",
			3351 => x"07045104",
			3352 => x"000934dd",
			3353 => x"fe6a34dd",
			3354 => x"02071704",
			3355 => x"042434dd",
			3356 => x"0c047e0c",
			3357 => x"06011904",
			3358 => x"020834dd",
			3359 => x"02088b04",
			3360 => x"fea734dd",
			3361 => x"020834dd",
			3362 => x"fe9334dd",
			3363 => x"fe6c34dd",
			3364 => x"07046c0c",
			3365 => x"02089304",
			3366 => x"fe6934dd",
			3367 => x"0f06ed04",
			3368 => x"02ce34dd",
			3369 => x"015934dd",
			3370 => x"0c043a08",
			3371 => x"08046904",
			3372 => x"ff8d34dd",
			3373 => x"008834dd",
			3374 => x"040ae810",
			3375 => x"040ae204",
			3376 => x"fe8634dd",
			3377 => x"0802f304",
			3378 => x"feb234dd",
			3379 => x"08030204",
			3380 => x"058b34dd",
			3381 => x"fef434dd",
			3382 => x"fe6634dd",
			3383 => x"01003c18",
			3384 => x"0c049914",
			3385 => x"03039408",
			3386 => x"07044a04",
			3387 => x"00003559",
			3388 => x"ff773559",
			3389 => x"04143608",
			3390 => x"0207df04",
			3391 => x"002f3559",
			3392 => x"016b3559",
			3393 => x"036a3559",
			3394 => x"fefe3559",
			3395 => x"0802f424",
			3396 => x"0c059e20",
			3397 => x"0e05c30c",
			3398 => x"09007f08",
			3399 => x"0304af04",
			3400 => x"ff1a3559",
			3401 => x"01083559",
			3402 => x"fed33559",
			3403 => x"0100e010",
			3404 => x"00034608",
			3405 => x"0b05a604",
			3406 => x"01843559",
			3407 => x"fedb3559",
			3408 => x"02088504",
			3409 => x"00003559",
			3410 => x"01d63559",
			3411 => x"00003559",
			3412 => x"fea83559",
			3413 => x"fe773559",
			3414 => x"06011920",
			3415 => x"0505f61c",
			3416 => x"0207670c",
			3417 => x"0304d804",
			3418 => x"fe9c35fd",
			3419 => x"01005904",
			3420 => x"017335fd",
			3421 => x"000035fd",
			3422 => x"0100530c",
			3423 => x"01004504",
			3424 => x"01aa35fd",
			3425 => x"06011204",
			3426 => x"01a035fd",
			3427 => x"000035fd",
			3428 => x"ffae35fd",
			3429 => x"fe9235fd",
			3430 => x"09004f10",
			3431 => x"020a500c",
			3432 => x"0414a408",
			3433 => x"02088b04",
			3434 => x"fea735fd",
			3435 => x"018935fd",
			3436 => x"fe8235fd",
			3437 => x"08ee35fd",
			3438 => x"0409c710",
			3439 => x"08028704",
			3440 => x"fe7e35fd",
			3441 => x"0e07dc04",
			3442 => x"ff3c35fd",
			3443 => x"0901bc04",
			3444 => x"028435fd",
			3445 => x"ffbb35fd",
			3446 => x"0802f410",
			3447 => x"0901830c",
			3448 => x"02099d08",
			3449 => x"040b2404",
			3450 => x"fe8b35fd",
			3451 => x"000035fd",
			3452 => x"021735fd",
			3453 => x"fe7635fd",
			3454 => x"fe6735fd",
			3455 => x"0601272c",
			3456 => x"02081520",
			3457 => x"0a022b18",
			3458 => x"0f05e604",
			3459 => x"ff4e3691",
			3460 => x"01009910",
			3461 => x"0a01f708",
			3462 => x"0801e404",
			3463 => x"00003691",
			3464 => x"01b63691",
			3465 => x"07049704",
			3466 => x"00f63691",
			3467 => x"ff693691",
			3468 => x"ffd63691",
			3469 => x"06010e04",
			3470 => x"002d3691",
			3471 => x"fe943691",
			3472 => x"0704aa08",
			3473 => x"01004b04",
			3474 => x"01903691",
			3475 => x"00003691",
			3476 => x"ff323691",
			3477 => x"02090004",
			3478 => x"fe6f3691",
			3479 => x"0c059e18",
			3480 => x"0003a210",
			3481 => x"0b063c08",
			3482 => x"0f090504",
			3483 => x"008c3691",
			3484 => x"ff6a3691",
			3485 => x"0b065b04",
			3486 => x"014b3691",
			3487 => x"00003691",
			3488 => x"0b049f04",
			3489 => x"008c3691",
			3490 => x"feae3691",
			3491 => x"fe8b3691",
			3492 => x"06011f24",
			3493 => x"01004b18",
			3494 => x"02071704",
			3495 => x"06dd3735",
			3496 => x"01001504",
			3497 => x"fe753735",
			3498 => x"0207f808",
			3499 => x"06011504",
			3500 => x"02e63735",
			3501 => x"fdcf3735",
			3502 => x"03058704",
			3503 => x"02c03735",
			3504 => x"03c93735",
			3505 => x"01005108",
			3506 => x"01004f04",
			3507 => x"feca3735",
			3508 => x"00b83735",
			3509 => x"fe673735",
			3510 => x"07046c0c",
			3511 => x"02089304",
			3512 => x"fe613735",
			3513 => x"0a02ed04",
			3514 => x"04573735",
			3515 => x"02d13735",
			3516 => x"04085204",
			3517 => x"04203735",
			3518 => x"040ae810",
			3519 => x"0705e60c",
			3520 => x"0d06d404",
			3521 => x"fe613735",
			3522 => x"0802cf04",
			3523 => x"032b3735",
			3524 => x"10983735",
			3525 => x"fe603735",
			3526 => x"0505000c",
			3527 => x"0d04f404",
			3528 => x"fe7f3735",
			3529 => x"0504e704",
			3530 => x"00b93735",
			3531 => x"fed53735",
			3532 => x"fe5e3735",
			3533 => x"06011f1c",
			3534 => x"09008a18",
			3535 => x"0207aa0c",
			3536 => x"06010e08",
			3537 => x"0304d604",
			3538 => x"003d37c9",
			3539 => x"01c837c9",
			3540 => x"fe6d37c9",
			3541 => x"0c047e08",
			3542 => x"06011904",
			3543 => x"01af37c9",
			3544 => x"00dc37c9",
			3545 => x"004a37c9",
			3546 => x"fe9737c9",
			3547 => x"04085204",
			3548 => x"043037c9",
			3549 => x"0003a214",
			3550 => x"0c059e10",
			3551 => x"0f089c04",
			3552 => x"feb637c9",
			3553 => x"0100e308",
			3554 => x"06013504",
			3555 => x"000037c9",
			3556 => x"031737c9",
			3557 => x"fee537c9",
			3558 => x"fe6d37c9",
			3559 => x"07046c08",
			3560 => x"02089304",
			3561 => x"fe8737c9",
			3562 => x"014337c9",
			3563 => x"0c04540c",
			3564 => x"0e037908",
			3565 => x"0d04ce04",
			3566 => x"ff7237c9",
			3567 => x"00a537c9",
			3568 => x"fef137c9",
			3569 => x"fe6637c9",
			3570 => x"06011f20",
			3571 => x"01004b1c",
			3572 => x"0f05c308",
			3573 => x"07045104",
			3574 => x"00033875",
			3575 => x"fe7a3875",
			3576 => x"06011508",
			3577 => x"0408cc04",
			3578 => x"03443875",
			3579 => x"01f33875",
			3580 => x"07048f08",
			3581 => x"040c9a04",
			3582 => x"ffe43875",
			3583 => x"01f03875",
			3584 => x"fdf73875",
			3585 => x"fe6d3875",
			3586 => x"07046c0c",
			3587 => x"0f05ee04",
			3588 => x"fe6d3875",
			3589 => x"01002d04",
			3590 => x"02803875",
			3591 => x"fe913875",
			3592 => x"0c043a08",
			3593 => x"08046904",
			3594 => x"ffa13875",
			3595 => x"00713875",
			3596 => x"040ae818",
			3597 => x"040ae20c",
			3598 => x"0c059e08",
			3599 => x"0c057f04",
			3600 => x"fe983875",
			3601 => x"01db3875",
			3602 => x"fe653875",
			3603 => x"0c057e08",
			3604 => x"0c04b404",
			3605 => x"ff193875",
			3606 => x"04b73875",
			3607 => x"feb33875",
			3608 => x"0c045e08",
			3609 => x"0c045c04",
			3610 => x"fe863875",
			3611 => x"02103875",
			3612 => x"fe633875",
			3613 => x"0c046328",
			3614 => x"0f05b604",
			3615 => x"fe5f3963",
			3616 => x"01003f14",
			3617 => x"02080e0c",
			3618 => x"0a028e04",
			3619 => x"030e3963",
			3620 => x"0004b804",
			3621 => x"fea23963",
			3622 => x"003c3963",
			3623 => x"0006ad04",
			3624 => x"032b3963",
			3625 => x"048c3963",
			3626 => x"0a025608",
			3627 => x"05051e04",
			3628 => x"039b3963",
			3629 => x"00383963",
			3630 => x"040d5504",
			3631 => x"fe563963",
			3632 => x"00b63963",
			3633 => x"07048f1c",
			3634 => x"0a024c08",
			3635 => x"0207c504",
			3636 => x"00a63963",
			3637 => x"03273963",
			3638 => x"02087e0c",
			3639 => x"0b045f08",
			3640 => x"0504d604",
			3641 => x"fe9a3963",
			3642 => x"00763963",
			3643 => x"fe613963",
			3644 => x"01003c04",
			3645 => x"03003963",
			3646 => x"fe913963",
			3647 => x"02076714",
			3648 => x"09006f08",
			3649 => x"040c4404",
			3650 => x"04ad3963",
			3651 => x"ff103963",
			3652 => x"0f067a04",
			3653 => x"fe583963",
			3654 => x"05066c04",
			3655 => x"04d03963",
			3656 => x"fe8d3963",
			3657 => x"0802d514",
			3658 => x"0705e610",
			3659 => x"02089008",
			3660 => x"0a01f704",
			3661 => x"01e63963",
			3662 => x"fed13963",
			3663 => x"0d073004",
			3664 => x"0d0b3963",
			3665 => x"00913963",
			3666 => x"fe5f3963",
			3667 => x"0d04e608",
			3668 => x"0504f204",
			3669 => x"fea13963",
			3670 => x"001c3963",
			3671 => x"fe5d3963",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1192, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(2454, initial_addr_3'length));
	end generate gen_rom_15;

	process (Clk)
	begin
		if rising_edge(Clk) then
			if (Re = '1') then
				-- Read from Addr
				Dout <= bank(to_integer(unsigned(Addr)));
			else
				Dout <= (others => '0');
			end if;
		end if;
	end process;
end Behavioral;
