-------------------------------------------------------------------------------
-- Synchronous ROM with generic memory and data sizes
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity rom is
    generic(ADDRESS_BITS: positive;
            DATA_LENGTH:  positive;
            SELECT_ROM:  integer := 0); -- Select which ROM to use
    port(-- Control signals
         Clk: in std_logic;
         Re:  in std_logic;
         
         -- Input signals
         Addr: in std_logic_vector (ADDRESS_BITS - 1 downto 0);
         
         -- Output
         Dout: out std_logic_vector (DATA_LENGTH - 1 downto 0);
         initial_addr_2: out std_logic_vector (ADDRESS_BITS - 1 downto 0);
         initial_addr_3: out std_logic_vector (ADDRESS_BITS - 1 downto 0));
end rom;

architecture Behavioral of rom is

    type MemoryBank is array(0 to 2**ADDRESS_BITS - 1)
                    of std_logic_vector(DATA_LENGTH - 1 downto 0);
    signal bank: MemoryBank;


begin

	gen_rom_0: if SELECT_ROM = 0 generate
		bank <= (
			0 => "00000000000000000000000000000101",
			1 => "00000000000000000000000000001001",
			2 => "00000000000000000000000000001101",
			3 => "00000000000000000000000000010001",
			4 => "00000000000000000000000000010101",
			5 => "00000000000000000000000000011001",
			6 => "00000000000000000000000000011101",
			7 => "00000000000000000000000000100001",
			8 => "00000000000000000000000000100101",
			9 => "00000000000000000000000000101001",
			10 => "00000000000000000000000000101101",
			11 => "00000000000000000000000000110001",
			12 => "00000000000000000000000000110101",
			13 => "00000000000000000000000000111001",
			14 => "00000000000000000000000000111101",
			15 => "00000000000000000000000001000001",
			16 => "00000000000000000000000001000101",
			17 => "00000000000000000000000001001001",
			18 => "00000000000000000000000001001101",
			19 => "00000000000000000000000001010001",
			20 => "00000000000000000000000001010101",
			21 => "00000000000000000000000001011001",
			22 => "00000000000000000000000001011101",
			23 => "00000000000000000000000001100001",
			24 => "00000000000000000000000001100101",
			25 => "00000000000000000000000001101001",
			26 => "00000000000000000000000001101101",
			27 => "00000000000000000000000001110001",
			28 => "00000000000000000000000001110101",
			29 => "00000000000000000000000001111001",
			30 => "00000000000000000000000001111101",
			31 => "00000000000000000000000010000001",
			32 => "00000000000000000000000010000101",
			33 => "00000000000000000000000010001001",
			34 => "00000000000000000000000010001101",
			35 => "00000000000000000000000010010001",
			36 => "00000000000000000000000010010101",
			37 => "0000001111000000001010111000000100",
			38 => "00000000000000000000000010100001",
			39 => "11111111111001100000000010100001",
			40 => "0000001111000000000000001100000100",
			41 => "00000000000000000000000010101101",
			42 => "11111111111100100000000010101101",
			43 => "0000000000000000001100100100000100",
			44 => "11111111111001110000000010111001",
			45 => "00000000000000000000000010111001",
			46 => "0000000000000000001100100100000100",
			47 => "11111111111011010000000011000101",
			48 => "00000000000000000000000011000101",
			49 => "0000001111000000000000001100000100",
			50 => "00000000000000000000000011010001",
			51 => "11111111111011100000000011010001",
			52 => "0000001111000000000111001000001000",
			53 => "0000001110000000001001101000000100",
			54 => "00000000000000000000000011100101",
			55 => "00000000000011100000000011100101",
			56 => "11111111111000010000000011100101",
			57 => "0000000000000000000110100000001000",
			58 => "0000001111000000001100101100000100",
			59 => "00000000000000000000000100000001",
			60 => "11111111100110010000000100000001",
			61 => "0000001110000000001001101000000100",
			62 => "00000000000000000000000100000001",
			63 => "00000000000101100000000100000001",
			64 => "0000000000000000000101100100000100",
			65 => "11111111000011000000000100011101",
			66 => "0000000110000000001100011000001000",
			67 => "0000001001000000001100100000000100",
			68 => "00000000011111110000000100011101",
			69 => "00000000000000000000000100011101",
			70 => "00000000000000000000000100011101",
			71 => "0000001001000000001100100000001100",
			72 => "0000000110000000001100011000001000",
			73 => "0000000101000000000100011000000100",
			74 => "00000000000000000000000100111001",
			75 => "00000000100010000000000100111001",
			76 => "00000000000000000000000100111001",
			77 => "11111111001100100000000100111001",
			78 => "0000000001000000001110011100001100",
			79 => "0000001110000000001100011100000100",
			80 => "00000000000000000000000101010101",
			81 => "0000001111000000001010111000000100",
			82 => "00000000000010110000000101010101",
			83 => "00000000000000000000000101010101",
			84 => "00000000000000000000000101010101",
			85 => "0000001111000000001010111000001100",
			86 => "0000001100000000001110001100000100",
			87 => "00000000000000000000000101110001",
			88 => "0000001100000000001101010100000100",
			89 => "00000000001000110000000101110001",
			90 => "00000000000000000000000101110001",
			91 => "00000000000000000000000101110001",
			92 => "0000001111000000001010111000001100",
			93 => "0000001100000000001101010100001000",
			94 => "0000001100000000001100110000000100",
			95 => "00000000000000000000000110001101",
			96 => "00000000000111100000000110001101",
			97 => "00000000000000000000000110001101",
			98 => "00000000000000000000000110001101",
			99 => "0000001001000000001100100000001100",
			100 => "0000001111000000001010111000001000",
			101 => "0000000000000000000101100100000100",
			102 => "00000000000000000000000110101001",
			103 => "00000000000001100000000110101001",
			104 => "00000000000000000000000110101001",
			105 => "00000000000000000000000110101001",
			106 => "0000000000000000000110100000001000",
			107 => "0000001001000000001100100000000100",
			108 => "00000000000000000000000111001101",
			109 => "11111110110001010000000111001101",
			110 => "0000001100000000000100001000001000",
			111 => "0000000010000000001110110100000100",
			112 => "00000000110011110000000111001101",
			113 => "00000000000000000000000111001101",
			114 => "00000000000000000000000111001101",
			115 => "0000000100000000000010100000000100",
			116 => "11111110100100110000000111110001",
			117 => "0000000010000000001110010000001100",
			118 => "0000000011000000000001110100000100",
			119 => "00000000000000000000000111110001",
			120 => "0000001001000000001100100000000100",
			121 => "00000001001100010000000111110001",
			122 => "00000000000000000000000111110001",
			123 => "00000000000000000000000111110001",
			124 => "0000000001000000001110011100010000",
			125 => "0000001100000000001101010100001100",
			126 => "0000000101000000001110110000000100",
			127 => "00000000000000000000001000010101",
			128 => "0000001111000000001010111000000100",
			129 => "00000000011101010000001000010101",
			130 => "00000000000000000000001000010101",
			131 => "00000000000000000000001000010101",
			132 => "11111111001000000000001000010101",
			133 => "0000001111000000001010111000010000",
			134 => "0000000111000000000111001000001100",
			135 => "0000001100000000001100110000000100",
			136 => "00000000000000000000001000111001",
			137 => "0000001001000000001100100000000100",
			138 => "00000000011000100000001000111001",
			139 => "00000000000000000000001000111001",
			140 => "00000000000000000000001000111001",
			141 => "11111111011000100000001000111001",
			142 => "0000000001000000001110011100010000",
			143 => "0000001100000000000001111100001100",
			144 => "0000000111000000000110000100000100",
			145 => "00000000000000000000001001011101",
			146 => "0000001111000000001010111000000100",
			147 => "00000000001011010000001001011101",
			148 => "00000000000000000000001001011101",
			149 => "00000000000000000000001001011101",
			150 => "11111111101111000000001001011101",
			151 => "0000001111000000000111001000010000",
			152 => "0000001110000000001001101000000100",
			153 => "00000000000000000000001010000001",
			154 => "0000001001000000001100100000001000",
			155 => "0000001100000000001101010100000100",
			156 => "00000000001001010000001010000001",
			157 => "00000000000000000000001010000001",
			158 => "00000000000000000000001010000001",
			159 => "11111111110110010000001010000001",
			160 => "0000001001000000001100100000010000",
			161 => "0000001100000000001110001100000100",
			162 => "00000000000000000000001010100101",
			163 => "0000001100000000001101010100001000",
			164 => "0000001111000000000111001000000100",
			165 => "00000000001010100000001010100101",
			166 => "00000000000000000000001010100101",
			167 => "00000000000000000000001010100101",
			168 => "00000000000000000000001010100101",
			169 => "0000000000000000000010110100001000",
			170 => "0000001001000000001100100000000100",
			171 => "00000000000000000000001011010001",
			172 => "11111111100001010000001011010001",
			173 => "0000001110000000001001101000000100",
			174 => "00000000000000000000001011010001",
			175 => "0000001100000000001101010100001000",
			176 => "0000001001000000001100100000000100",
			177 => "00000000010000010000001011010001",
			178 => "00000000000000000000001011010001",
			179 => "00000000000000000000001011010001",
			180 => "0000000000000000000101100100000100",
			181 => "11111110011011010000001011111101",
			182 => "0000000001000000001110011100001100",
			183 => "0000001111000000000111001000001000",
			184 => "0000000010000000001001100000000100",
			185 => "00000001011011010000001011111101",
			186 => "00000000000000000000001011111101",
			187 => "00000000000000000000001011111101",
			188 => "0000001111000000000000001100000100",
			189 => "00000000010000110000001011111101",
			190 => "11111111001100100000001011111101",
			191 => "0000000000000000001101000100001100",
			192 => "0000000001000000001110011100001000",
			193 => "0000001110000000001011010100000100",
			194 => "11111110101001010000001100110001",
			195 => "00000001101110100000001100110001",
			196 => "11111110011001100000001100110001",
			197 => "0000000010000000001100010100000100",
			198 => "00000001101000100000001100110001",
			199 => "0000000100000000000001100000000100",
			200 => "11111110100001100000001100110001",
			201 => "0000000010000000001110110100000100",
			202 => "00000001111001010000001100110001",
			203 => "11111111100001110000001100110001",
			204 => "0000000000000000001100100100001100",
			205 => "0000001001000000001100100000001000",
			206 => "0000000011000000000111000000000100",
			207 => "11111110011011000000001101101101",
			208 => "00000100101000110000001101101101",
			209 => "11111110010111010000001101101101",
			210 => "0000000010000000000110010000001100",
			211 => "0000001111000000001010111100001000",
			212 => "0000001111000000000100001000000100",
			213 => "00000010111000110000001101101101",
			214 => "00000001110110000000001101101101",
			215 => "00000101001110100000001101101101",
			216 => "0000000111000000001101010100000100",
			217 => "00000001110010100000001101101101",
			218 => "11111110010010010000001101101101",
			219 => "0000000000000000000010110100001000",
			220 => "0000001001000000001100100000000100",
			221 => "00000000000000000000001110100001",
			222 => "11111110011010000000001110100001",
			223 => "0000001111000000000000001100000100",
			224 => "00000001100101110000001110100001",
			225 => "0000000110000000001100011000001000",
			226 => "0000000010000000000010000100000100",
			227 => "00000001101010100000001110100001",
			228 => "00000000000000000000001110100001",
			229 => "0000001010000000000010111100000100",
			230 => "11111110100110010000001110100001",
			231 => "00000001000011000000001110100001",
			232 => "0000000000000000000010110100001000",
			233 => "0000001001000000001100100000000100",
			234 => "00000000000000000000001111011101",
			235 => "11111110011101000000001111011101",
			236 => "0000001100000000000100001000001100",
			237 => "0000000010000000001110110100001000",
			238 => "0000000000000000000110100000000100",
			239 => "00000000000000000000001111011101",
			240 => "00000001110101100000001111011101",
			241 => "00000000000000000000001111011101",
			242 => "0000000010000000000011001000000100",
			243 => "00000000110001000000001111011101",
			244 => "0000000110000000001100011000000100",
			245 => "00000000000000000000001111011101",
			246 => "11111111011010000000001111011101",
			247 => "0000001000000000000101101100001000",
			248 => "0000001001000000001100100000000100",
			249 => "00000000000000000000010000010001",
			250 => "11111110011001110000010000010001",
			251 => "0000000010000000001100010100000100",
			252 => "00000001100110010000010000010001",
			253 => "0000000110000000001100011000000100",
			254 => "00000001111101010000010000010001",
			255 => "0000001010000000000010111100001000",
			256 => "0000001011000000001010111100000100",
			257 => "00000000000000000000010000010001",
			258 => "11111110100000100000010000010001",
			259 => "00000000111100110000010000010001",
			260 => "0000000000000000000110100000001000",
			261 => "0000001111000000000000001100000100",
			262 => "00000000000000000000010001000101",
			263 => "11111111010110010000010001000101",
			264 => "0000000111000000000111001000010000",
			265 => "0000001111000000000111001000001100",
			266 => "0000001001000000001100100000000100",
			267 => "00000000000000000000010001000101",
			268 => "0000001001000000001100100000000100",
			269 => "00000000010011100000010001000101",
			270 => "00000000000000000000010001000101",
			271 => "00000000000000000000010001000101",
			272 => "00000000000000000000010001000101",
			273 => "0000000000000000000010110100001000",
			274 => "0000001001000000001100100000000100",
			275 => "00000000000000000000010001111001",
			276 => "11111111011111000000010001111001",
			277 => "0000001110000000001001101000000100",
			278 => "00000000000000000000010001111001",
			279 => "0000001100000000001101010100001100",
			280 => "0000001111000000000111001000001000",
			281 => "0000001001000000001100100000000100",
			282 => "00000000010010110000010001111001",
			283 => "00000000000000000000010001111001",
			284 => "00000000000000000000010001111001",
			285 => "00000000000000000000010001111001",
			286 => "0000001001000000001100100000010100",
			287 => "0000000111000000000111001000010000",
			288 => "0000000101000000001110110000000100",
			289 => "00000000000000000000010010100101",
			290 => "0000001111000000001010111000001000",
			291 => "0000001011000000001110110000000100",
			292 => "00000000010100110000010010100101",
			293 => "00000000000000000000010010100101",
			294 => "00000000000000000000010010100101",
			295 => "00000000000000000000010010100101",
			296 => "11111111010001100000010010100101",
			297 => "0000001111000000001010111000010100",
			298 => "0000001110000000001001101000000100",
			299 => "00000000000000000000010011010001",
			300 => "0000001100000000001101010100001100",
			301 => "0000000001000000001110011100001000",
			302 => "0000000001000000001110011100000100",
			303 => "00000000000000000000010011010001",
			304 => "00000000001001010000010011010001",
			305 => "00000000000000000000010011010001",
			306 => "00000000000000000000010011010001",
			307 => "11111111110000110000010011010001",
			308 => "0000000000000000001101000100001100",
			309 => "0000001001000000001100100000001000",
			310 => "0000000011000000001111001000000100",
			311 => "11111110100011010000010100010101",
			312 => "00000001110111010000010100010101",
			313 => "11111110011000110000010100010101",
			314 => "0000000010000000000010000000001100",
			315 => "0000000100000000000000100100000100",
			316 => "00000010111110100000010100010101",
			317 => "0000000000000000000111100000000100",
			318 => "00000001000110110000010100010101",
			319 => "00000001111000100000010100010101",
			320 => "0000000110000000001100011000000100",
			321 => "00000011011000110000010100010101",
			322 => "0000001101000000001000011000000100",
			323 => "00000001000001110000010100010101",
			324 => "11111110010101010000010100010101",
			325 => "0000000000000000001100100100001100",
			326 => "0000001001000000001100100000001000",
			327 => "0000000011000000000111000000000100",
			328 => "11111110011100000000010101011001",
			329 => "00000011011100100000010101011001",
			330 => "11111110010111100000010101011001",
			331 => "0000000010000000000110010000010000",
			332 => "0000001110000000001011010100001100",
			333 => "0000000011000000000010111100000100",
			334 => "00000010100100100000010101011001",
			335 => "0000001111000000000001111100000100",
			336 => "00000001101000000000010101011001",
			337 => "11111110101110100000010101011001",
			338 => "00000011100100000000010101011001",
			339 => "0000000110000000001010011000000100",
			340 => "00000001101100110000010101011001",
			341 => "11111110010011010000010101011001",
			342 => "0000000000000000000010110100001000",
			343 => "0000001001000000001100100000000100",
			344 => "00000000000000000000010110011101",
			345 => "11111110011100110000010110011101",
			346 => "0000001100000000000100001000001100",
			347 => "0000000010000000001110110100001000",
			348 => "0000000000000000000110100000000100",
			349 => "00000000000000000000010110011101",
			350 => "00000001111001000000010110011101",
			351 => "00000000000000000000010110011101",
			352 => "0000000010000000000011001000000100",
			353 => "00000000110101010000010110011101",
			354 => "0000000110000000001100011000000100",
			355 => "00000000000000000000010110011101",
			356 => "0000001101000000001000011000000100",
			357 => "00000000000000000000010110011101",
			358 => "11111111010011110000010110011101",
			359 => "0000000000000000001101000100001100",
			360 => "0000001001000000001100100000001000",
			361 => "0000000011000000001111001000000100",
			362 => "11111110100111110000010111101001",
			363 => "00000001011110010000010111101001",
			364 => "11111110011001000000010111101001",
			365 => "0000000010000000000010000000010000",
			366 => "0000000100000000000000100100000100",
			367 => "00000010101110000000010111101001",
			368 => "0000001111000000000000001100000100",
			369 => "00000001110010010000010111101001",
			370 => "0000000000000000000111100000000100",
			371 => "00000000000000000000010111101001",
			372 => "00000001010110110000010111101001",
			373 => "0000000110000000001100011000000100",
			374 => "00000010111010100000010111101001",
			375 => "0000001101000000001000011000000100",
			376 => "00000000101110110000010111101001",
			377 => "11111110010111110000010111101001",
			378 => "0000001001000000001100100000011000",
			379 => "0000000101000000001110110000000100",
			380 => "11111111010101010000011000100101",
			381 => "0000000010000000001100010100000100",
			382 => "00000001100100010000011000100101",
			383 => "0000001101000000000100000100001000",
			384 => "0000000001000000001110011100000100",
			385 => "00000000000000000000011000100101",
			386 => "11111111011000100000011000100101",
			387 => "0000001101000000000000011100000100",
			388 => "00000000101001000000011000100101",
			389 => "00000000000000000000011000100101",
			390 => "0000001010000000000010111100000100",
			391 => "11111110011010110000011000100101",
			392 => "00000000000000000000011000100101",
			393 => "0000001001000000001100100000011000",
			394 => "0000000111000000000111001000010100",
			395 => "0000000101000000001110110000000100",
			396 => "00000000000000000000011001100001",
			397 => "0000001111000000000111001000001100",
			398 => "0000000001000000001110011100001000",
			399 => "0000000010000000001001100000000100",
			400 => "00000001000010010000011001100001",
			401 => "00000000000000000000011001100001",
			402 => "00000000000000000000011001100001",
			403 => "00000000000000000000011001100001",
			404 => "00000000000000000000011001100001",
			405 => "0000001010000000000010111100000100",
			406 => "11111110100011110000011001100001",
			407 => "00000000000000000000011001100001",
			408 => "0000001001000000001100100000011100",
			409 => "0000000101000000000100011000000100",
			410 => "11111110111101100000011010100101",
			411 => "0000001111000000000000001100000100",
			412 => "00000001101000010000011010100101",
			413 => "0000000110000000001100011000001000",
			414 => "0000000000000000000111100000000100",
			415 => "00000000000000000000011010100101",
			416 => "00000001101010010000011010100101",
			417 => "0000000111000000000001111100000100",
			418 => "00000001001011110000011010100101",
			419 => "0000001010000000000010111100000100",
			420 => "11111110100111110000011010100101",
			421 => "00000000000000000000011010100101",
			422 => "0000001010000000000010111100000100",
			423 => "11111110011010010000011010100101",
			424 => "00000000000000000000011010100101",
			425 => "0000000000000000001110101000001100",
			426 => "0000001001000000001100100000001000",
			427 => "0000000000000000000101100100000100",
			428 => "11111110011110000000011011111001",
			429 => "00000001110011100000011011111001",
			430 => "11111110011000000000011011111001",
			431 => "0000001001000000001100100000011000",
			432 => "0000001101000000000100000100010100",
			433 => "0000000011000000000010111100001000",
			434 => "0000001111000000000100001000000100",
			435 => "00000010001011110000011011111001",
			436 => "00000001010010100000011011111001",
			437 => "0000000110000000001010011000000100",
			438 => "00000010110111010000011011111001",
			439 => "0000000010000000000110010000000100",
			440 => "00000000011000100000011011111001",
			441 => "11111110010100010000011011111001",
			442 => "00000100100101010000011011111001",
			443 => "0000000010000000000010000000000100",
			444 => "00000001010010100000011011111001",
			445 => "11111110011000000000011011111001",
			446 => "0000001001000000001100100000100100",
			447 => "0000000000000000000110100000010000",
			448 => "0000001110000000001011010100001000",
			449 => "0000001001000000001100100000000100",
			450 => "00000000000000000000011101001101",
			451 => "11111111110000110000011101001101",
			452 => "0000000110000000000100110100000100",
			453 => "00000000100000110000011101001101",
			454 => "00000000000000000000011101001101",
			455 => "0000000110000000001101111100000100",
			456 => "00000011101011100000011101001101",
			457 => "0000001100000000001010111100001100",
			458 => "0000000000000000001101000100000100",
			459 => "00000000000000000000011101001101",
			460 => "0000001111000000001010111000000100",
			461 => "00000001010111100000011101001101",
			462 => "00000000000000000000011101001101",
			463 => "00000000000000000000011101001101",
			464 => "0000001010000000000010111100000100",
			465 => "11111110011100010000011101001101",
			466 => "00000000000000000000011101001101",
			467 => "0000000000000000001110101000010100",
			468 => "0000000001000000001110011100010000",
			469 => "0000001110000000001011010100001000",
			470 => "0000000000000000001001010100000100",
			471 => "11111110011110100000011110101001",
			472 => "11111111111001010000011110101001",
			473 => "0000001010000000001000110000000100",
			474 => "00000010101101110000011110101001",
			475 => "11111111101100000000011110101001",
			476 => "11111110011000100000011110101001",
			477 => "0000000010000000001110110100011000",
			478 => "0000001110000000000110001000010100",
			479 => "0000000011000000000010111100001000",
			480 => "0000001111000000000100001000000100",
			481 => "00000001111101100000011110101001",
			482 => "00000000110110000000011110101001",
			483 => "0000000000000000000101001000001000",
			484 => "0000000001000000001110011100000100",
			485 => "11111110100001000000011110101001",
			486 => "00000000000000000000011110101001",
			487 => "00000000111000100000011110101001",
			488 => "00000011011101110000011110101001",
			489 => "11111110100011000000011110101001",
			490 => "0000001001000000001100100000101100",
			491 => "0000000001000000001110011100100000",
			492 => "0000000000000000001101000100010000",
			493 => "0000001110000000001011010100001000",
			494 => "0000001001000000001100100000000100",
			495 => "00000000000000000000100000001101",
			496 => "11111111101010110000100000001101",
			497 => "0000000110000000000100110100000100",
			498 => "00000000101010000000100000001101",
			499 => "00000000000000000000100000001101",
			500 => "0000001100000000001101010100001100",
			501 => "0000000001000000001110011100001000",
			502 => "0000000010000000001110110100000100",
			503 => "00000001011110000000100000001101",
			504 => "00000000000000000000100000001101",
			505 => "00000000000000000000100000001101",
			506 => "00000000000000000000100000001101",
			507 => "0000000101000000001010001100000100",
			508 => "00000000000000000000100000001101",
			509 => "0000001000000000000110000100000100",
			510 => "00000100111110010000100000001101",
			511 => "00000000000000000000100000001101",
			512 => "0000001000000000001101111000000100",
			513 => "11111110011011110000100000001101",
			514 => "00000000000000000000100000001101",
			515 => "0000000000000000000101100100000100",
			516 => "11111110100010110000100001001011",
			517 => "0000000111000000000111001000011000",
			518 => "0000001001000000001100100000010100",
			519 => "0000001111000000000111001000010000",
			520 => "0000000001000000001110011100001100",
			521 => "0000000010000000001001100000001000",
			522 => "0000001100000000001100110000000100",
			523 => "00000000000000000000100001001011",
			524 => "00000001000111000000100001001011",
			525 => "00000000000000000000100001001011",
			526 => "00000000000000000000100001001011",
			527 => "00000000000000000000100001001011",
			528 => "00000000000000000000100001001011",
			529 => "00000000000000000000100001001011",
			530 => "00000000000000000000100001001101",
			531 => "00000000000000000000100001010001",
			532 => "00000000000000000000100001010101",
			533 => "00000000000000000000100001011001",
			534 => "00000000000000000000100001011101",
			535 => "00000000000000000000100001100001",
			536 => "00000000000000000000100001100101",
			537 => "00000000000000000000100001101001",
			538 => "00000000000000000000100001101101",
			539 => "00000000000000000000100001110001",
			540 => "00000000000000000000100001110101",
			541 => "00000000000000000000100001111001",
			542 => "00000000000000000000100001111101",
			543 => "00000000000000000000100010000001",
			544 => "00000000000000000000100010000101",
			545 => "00000000000000000000100010001001",
			546 => "00000000000000000000100010001101",
			547 => "00000000000000000000100010010001",
			548 => "00000000000000000000100010010101",
			549 => "00000000000000000000100010011001",
			550 => "00000000000000000000100010011101",
			551 => "00000000000000000000100010100001",
			552 => "00000000000000000000100010100101",
			553 => "00000000000000000000100010101001",
			554 => "00000000000000000000100010101101",
			555 => "00000000000000000000100010110001",
			556 => "00000000000000000000100010110101",
			557 => "00000000000000000000100010111001",
			558 => "00000000000000000000100010111101",
			559 => "00000000000000000000100011000001",
			560 => "00000000000000000000100011000101",
			561 => "00000000000000000000100011001001",
			562 => "00000000000000000000100011001101",
			563 => "00000000000000000000100011010001",
			564 => "00000000000000000000100011010101",
			565 => "00000000000000000000100011011001",
			566 => "00000000000000000000100011011101",
			567 => "0000001111000000001010111000000100",
			568 => "00000000000000000000100011101001",
			569 => "11111111111010100000100011101001",
			570 => "0000001111000000000000001100000100",
			571 => "00000000000000000000100011110101",
			572 => "11111111111101000000100011110101",
			573 => "0000000000000000001100100100000100",
			574 => "11111111111010100000100100000001",
			575 => "00000000000000000000100100000001",
			576 => "0000000000000000001100100100000100",
			577 => "11111111111011110000100100001101",
			578 => "00000000000000000000100100001101",
			579 => "0000001111000000000000001100000100",
			580 => "00000000000000000000100100011001",
			581 => "11111111111010010000100100011001",
			582 => "0000000000000000000110100000001000",
			583 => "0000001111000000000000001100000100",
			584 => "00000000000000000000100100101101",
			585 => "11111111111000100000100100101101",
			586 => "00000000000000000000100100101101",
			587 => "0000000000000000000110100000001000",
			588 => "0000001111000000001100101100000100",
			589 => "00000000000000000000100101001001",
			590 => "11111111101000000000100101001001",
			591 => "0000001110000000001001101000000100",
			592 => "00000000000000000000100101001001",
			593 => "00000000000100110000100101001001",
			594 => "0000000001000000001110011100001100",
			595 => "0000000010000000001001100000001000",
			596 => "0000000101000000001110110000000100",
			597 => "00000000000000000000100101100101",
			598 => "00000000011110100000100101100101",
			599 => "00000000000000000000100101100101",
			600 => "11111111000101100000100101100101",
			601 => "0000000000000000000111100000001100",
			602 => "0000001111000000001110001100000100",
			603 => "00000000000000000000100110000001",
			604 => "0000001010000000000010111100000100",
			605 => "11111111100010100000100110000001",
			606 => "00000000000000000000100110000001",
			607 => "00000000000000000000100110000001",
			608 => "0000000001000000001110011100001100",
			609 => "0000001110000000001100011100000100",
			610 => "00000000000000000000100110011101",
			611 => "0000001111000000001010111000000100",
			612 => "00000000000010110000100110011101",
			613 => "00000000000000000000100110011101",
			614 => "00000000000000000000100110011101",
			615 => "0000001111000000001010111000001100",
			616 => "0000001100000000001101010100001000",
			617 => "0000001100000000001100110000000100",
			618 => "00000000000000000000100110111001",
			619 => "00000000001001010000100110111001",
			620 => "00000000000000000000100110111001",
			621 => "00000000000000000000100110111001",
			622 => "0000001001000000001100100000001100",
			623 => "0000001111000000001010111000001000",
			624 => "0000001000000000001011000100000100",
			625 => "00000000000000000000100111010101",
			626 => "00000000000001100000100111010101",
			627 => "00000000000000000000100111010101",
			628 => "00000000000000000000100111010101",
			629 => "0000001111000000001010111000001100",
			630 => "0000000111000000000110000100000100",
			631 => "00000000000000000000100111110001",
			632 => "0000000001000000001110011100000100",
			633 => "00000000000100100000100111110001",
			634 => "00000000000000000000100111110001",
			635 => "00000000000000000000100111110001",
			636 => "0000000000000000000110100000001000",
			637 => "0000001001000000001100100000000100",
			638 => "00000000000000000000101000010101",
			639 => "11111110110011000000101000010101",
			640 => "0000001100000000000100001000001000",
			641 => "0000000010000000001110110100000100",
			642 => "00000000110000010000101000010101",
			643 => "00000000000000000000101000010101",
			644 => "00000000000000000000101000010101",
			645 => "0000001111000000001010111000010000",
			646 => "0000000110000000001100011000001100",
			647 => "0000000111000000000110000100000100",
			648 => "00000000000000000000101000111001",
			649 => "0000001001000000001100100000000100",
			650 => "00000000100100100000101000111001",
			651 => "00000000000000000000101000111001",
			652 => "00000000000000000000101000111001",
			653 => "11111110111110010000101000111001",
			654 => "0000000000000000000101100100000100",
			655 => "11111111001110110000101001011101",
			656 => "0000000110000000001100011000001100",
			657 => "0000001001000000001100100000001000",
			658 => "0000000111000000001101111000000100",
			659 => "00000000000000000000101001011101",
			660 => "00000000100000010000101001011101",
			661 => "00000000000000000000101001011101",
			662 => "00000000000000000000101001011101",
			663 => "0000000001000000001110011100010000",
			664 => "0000001100000000000001111100001100",
			665 => "0000000111000000000110000100000100",
			666 => "00000000000000000000101010000001",
			667 => "0000001111000000001010111000000100",
			668 => "00000000001101110000101010000001",
			669 => "00000000000000000000101010000001",
			670 => "00000000000000000000101010000001",
			671 => "11111111101100000000101010000001",
			672 => "0000001111000000001010111000010000",
			673 => "0000001100000000000100001000001100",
			674 => "0000000111000000000111001000001000",
			675 => "0000001100000000001100110000000100",
			676 => "00000000000000000000101010100101",
			677 => "00000000001001000000101010100101",
			678 => "00000000000000000000101010100101",
			679 => "00000000000000000000101010100101",
			680 => "11111111101111100000101010100101",
			681 => "0000001111000000000111001000010000",
			682 => "0000001110000000001001101000000100",
			683 => "00000000000000000000101011001001",
			684 => "0000001100000000001101010100001000",
			685 => "0000000111000000001110001100000100",
			686 => "00000000000000000000101011001001",
			687 => "00000000000110000000101011001001",
			688 => "00000000000000000000101011001001",
			689 => "11111111110110110000101011001001",
			690 => "0000001001000000001100100000010000",
			691 => "0000001100000000001110001100000100",
			692 => "00000000000000000000101011101101",
			693 => "0000001100000000001101010100001000",
			694 => "0000001111000000000111001000000100",
			695 => "00000000001000110000101011101101",
			696 => "00000000000000000000101011101101",
			697 => "00000000000000000000101011101101",
			698 => "00000000000000000000101011101101",
			699 => "0000000000000000000110100000001000",
			700 => "0000001111000000001100101100000100",
			701 => "00000000000000000000101100011001",
			702 => "11111111100100100000101100011001",
			703 => "0000001110000000001001101000000100",
			704 => "00000000000000000000101100011001",
			705 => "0000001100000000001101010100001000",
			706 => "0000001100000000000000001100000100",
			707 => "00000000000000000000101100011001",
			708 => "00000000000111110000101100011001",
			709 => "00000000000000000000101100011001",
			710 => "0000001001000000001100100000010100",
			711 => "0000000010000000001010001000001000",
			712 => "0000000101000000001110110000000100",
			713 => "00000000000000000000101101000101",
			714 => "00000000111011100000101101000101",
			715 => "0000000111000000000001111100000100",
			716 => "00000000000001100000101101000101",
			717 => "0000001101000000000100000100000100",
			718 => "11111111111010000000101101000101",
			719 => "00000000000000000000101101000101",
			720 => "11111110101011000000101101000101",
			721 => "0000000001000000001110011100010000",
			722 => "0000000101000000001110110000000100",
			723 => "11111111101100010000101101111001",
			724 => "0000001111000000001010111100001000",
			725 => "0000001100000000001101010100000100",
			726 => "00000001011111000000101101111001",
			727 => "00000000000000000000101101111001",
			728 => "00000000000000000000101101111001",
			729 => "0000001010000000000010011000000100",
			730 => "11111110011011000000101101111001",
			731 => "0000001111000000000100001000000100",
			732 => "00000000010101110000101101111001",
			733 => "00000000000000000000101101111001",
			734 => "0000000000000000000010110100001000",
			735 => "0000001001000000001100100000000100",
			736 => "00000000000000000000101110101101",
			737 => "11111110011001110000101110101101",
			738 => "0000001111000000000000001100000100",
			739 => "00000001100111000000101110101101",
			740 => "0000000110000000001100011000001000",
			741 => "0000000010000000000010000100000100",
			742 => "00000001101111000000101110101101",
			743 => "00000000000000000000101110101101",
			744 => "0000001010000000000010111100000100",
			745 => "11111110100001100000101110101101",
			746 => "00000001010000110000101110101101",
			747 => "0000000000000000000110100000001000",
			748 => "0000001001000000001100100000000100",
			749 => "00000000000000000000101111100001",
			750 => "11111110011110000000101111100001",
			751 => "0000000010000000000011001000000100",
			752 => "00000001101110100000101111100001",
			753 => "0000000111000000001101010100001000",
			754 => "0000000111000000001010111100000100",
			755 => "00000000001111010000101111100001",
			756 => "00000000000000000000101111100001",
			757 => "0000000110000000001100011000000100",
			758 => "00000000000000000000101111100001",
			759 => "11111111011101110000101111100001",
			760 => "0000000001000000001110011100011000",
			761 => "0000000110000000001100011000001100",
			762 => "0000000101000000000100011000000100",
			763 => "00000000000000000000110000011101",
			764 => "0000001001000000001100100000000100",
			765 => "00000001100100000000110000011101",
			766 => "00000000000000000000110000011101",
			767 => "0000001010000000000010111100001000",
			768 => "0000000010000000001010001000000100",
			769 => "00000000000000000000110000011101",
			770 => "11111111011001010000110000011101",
			771 => "00000000101010000000110000011101",
			772 => "0000001010000000000010111100000100",
			773 => "11111110011111110000110000011101",
			774 => "00000000000000000000110000011101",
			775 => "0000001001000000001100100000010100",
			776 => "0000000111000000000111001000010000",
			777 => "0000000101000000001110110000000100",
			778 => "00000000000000000000110001010001",
			779 => "0000001111000000000111001000001000",
			780 => "0000000001000000001110011100000100",
			781 => "00000001001010010000110001010001",
			782 => "00000000000000000000110001010001",
			783 => "00000000000000000000110001010001",
			784 => "00000000000000000000110001010001",
			785 => "0000001010000000000010111100000100",
			786 => "11111110100010000000110001010001",
			787 => "00000000000000000000110001010001",
			788 => "0000001000000000000101101100001000",
			789 => "0000001001000000001100100000000100",
			790 => "00000000000000000000110010000101",
			791 => "11111111011010100000110010000101",
			792 => "0000000111000000000111001000010000",
			793 => "0000001001000000001100100000000100",
			794 => "00000000000000000000110010000101",
			795 => "0000001111000000000111001000001000",
			796 => "0000001001000000001100100000000100",
			797 => "00000000001110010000110010000101",
			798 => "00000000000000000000110010000101",
			799 => "00000000000000000000110010000101",
			800 => "00000000000000000000110010000101",
			801 => "0000001100000000001110001100001000",
			802 => "0000001000000000001110001100000100",
			803 => "11111111101111110000110010111001",
			804 => "00000000000000000000110010111001",
			805 => "0000000111000000000111001000010000",
			806 => "0000001001000000001100100000001100",
			807 => "0000001100000000000100001000001000",
			808 => "0000001111000000000111001000000100",
			809 => "00000000001010110000110010111001",
			810 => "00000000000000000000110010111001",
			811 => "00000000000000000000110010111001",
			812 => "00000000000000000000110010111001",
			813 => "00000000000000000000110010111001",
			814 => "0000000000000000000101100100000100",
			815 => "11111111010011110000110011100101",
			816 => "0000000111000000000111001000010000",
			817 => "0000001001000000001100100000001100",
			818 => "0000000001000000001110011100001000",
			819 => "0000001100000000001100110000000100",
			820 => "00000000000000000000110011100101",
			821 => "00000000011100100000110011100101",
			822 => "00000000000000000000110011100101",
			823 => "00000000000000000000110011100101",
			824 => "00000000000000000000110011100101",
			825 => "0000001111000000001010111000010100",
			826 => "0000001001000000001100100000010000",
			827 => "0000001100000000001101010100001100",
			828 => "0000000101000000000100011000000100",
			829 => "00000000000000000000110100010001",
			830 => "0000000001000000001110011100000100",
			831 => "00000000000110110000110100010001",
			832 => "00000000000000000000110100010001",
			833 => "00000000000000000000110100010001",
			834 => "00000000000000000000110100010001",
			835 => "00000000000000000000110100010001",
			836 => "0000000000000000000101100100000100",
			837 => "11111110011011110000110101000101",
			838 => "0000000001000000001110011100010000",
			839 => "0000001100000000001101010100001100",
			840 => "0000001111000000000111001000001000",
			841 => "0000000010000000001001100000000100",
			842 => "00000001010110000000110101000101",
			843 => "00000000000000000000110101000101",
			844 => "00000000000000000000110101000101",
			845 => "00000000000000000000110101000101",
			846 => "0000001111000000000000001100000100",
			847 => "00000000000100010000110101000101",
			848 => "11111111011001010000110101000101",
			849 => "0000000000000000001100100100001100",
			850 => "0000001001000000001100100000001000",
			851 => "0000000011000000000111000000000100",
			852 => "11111110011101010000110110001001",
			853 => "00000010110001000000110110001001",
			854 => "11111110010111110000110110001001",
			855 => "0000000010000000000110010000010000",
			856 => "0000001110000000001011010100001100",
			857 => "0000000011000000000010111100000100",
			858 => "00000010010110000000110110001001",
			859 => "0000001111000000000001111100000100",
			860 => "00000001011001110000110110001001",
			861 => "11111110110010010000110110001001",
			862 => "00000011010000010000110110001001",
			863 => "0000000111000000001101010100000100",
			864 => "00000001011101110000110110001001",
			865 => "11111110010100100000110110001001",
			866 => "0000000000000000000010110100001000",
			867 => "0000000001000000001110011100000100",
			868 => "00000000000000000000110111001101",
			869 => "11111110011101100000110111001101",
			870 => "0000001100000000000100001000001100",
			871 => "0000000010000000001110110100001000",
			872 => "0000000000000000000110100000000100",
			873 => "00000000000000000000110111001101",
			874 => "00000001110001010000110111001101",
			875 => "00000000000000000000110111001101",
			876 => "0000000010000000000011001000000100",
			877 => "00000000101100110000110111001101",
			878 => "0000000110000000001100011000000100",
			879 => "00000000000000000000110111001101",
			880 => "0000001101000000001000011000000100",
			881 => "00000000000000000000110111001101",
			882 => "11111111011110010000110111001101",
			883 => "0000001001000000001100100000011000",
			884 => "0000000101000000000100011000000100",
			885 => "11111111001001010000111000001001",
			886 => "0000001111000000000000001100000100",
			887 => "00000001100110010000111000001001",
			888 => "0000000110000000001100011000001000",
			889 => "0000000000000000000111100000000100",
			890 => "00000000000000000000111000001001",
			891 => "00000001011111010000111000001001",
			892 => "0000000111000000000001111100000100",
			893 => "00000001000000110000111000001001",
			894 => "11111110110101010000111000001001",
			895 => "0000001010000000000010111100000100",
			896 => "11111110011010100000111000001001",
			897 => "00000000000000000000111000001001",
			898 => "0000000000000000001101000100011000",
			899 => "0000001001000000001100100000010100",
			900 => "0000000110000000000111101000001000",
			901 => "0000001111000000001001110000000100",
			902 => "00000000000000000000111001010101",
			903 => "00000010010111010000111001010101",
			904 => "0000000001000000001110011100001000",
			905 => "0000001001000000001100100000000100",
			906 => "00000000001101010000111001010101",
			907 => "00000000000000000000111001010101",
			908 => "11111110100100110000111001010101",
			909 => "11111110011001010000111001010101",
			910 => "0000000010000000001100010100000100",
			911 => "00000001101011100000111001010101",
			912 => "0000000110000000001100011000000100",
			913 => "00000010010000100000111001010101",
			914 => "0000000100000000000011100100000100",
			915 => "11111110011100100000111001010101",
			916 => "00000000000000000000111001010101",
			917 => "0000000000000000000101100100000100",
			918 => "11111110101100100000111010011001",
			919 => "0000000110000000001100011000001100",
			920 => "0000001001000000001100100000001000",
			921 => "0000000111000000001101111000000100",
			922 => "00000000000000000000111010011001",
			923 => "00000001000000000000111010011001",
			924 => "00000000000000000000111010011001",
			925 => "0000000111000000000001111100001000",
			926 => "0000000011000000000010011000000100",
			927 => "00000000010010000000111010011001",
			928 => "00000000000000000000111010011001",
			929 => "0000000110000000001101011000001000",
			930 => "0000000011000000001111000100000100",
			931 => "00000000000000000000111010011001",
			932 => "11111111111000100000111010011001",
			933 => "00000000000000000000111010011001",
			934 => "0000001001000000001100100000011100",
			935 => "0000000101000000000100011000000100",
			936 => "11111111000011000000111011011101",
			937 => "0000001111000000000000001100000100",
			938 => "00000001100111010000111011011101",
			939 => "0000000110000000001100011000001000",
			940 => "0000000000000000000111100000000100",
			941 => "00000000000000000000111011011101",
			942 => "00000001100100100000111011011101",
			943 => "0000000111000000000001111100000100",
			944 => "00000001000110110000111011011101",
			945 => "0000001010000000000010111100000100",
			946 => "11111110101011010000111011011101",
			947 => "00000000000000000000111011011101",
			948 => "0000001010000000000010111100000100",
			949 => "11111110011010010000111011011101",
			950 => "00000000000000000000111011011101",
			951 => "0000000000000000001110101000010100",
			952 => "0000000001000000001110011100010000",
			953 => "0000001110000000001011010100001000",
			954 => "0000000000000000001001010100000100",
			955 => "11111110011101100000111100110001",
			956 => "11111111110110110000111100110001",
			957 => "0000001010000000001000110000000100",
			958 => "00000011000101000000111100110001",
			959 => "11111111100101110000111100110001",
			960 => "11111110011000010000111100110001",
			961 => "0000000010000000001110110100010100",
			962 => "0000001110000000000110001000010000",
			963 => "0000000010000000001100010100000100",
			964 => "00000010000011100000111100110001",
			965 => "0000000110000000001010011000000100",
			966 => "00000010101101110000111100110001",
			967 => "0000001011000000000111001000000100",
			968 => "00000001000000100000111100110001",
			969 => "11111110001111110000111100110001",
			970 => "00000011101110010000111100110001",
			971 => "11111110100001000000111100110001",
			972 => "0000000000000000001100100100010100",
			973 => "0000001001000000001100100000001000",
			974 => "0000000000000000001001010100000100",
			975 => "11111110011001000000111110001101",
			976 => "00001011000010100000111110001101",
			977 => "0000001010000000000010011000000100",
			978 => "11111110010110100000111110001101",
			979 => "0000001000000000001100110000000100",
			980 => "11111110100101010000111110001101",
			981 => "00000010010100110000111110001101",
			982 => "0000000010000000001110110100011000",
			983 => "0000001111000000000111001000010100",
			984 => "0000001100000000001010111100001100",
			985 => "0000001111000000000001111100001000",
			986 => "0000001111000000000100001000000100",
			987 => "00000100001001110000111110001101",
			988 => "00000010101111000000111110001101",
			989 => "00001001111000100000111110001101",
			990 => "0000000010000000001100010100000100",
			991 => "00000011111110100000111110001101",
			992 => "11111110011011010000111110001101",
			993 => "00001001101000010000111110001101",
			994 => "11111110011011110000111110001101",
			995 => "0000000000000000001101000100001100",
			996 => "0000001001000000001100100000001000",
			997 => "0000000011000000001111001000000100",
			998 => "11111110100101010000111111100001",
			999 => "00000001101001110000111111100001",
			1000 => "11111110011000110000111111100001",
			1001 => "0000000010000000001001100000011100",
			1002 => "0000001100000000001010111100010100",
			1003 => "0000001001000000001100100000010000",
			1004 => "0000001111000000000001111100001000",
			1005 => "0000000010000000001100010100000100",
			1006 => "00000001110101010000111111100001",
			1007 => "00000000000111100000111111100001",
			1008 => "0000001000000000001110001100000100",
			1009 => "00000110011111000000111111100001",
			1010 => "00000010011100100000111111100001",
			1011 => "11111110110010100000111111100001",
			1012 => "0000000010000000001100010100000100",
			1013 => "00000001100001000000111111100001",
			1014 => "11111110011001000000111111100001",
			1015 => "11111110100001100000111111100001",
			1016 => "0000000000000000000101001000101100",
			1017 => "0000000000000000001100100100011100",
			1018 => "0000001001000000001100100000001000",
			1019 => "0000001010000000000111000100000100",
			1020 => "11001001110001010001000001000101",
			1021 => "11011101000101100001000001000101",
			1022 => "0000001001000000001100100000001000",
			1023 => "0000001010000000000111000100000100",
			1024 => "11001001101110000001000001000101",
			1025 => "11010101001111000001000001000101",
			1026 => "0000001010000000000010011000000100",
			1027 => "11001001101001100001000001000101",
			1028 => "0000001010000000000010111100000100",
			1029 => "11001100011010100001000001000101",
			1030 => "11001001111000010001000001000101",
			1031 => "0000000010000000001100010100000100",
			1032 => "11110100100001000001000001000101",
			1033 => "0000001100000000000100001000000100",
			1034 => "11010111001010010001000001000101",
			1035 => "0000000010000000000010000000000100",
			1036 => "11001101011000100001000001000101",
			1037 => "11001001101110000001000001000101",
			1038 => "0000001111000000001010111100000100",
			1039 => "11110110001110110001000001000101",
			1040 => "11010101001111000001000001000101",
			1041 => "0000000000000000001101000100001100",
			1042 => "0000001001000000001100100000001000",
			1043 => "0000000011000000001011010100000100",
			1044 => "11111110101011000001000010011011",
			1045 => "00000001011110100001000010011011",
			1046 => "11111110011001000001000010011011",
			1047 => "0000001111000000000111001000011100",
			1048 => "0000001001000000001100100000011000",
			1049 => "0000000000000000001101000100000100",
			1050 => "00000100110100000001000010011011",
			1051 => "0000000000000000000111100000001000",
			1052 => "0000000010000000001100010100000100",
			1053 => "00000001110110100001000010011011",
			1054 => "11111110100110010001000010011011",
			1055 => "0000001101000000000100000100001000",
			1056 => "0000001101000000001010011100000100",
			1057 => "00000001110010000001000010011011",
			1058 => "00000001000011000001000010011011",
			1059 => "00000010110100000001000010011011",
			1060 => "11111111011001110001000010011011",
			1061 => "11111110100110100001000010011011",
			1062 => "00000000000000000001000010011101",
			1063 => "00000000000000000001000010100001",
			1064 => "00000000000000000001000010100101",
			1065 => "00000000000000000001000010101001",
			1066 => "00000000000000000001000010101101",
			1067 => "00000000000000000001000010110001",
			1068 => "00000000000000000001000010110101",
			1069 => "00000000000000000001000010111001",
			1070 => "00000000000000000001000010111101",
			1071 => "00000000000000000001000011000001",
			1072 => "00000000000000000001000011000101",
			1073 => "00000000000000000001000011001001",
			1074 => "00000000000000000001000011001101",
			1075 => "00000000000000000001000011010001",
			1076 => "00000000000000000001000011010101",
			1077 => "00000000000000000001000011011001",
			1078 => "00000000000000000001000011011101",
			1079 => "00000000000000000001000011100001",
			1080 => "00000000000000000001000011100101",
			1081 => "00000000000000000001000011101001",
			1082 => "00000000000000000001000011101101",
			1083 => "00000000000000000001000011110001",
			1084 => "00000000000000000001000011110101",
			1085 => "00000000000000000001000011111001",
			1086 => "00000000000000000001000011111101",
			1087 => "00000000000000000001000100000001",
			1088 => "00000000000000000001000100000101",
			1089 => "00000000000000000001000100001001",
			1090 => "00000000000000000001000100001101",
			1091 => "00000000000000000001000100010001",
			1092 => "00000000000000000001000100010101",
			1093 => "00000000000000000001000100011001",
			1094 => "00000000000000000001000100011101",
			1095 => "00000000000000000001000100100001",
			1096 => "00000000000000000001000100100101",
			1097 => "00000000000000000001000100101001",
			1098 => "00000000000000000001000100101101",
			1099 => "0000001111000000001010111000000100",
			1100 => "00000000000000000001000100111001",
			1101 => "11111111111011000001000100111001",
			1102 => "0000001111000000000000001100000100",
			1103 => "00000000000000000001000101000101",
			1104 => "11111111111111110001000101000101",
			1105 => "0000000000000000001100100100000100",
			1106 => "11111111111011010001000101010001",
			1107 => "00000000000000000001000101010001",
			1108 => "0000001111000000000000001100000100",
			1109 => "00000000000000000001000101011101",
			1110 => "11111111111011000001000101011101",
			1111 => "0000000000000000001001010100000100",
			1112 => "11111110111100100001000101110001",
			1113 => "0000000010000000001010001000000100",
			1114 => "00000000011011110001000101110001",
			1115 => "00000000000000000001000101110001",
			1116 => "0000001111000000000000001100000100",
			1117 => "00000000000000000001000110000101",
			1118 => "0000001001000000001100100000000100",
			1119 => "00000000000000000001000110000101",
			1120 => "11111111110110000001000110000101",
			1121 => "0000000000000000000101100100000100",
			1122 => "11111110100111000001000110100001",
			1123 => "0000000010000000001110010000001000",
			1124 => "0000001001000000001100100000000100",
			1125 => "00000001000100010001000110100001",
			1126 => "00000000000000000001000110100001",
			1127 => "00000000000000000001000110100001",
			1128 => "0000000001000000001110011100001100",
			1129 => "0000000101000000001110110000000100",
			1130 => "00000000000000000001000110111101",
			1131 => "0000000110000000001100011000000100",
			1132 => "00000000100010000001000110111101",
			1133 => "00000000000000000001000110111101",
			1134 => "11111111001010010001000110111101",
			1135 => "0000000000000000000111100000001100",
			1136 => "0000001111000000001110001100000100",
			1137 => "00000000000000000001000111011001",
			1138 => "0000001010000000000010111100000100",
			1139 => "11111111100100100001000111011001",
			1140 => "00000000000000000001000111011001",
			1141 => "00000000000000000001000111011001",
			1142 => "0000000001000000001110011100001100",
			1143 => "0000000100000000000010100000000100",
			1144 => "00000000000000000001000111110101",
			1145 => "0000001111000000001010111000000100",
			1146 => "00000000000010010001000111110101",
			1147 => "00000000000000000001000111110101",
			1148 => "00000000000000000001000111110101",
			1149 => "0000001111000000001010111000001100",
			1150 => "0000001100000000001101010100001000",
			1151 => "0000001100000000001100110000000100",
			1152 => "00000000000000000001001000010001",
			1153 => "00000000001000100001001000010001",
			1154 => "00000000000000000001001000010001",
			1155 => "00000000000000000001001000010001",
			1156 => "0000001001000000001100100000001100",
			1157 => "0000001111000000001010111000001000",
			1158 => "0000000000000000000101100100000100",
			1159 => "00000000000000000001001000101101",
			1160 => "00000000000001100001001000101101",
			1161 => "00000000000000000001001000101101",
			1162 => "00000000000000000001001000101101",
			1163 => "0000001001000000001100100000001100",
			1164 => "0000000010000000001110010000001000",
			1165 => "0000000101000000000100011000000100",
			1166 => "00000000000000000001001001010001",
			1167 => "00000001001000010001001001010001",
			1168 => "00000000000000000001001001010001",
			1169 => "0000001010000000000010111100000100",
			1170 => "11111110100101110001001001010001",
			1171 => "00000000000000000001001001010001",
			1172 => "0000000000000000000110100000001000",
			1173 => "0000001111000000001100101100000100",
			1174 => "00000000000000000001001001110101",
			1175 => "11111110110101000001001001110101",
			1176 => "0000001100000000000100001000001000",
			1177 => "0000000010000000001110110100000100",
			1178 => "00000000101100000001001001110101",
			1179 => "00000000000000000001001001110101",
			1180 => "00000000000000000001001001110101",
			1181 => "0000001111000000001010111000010000",
			1182 => "0000000110000000001100011000001100",
			1183 => "0000001100000000001100110000000100",
			1184 => "00000000000000000001001010011001",
			1185 => "0000001001000000001100100000000100",
			1186 => "00000000100010010001001010011001",
			1187 => "00000000000000000001001010011001",
			1188 => "00000000000000000001001010011001",
			1189 => "11111111000000100001001010011001",
			1190 => "0000001111000000001010111000010000",
			1191 => "0000000111000000000111001000001100",
			1192 => "0000001100000000001100110000000100",
			1193 => "00000000000000000001001010111101",
			1194 => "0000001001000000001100100000000100",
			1195 => "00000000011010100001001010111101",
			1196 => "00000000000000000001001010111101",
			1197 => "00000000000000000001001010111101",
			1198 => "11111111010110010001001010111101",
			1199 => "0000000001000000001110011100010000",
			1200 => "0000001100000000000001111100001100",
			1201 => "0000000101000000001110110000000100",
			1202 => "00000000000000000001001011100001",
			1203 => "0000001111000000001010111000000100",
			1204 => "00000000001100100001001011100001",
			1205 => "00000000000000000001001011100001",
			1206 => "00000000000000000001001011100001",
			1207 => "11111111101101100001001011100001",
			1208 => "0000001111000000001010111000010000",
			1209 => "0000001110000000001001101000000100",
			1210 => "00000000000000000001001100000101",
			1211 => "0000001001000000001100100000001000",
			1212 => "0000001100000000001101010100000100",
			1213 => "00000000001000100001001100000101",
			1214 => "00000000000000000001001100000101",
			1215 => "00000000000000000001001100000101",
			1216 => "11111111110010000001001100000101",
			1217 => "0000001111000000000111001000010000",
			1218 => "0000001110000000001001101000000100",
			1219 => "00000000000000000001001100101001",
			1220 => "0000001100000000001101010100001000",
			1221 => "0000000111000000001110001100000100",
			1222 => "00000000000000000001001100101001",
			1223 => "00000000000101010001001100101001",
			1224 => "00000000000000000001001100101001",
			1225 => "11111111110111100001001100101001",
			1226 => "0000000000000000000110100000001000",
			1227 => "0000001001000000001100100000000100",
			1228 => "00000000000000000001001101010101",
			1229 => "11111110011111010001001101010101",
			1230 => "0000000010000000000011001000000100",
			1231 => "00000001100101010001001101010101",
			1232 => "0000000101000000000001101000000100",
			1233 => "00000000001000100001001101010101",
			1234 => "0000000011000000000011010000000100",
			1235 => "11111111101111010001001101010101",
			1236 => "00000000000000000001001101010101",
			1237 => "0000001100000000001110001100001000",
			1238 => "0000001000000000001110001100000100",
			1239 => "11111111110001000001001110000001",
			1240 => "00000000000000000001001110000001",
			1241 => "0000000111000000000111001000001100",
			1242 => "0000001001000000001100100000001000",
			1243 => "0000001100000000000100001000000100",
			1244 => "00000000001001100001001110000001",
			1245 => "00000000000000000001001110000001",
			1246 => "00000000000000000001001110000001",
			1247 => "00000000000000000001001110000001",
			1248 => "0000000100000000001101110000000100",
			1249 => "11111110111010010001001110101101",
			1250 => "0000000110000000001100011000001000",
			1251 => "0000001001000000001100100000000100",
			1252 => "00000000011111000001001110101101",
			1253 => "00000000000000000001001110101101",
			1254 => "0000000010000000001010001000000100",
			1255 => "00000000000000000001001110101101",
			1256 => "0000001111000000001101111000000100",
			1257 => "00000000000000000001001110101101",
			1258 => "11111111111000000001001110101101",
			1259 => "0000001001000000001100100000010100",
			1260 => "0000000110000000001100011000001000",
			1261 => "0000000000000000000001001000000100",
			1262 => "00000000000000000001001111100001",
			1263 => "00000000100001000001001111100001",
			1264 => "0000001111000000001101111000000100",
			1265 => "00000000000000000001001111100001",
			1266 => "0000000000000000000010011100000100",
			1267 => "11111111111000000001001111100001",
			1268 => "00000000000000000001001111100001",
			1269 => "0000001111000000000000001100000100",
			1270 => "00000000000000000001001111100001",
			1271 => "11111110110111100001001111100001",
			1272 => "0000000000000000000010110100001000",
			1273 => "0000001001000000001100100000000100",
			1274 => "00000000000000000001010000010101",
			1275 => "11111110011010000001010000010101",
			1276 => "0000001111000000000000001100000100",
			1277 => "00000001100110010001010000010101",
			1278 => "0000000110000000001100011000001000",
			1279 => "0000000010000000000010000100000100",
			1280 => "00000001101101000001010000010101",
			1281 => "00000000000000000001010000010101",
			1282 => "0000000111000000000001111100000100",
			1283 => "00000001010110000001010000010101",
			1284 => "11111110101000010001010000010101",
			1285 => "0000001000000000000101101100001000",
			1286 => "0000000001000000001110011100000100",
			1287 => "00000000000000000001010001001001",
			1288 => "11111110011110100001010001001001",
			1289 => "0000000010000000000011001000000100",
			1290 => "00000001101001100001010001001001",
			1291 => "0000000111000000001101010100001000",
			1292 => "0000001100000000000100001000000100",
			1293 => "00000000001011000001010001001001",
			1294 => "00000000000000000001010001001001",
			1295 => "0000000110000000001100011000000100",
			1296 => "00000000000000000001010001001001",
			1297 => "11111111011111000001010001001001",
			1298 => "0000000001000000001110011100011000",
			1299 => "0000000110000000001100011000001100",
			1300 => "0000000101000000000100011000000100",
			1301 => "00000000000000000001010010000101",
			1302 => "0000001001000000001100100000000100",
			1303 => "00000001011011110001010010000101",
			1304 => "00000000000000000001010010000101",
			1305 => "0000001010000000000010111100001000",
			1306 => "0000000010000000001010001000000100",
			1307 => "00000000000000000001010010000101",
			1308 => "11111111011111100001010010000101",
			1309 => "00000000100001000001010010000101",
			1310 => "0000001010000000000010111100000100",
			1311 => "11111110100001010001010010000101",
			1312 => "00000000000000000001010010000101",
			1313 => "0000001111000000001010111000011000",
			1314 => "0000000110000000001100011000001100",
			1315 => "0000000111000000001110001100000100",
			1316 => "00000000000000000001010010111001",
			1317 => "0000001001000000001100100000000100",
			1318 => "00000000111010000001010010111001",
			1319 => "00000000000000000001010010111001",
			1320 => "0000000111000000000001111100001000",
			1321 => "0000000101000000000001101000000100",
			1322 => "00000000001000010001010010111001",
			1323 => "00000000000000000001010010111001",
			1324 => "00000000000000000001010010111001",
			1325 => "11111110110000000001010010111001",
			1326 => "0000000000000000000110100000001000",
			1327 => "0000001111000000000000001100000100",
			1328 => "00000000000000000001010011101101",
			1329 => "11111111011010100001010011101101",
			1330 => "0000000001000000001110011100000100",
			1331 => "00000000000000000001010011101101",
			1332 => "0000001111000000000111001000001100",
			1333 => "0000001001000000001100100000001000",
			1334 => "0000000001000000001110011100000100",
			1335 => "00000000001110000001010011101101",
			1336 => "00000000000000000001010011101101",
			1337 => "00000000000000000001010011101101",
			1338 => "00000000000000000001010011101101",
			1339 => "0000000000000000000101100100000100",
			1340 => "11111110101110010001010100011001",
			1341 => "0000001100000000000100001000010000",
			1342 => "0000000010000000001110110100001100",
			1343 => "0000001001000000001100100000001000",
			1344 => "0000000111000000000111001000000100",
			1345 => "00000000110110100001010100011001",
			1346 => "00000000000000000001010100011001",
			1347 => "00000000000000000001010100011001",
			1348 => "00000000000000000001010100011001",
			1349 => "00000000000000000001010100011001",
			1350 => "0000001000000000000011011100000100",
			1351 => "11111111100000100001010101000101",
			1352 => "0000001110000000001001101000000100",
			1353 => "00000000000000000001010101000101",
			1354 => "0000001000000000001100110000000100",
			1355 => "00000000000000000001010101000101",
			1356 => "0000001100000000001101010100001000",
			1357 => "0000001111000000000111001000000100",
			1358 => "00000000010100100001010101000101",
			1359 => "00000000000000000001010101000101",
			1360 => "00000000000000000001010101000101",
			1361 => "0000001111000000001010111000010100",
			1362 => "0000001001000000001100100000010000",
			1363 => "0000001100000000001101010100001100",
			1364 => "0000000101000000000100011000000100",
			1365 => "00000000000000000001010101110001",
			1366 => "0000000001000000001110011100000100",
			1367 => "00000000000110000001010101110001",
			1368 => "00000000000000000001010101110001",
			1369 => "00000000000000000001010101110001",
			1370 => "00000000000000000001010101110001",
			1371 => "00000000000000000001010101110001",
			1372 => "0000001001000000001100100000011000",
			1373 => "0000000010000000001010001000001000",
			1374 => "0000000101000000001110110000000100",
			1375 => "00000000000000000001010110100101",
			1376 => "00000000111111010001010110100101",
			1377 => "0000001111000000000001111100000100",
			1378 => "00000000000000000001010110100101",
			1379 => "0000001111000000001010111000001000",
			1380 => "0000000111000000001110110000000100",
			1381 => "00000000001011100001010110100101",
			1382 => "00000000000000000001010110100101",
			1383 => "00000000000000000001010110100101",
			1384 => "11111110101001110001010110100101",
			1385 => "0000000000000000000110100000001100",
			1386 => "0000001001000000001100100000001000",
			1387 => "0000001000000000001011000100000100",
			1388 => "11111111010000000001010111110001",
			1389 => "00000000000000000001010111110001",
			1390 => "11111110011001110001010111110001",
			1391 => "0000001101000000001010011100001100",
			1392 => "0000001001000000001100100000001000",
			1393 => "0000001011000000001010111000000100",
			1394 => "00000001101011100001010111110001",
			1395 => "00000000000111110001010111110001",
			1396 => "00000000000000000001010111110001",
			1397 => "0000000110000000001100011000001000",
			1398 => "0000000010000000000010000100000100",
			1399 => "00000001101101100001010111110001",
			1400 => "00000000000000000001010111110001",
			1401 => "0000000010000000000011001000000100",
			1402 => "00000001010111110001010111110001",
			1403 => "11111110011110100001010111110001",
			1404 => "0000001001000000001100100000011100",
			1405 => "0000001110000000001001101000001100",
			1406 => "0000000000000000001111010000001000",
			1407 => "0000001001000000001100100000000100",
			1408 => "00000000000000000001011000110101",
			1409 => "11111111101000110001011000110101",
			1410 => "00000000100100100001011000110101",
			1411 => "0000000010000000001001100000001100",
			1412 => "0000001100000000001101010100001000",
			1413 => "0000000001000000001110011100000100",
			1414 => "00000001011001100001011000110101",
			1415 => "00000000000000000001011000110101",
			1416 => "00000000000000000001011000110101",
			1417 => "00000000000000000001011000110101",
			1418 => "0000001010000000000010111100000100",
			1419 => "11111110100000100001011000110101",
			1420 => "00000000000000000001011000110101",
			1421 => "0000001001000000001100100000011000",
			1422 => "0000000111000000001110001100000100",
			1423 => "11111111001110100001011001110001",
			1424 => "0000000010000000001100010100000100",
			1425 => "00000001100110100001011001110001",
			1426 => "0000001101000000000100000100001000",
			1427 => "0000000001000000001110011100000100",
			1428 => "00000000000000000001011001110001",
			1429 => "11111111010011000001011001110001",
			1430 => "0000001101000000000000011100000100",
			1431 => "00000000101100010001011001110001",
			1432 => "00000000000000000001011001110001",
			1433 => "0000001010000000000010111100000100",
			1434 => "11111110011010110001011001110001",
			1435 => "00000000000000000001011001110001",
			1436 => "0000000000000000001101000100011000",
			1437 => "0000001001000000001100100000010100",
			1438 => "0000000110000000000111101000001000",
			1439 => "0000001111000000001001110000000100",
			1440 => "00000000000000000001011010111101",
			1441 => "00000010000000110001011010111101",
			1442 => "0000000001000000001110011100001000",
			1443 => "0000001001000000001100100000000100",
			1444 => "00000000001001110001011010111101",
			1445 => "00000000000000000001011010111101",
			1446 => "11111110101001100001011010111101",
			1447 => "11111110011001100001011010111101",
			1448 => "0000000010000000001100010100000100",
			1449 => "00000001101010000001011010111101",
			1450 => "0000000110000000001100011000000100",
			1451 => "00000010001001000001011010111101",
			1452 => "0000000100000000000011100100000100",
			1453 => "11111110011110100001011010111101",
			1454 => "00000000000000000001011010111101",
			1455 => "0000000000000000000101100100000100",
			1456 => "11111110011011100001011011111001",
			1457 => "0000000001000000001110011100010100",
			1458 => "0000001100000000001101010100010000",
			1459 => "0000001111000000000111001000001100",
			1460 => "0000000000000000000110100000001000",
			1461 => "0000000000000000001110101100000100",
			1462 => "00000000100111100001011011111001",
			1463 => "00000000000000000001011011111001",
			1464 => "00000001011111000001011011111001",
			1465 => "00000000000000000001011011111001",
			1466 => "00000000000000000001011011111001",
			1467 => "0000001111000000000000001100000100",
			1468 => "00000000001010010001011011111001",
			1469 => "11111111010010110001011011111001",
			1470 => "0000000100000000000010100000000100",
			1471 => "11111110011100100001011100111101",
			1472 => "0000000010000000001010001000001100",
			1473 => "0000000011000000000001110100000100",
			1474 => "00000000000000000001011100111101",
			1475 => "0000001001000000001100100000000100",
			1476 => "00000001111100000001011100111101",
			1477 => "00000000000000000001011100111101",
			1478 => "0000001000000000001100101100000100",
			1479 => "11111111100101110001011100111101",
			1480 => "0000000001000000001110011100001100",
			1481 => "0000001100000000000001111100001000",
			1482 => "0000000010000000001110110100000100",
			1483 => "00000001001011000001011100111101",
			1484 => "00000000000000000001011100111101",
			1485 => "00000000000000000001011100111101",
			1486 => "00000000000000000001011100111101",
			1487 => "0000000000000000000110100000001100",
			1488 => "0000001001000000001100100000001000",
			1489 => "0000001111000000000101101100000100",
			1490 => "11111111001001000001011110010001",
			1491 => "00000000000000000001011110010001",
			1492 => "11111110011001100001011110010001",
			1493 => "0000001101000000001010011100001000",
			1494 => "0000001001000000001100100000000100",
			1495 => "00000001101011110001011110010001",
			1496 => "00000000000000000001011110010001",
			1497 => "0000000010000000000011001000000100",
			1498 => "00000001100010100001011110010001",
			1499 => "0000000100000000000101101000001100",
			1500 => "0000001110000000000111000100000100",
			1501 => "11111110011100100001011110010001",
			1502 => "0000001101000000000001011000000100",
			1503 => "00000000001111010001011110010001",
			1504 => "00000000000000000001011110010001",
			1505 => "0000000010000000000010000100000100",
			1506 => "00000001110010100001011110010001",
			1507 => "00000000000000000001011110010001",
			1508 => "0000000000000000001101000100001100",
			1509 => "0000001001000000001100100000001000",
			1510 => "0000000011000000001011010100000100",
			1511 => "11111110101110010001011111110101",
			1512 => "00000001010100100001011111110101",
			1513 => "11111110011001010001011111110101",
			1514 => "0000000010000000000110010000011100",
			1515 => "0000001100000000001010111100010000",
			1516 => "0000001111000000000001111100001100",
			1517 => "0000001111000000000000001100000100",
			1518 => "00000001101110100001011111110101",
			1519 => "0000001101000000001010011100000100",
			1520 => "00000001011001100001011111110101",
			1521 => "00000000000000000001011111110101",
			1522 => "00000011000000010001011111110101",
			1523 => "0000000010000000000011001000000100",
			1524 => "00000001011011100001011111110101",
			1525 => "0000001011000000001110110000000100",
			1526 => "00000000100101110001011111110101",
			1527 => "11111111000001100001011111110101",
			1528 => "0000000111000000000111001000001000",
			1529 => "0000001001000000001100100000000100",
			1530 => "00000010011100000001011111110101",
			1531 => "11111110111011000001011111110101",
			1532 => "11111110011110000001011111110101",
			1533 => "0000001001000000001100100000100100",
			1534 => "0000000010000000001010001000001000",
			1535 => "0000000101000000001110110000000100",
			1536 => "00000000000000000001100001000001",
			1537 => "00000001000010110001100001000001",
			1538 => "0000001111000000000001111100001100",
			1539 => "0000000110000000001100011000000100",
			1540 => "00000000000000000001100001000001",
			1541 => "0000001010000000000010111100000100",
			1542 => "11111111110101010001100001000001",
			1543 => "00000000000000000001100001000001",
			1544 => "0000001010000000001111000100000100",
			1545 => "00000000000000000001100001000001",
			1546 => "0000001111000000001010111000001000",
			1547 => "0000000111000000001110110000000100",
			1548 => "00000000010000000001100001000001",
			1549 => "00000000000000000001100001000001",
			1550 => "00000000000000000001100001000001",
			1551 => "11111110101000010001100001000001",
			1552 => "0000000000000000001110101000011000",
			1553 => "0000000001000000001110011100001100",
			1554 => "0000000000000000001001010100000100",
			1555 => "11111110011001000001100010101101",
			1556 => "0000001010000000001101010000000100",
			1557 => "00000101011101010001100010101101",
			1558 => "11111110110001010001100010101101",
			1559 => "0000001010000000000010011000000100",
			1560 => "11111110010110110001100010101101",
			1561 => "0000001000000000001100110000000100",
			1562 => "11111110100111110001100010101101",
			1563 => "00000001111101110001100010101101",
			1564 => "0000000010000000001110110100011100",
			1565 => "0000001100000000001101010100010100",
			1566 => "0000001110000000000110001000010000",
			1567 => "0000000011000000000011111100001100",
			1568 => "0000001111000000001010111100001000",
			1569 => "0000001111000000000100001000000100",
			1570 => "00000011010111100001100010101101",
			1571 => "00000001010110100001100010101101",
			1572 => "00000110110000010001100010101101",
			1573 => "00000000101010000001100010101101",
			1574 => "00000101110011000001100010101101",
			1575 => "0000000010000000000010000000000100",
			1576 => "00000010110101110001100010101101",
			1577 => "11111110011101000001100010101101",
			1578 => "11111110011011100001100010101101",
			1579 => "0000000000000000001101000100001100",
			1580 => "0000001001000000001100100000001000",
			1581 => "0000000011000000001011010100000100",
			1582 => "11111110110010000001100100100011",
			1583 => "00000001001011100001100100100011",
			1584 => "11111110011001010001100100100011",
			1585 => "0000001111000000000111001000101100",
			1586 => "0000001100000000001010111100011100",
			1587 => "0000000001000000001110011100010000",
			1588 => "0000001110000000000110001000001100",
			1589 => "0000000011000000000010011000000100",
			1590 => "00000001101110010001100100100011",
			1591 => "0000000011000000000010111100000100",
			1592 => "00000000111000010001100100100011",
			1593 => "00000000000000000001100100100011",
			1594 => "00000010100110100001100100100011",
			1595 => "0000000011000000000010011000000100",
			1596 => "00000001100100010001100100100011",
			1597 => "0000000100000000000101111100000100",
			1598 => "00000000000000000001100100100011",
			1599 => "11111110101001100001100100100011",
			1600 => "0000000110000000001010011000000100",
			1601 => "00000001100011100001100100100011",
			1602 => "0000000110000000001101011000001000",
			1603 => "0000001011000000001010111000000100",
			1604 => "00000000000000000001100100100011",
			1605 => "11111110100111010001100100100011",
			1606 => "00000000000000000001100100100011",
			1607 => "11111110101100010001100100100011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(530, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(1062, initial_addr_3'length));
	end generate gen_rom_0;

	gen_rom_1: if SELECT_ROM = 1 generate
		bank <= (
			0 => "00000000000000000000000000000101",
			1 => "00000000000000000000000000001001",
			2 => "00000000000000000000000000001101",
			3 => "00000000000000000000000000010001",
			4 => "00000000000000000000000000010101",
			5 => "00000000000000000000000000011001",
			6 => "00000000000000000000000000011101",
			7 => "00000000000000000000000000100001",
			8 => "00000000000000000000000000100101",
			9 => "00000000000000000000000000101001",
			10 => "00000000000000000000000000101101",
			11 => "00000000000000000000000000110001",
			12 => "00000000000000000000000000110101",
			13 => "00000000000000000000000000111001",
			14 => "00000000000000000000000000111101",
			15 => "00000000000000000000000001000001",
			16 => "00000000000000000000000001000101",
			17 => "00000000000000000000000001001001",
			18 => "00000000000000000000000001001101",
			19 => "00000000000000000000000001010001",
			20 => "00000000000000000000000001010101",
			21 => "00000000000000000000000001011001",
			22 => "00000000000000000000000001011101",
			23 => "00000000000000000000000001100001",
			24 => "00000000000000000000000001100101",
			25 => "00000000000000000000000001101001",
			26 => "00000000000000000000000001101101",
			27 => "00000000000000000000000001110001",
			28 => "00000000000000000000000001110101",
			29 => "00000000000000000000000001111001",
			30 => "00000000000000000000000001111101",
			31 => "00000000000000000000000010000001",
			32 => "00000000000000000000000010000101",
			33 => "00000000000000000000000010001001",
			34 => "00000000000000000000000010001101",
			35 => "00000000000000000000000010010001",
			36 => "00000000000000000000000010010101",
			37 => "00000000000000000000000010011001",
			38 => "0000000111000000000001111100000100",
			39 => "11111111001101110000000010100101",
			40 => "00000000000000000000000010100101",
			41 => "0000000100000000000010010000000100",
			42 => "11111111101001000000000010110001",
			43 => "00000000000000000000000010110001",
			44 => "0000000001000000000110000000000100",
			45 => "00000000000000000000000010111101",
			46 => "11111111101010010000000010111101",
			47 => "0000001001000000001110100000000100",
			48 => "00000000000000000000000011001001",
			49 => "11111111110100010000000011001001",
			50 => "0000001001000000000000011000000100",
			51 => "00000000000000000000000011010101",
			52 => "11111111110111010000000011010101",
			53 => "0000000111000000000001111100000100",
			54 => "11111111111001010000000011100001",
			55 => "00000000000000000000000011100001",
			56 => "0000000101000000000110100100001000",
			57 => "0000000100000000001111111000000100",
			58 => "11111111001011010000000011110101",
			59 => "00000000000000000000000011110101",
			60 => "00000000000000000000000011110101",
			61 => "0000000001000000000000011000001000",
			62 => "0000000010000000001010001000000100",
			63 => "00000000000000000000000100001001",
			64 => "00000000000001100000000100001001",
			65 => "11111111010110010000000100001001",
			66 => "0000000111000000000111001000001000",
			67 => "0000000010000000001100010000000100",
			68 => "11111111111011110000000100011101",
			69 => "00000000000000000000000100011101",
			70 => "00000000000000000000000100011101",
			71 => "0000001011000000001110001100001000",
			72 => "0000001110000000001001101000000100",
			73 => "00000000000000000000000100111001",
			74 => "11111111100000010000000100111001",
			75 => "0000000110000000001101011000000100",
			76 => "00000000000001110000000100111001",
			77 => "00000000000000000000000100111001",
			78 => "0000001001000000001110100000001000",
			79 => "0000000000000000000111100000000100",
			80 => "00000000000100100000000101010101",
			81 => "00000000000000000000000101010101",
			82 => "0000000100000000000101001100000100",
			83 => "11111111110100100000000101010101",
			84 => "00000000000000000000000101010101",
			85 => "0000001011000000001110001100000100",
			86 => "11111111100011100000000101110001",
			87 => "0000000110000000001101011000001000",
			88 => "0000000110000000001100011000000100",
			89 => "00000000000000000000000101110001",
			90 => "00000000001010110000000101110001",
			91 => "00000000000000000000000101110001",
			92 => "0000000111000000000001111100000100",
			93 => "11111111100111100000000110001101",
			94 => "0000000010000000001010001000000100",
			95 => "00000000000000000000000110001101",
			96 => "0000000010000000001100111000000100",
			97 => "00000000001010110000000110001101",
			98 => "00000000000000000000000110001101",
			99 => "0000001101000000001010011100001100",
			100 => "0000001100000000000100001000001000",
			101 => "0000001011000000001010111000000100",
			102 => "11111111111000000000000110101001",
			103 => "00000000000000000000000110101001",
			104 => "00000000000000000000000110101001",
			105 => "00000000000000000000000110101001",
			106 => "0000000111000000001110001100001000",
			107 => "0000000100000000001111111000000100",
			108 => "11111111001000000000000111001101",
			109 => "00000000000000000000000111001101",
			110 => "0000000110000000001101011000001000",
			111 => "0000000110000000001100011000000100",
			112 => "00000000000000000000000111001101",
			113 => "00000000001101010000000111001101",
			114 => "00000000000000000000000111001101",
			115 => "0000000100000000000010010000000100",
			116 => "11111110111001100000000111110001",
			117 => "0000001111000000001010111000000100",
			118 => "00000000000000000000000111110001",
			119 => "0000001100000000001001110000000100",
			120 => "00000000000000000000000111110001",
			121 => "0000000001000000000010001100000100",
			122 => "00000000100101100000000111110001",
			123 => "00000000000000000000000111110001",
			124 => "0000000010000000000011001000000100",
			125 => "11111111110110010000001000010101",
			126 => "0000000001000000000110000000001100",
			127 => "0000001001000000001100100000000100",
			128 => "00000000000000000000001000010101",
			129 => "0000001110000000000001110000000100",
			130 => "00000000000000000000001000010101",
			131 => "00000000000110110000001000010101",
			132 => "00000000000000000000001000010101",
			133 => "0000000111000000000001111100000100",
			134 => "11111111110011000000001000111001",
			135 => "0000000001000000001001111000001100",
			136 => "0000001001000000001100100000000100",
			137 => "00000000000000000000001000111001",
			138 => "0000001101000000000001101000000100",
			139 => "00000000000000000000001000111001",
			140 => "00000000000101110000001000111001",
			141 => "00000000000000000000001000111001",
			142 => "0000000111000000001110001100001000",
			143 => "0000000100000000000000100100000100",
			144 => "11111110110010010000001001100101",
			145 => "00000000000000000000001001100101",
			146 => "0000000001000000000010001100001100",
			147 => "0000001111000000000100001000000100",
			148 => "00000000000000000000001001100101",
			149 => "0000001000000000001101111000000100",
			150 => "00000000101010110000001001100101",
			151 => "00000000000000000000001001100101",
			152 => "00000000000000000000001001100101",
			153 => "0000000001000000000110000000010100",
			154 => "0000001111000000001101010100001000",
			155 => "0000000110000000001100011000000100",
			156 => "11111111111010110000001010010001",
			157 => "00000000000000000000001010010001",
			158 => "0000001100000000000011011100000100",
			159 => "00000000000000000000001010010001",
			160 => "0000000001000000001110011100000100",
			161 => "00000000000000000000001010010001",
			162 => "00000000011010110000001010010001",
			163 => "11111110111101000000001010010001",
			164 => "0000000100000000000101001100000100",
			165 => "11111110101110000000001010111101",
			166 => "0000000110000000001100011000000100",
			167 => "00000000000000000000001010111101",
			168 => "0000000000000000001111010000001100",
			169 => "0000001111000000000100010000001000",
			170 => "0000001111000000001101111000000100",
			171 => "00000000000000000000001010111101",
			172 => "00000000110111010000001010111101",
			173 => "00000000000000000000001010111101",
			174 => "00000000000000000000001010111101",
			175 => "0000000001000000000110000000011000",
			176 => "0000001111000000001101010100001000",
			177 => "0000000110000000001100011000000100",
			178 => "11111111111101010000001011110001",
			179 => "00000000000000000000001011110001",
			180 => "0000000010000000000101110000000100",
			181 => "00000000000000000000001011110001",
			182 => "0000000011000000001111000100000100",
			183 => "00000000000000000000001011110001",
			184 => "0000000000000000001011000100000100",
			185 => "00000000000000000000001011110001",
			186 => "00000000010111000000001011110001",
			187 => "11111110111111010000001011110001",
			188 => "0000001001000000001100110100011100",
			189 => "0000001101000000000110100100001100",
			190 => "0000000011000000000011111100001000",
			191 => "0000001011000000001010111100000100",
			192 => "11111111011000110000001100101101",
			193 => "00000000000000000000001100101101",
			194 => "00000000000000000000001100101101",
			195 => "0000000010000000001010001000000100",
			196 => "00000000000000000000001100101101",
			197 => "0000000100000000000101101000001000",
			198 => "0000001001000000001100100000000100",
			199 => "00000000000000000000001100101101",
			200 => "00000001000010100000001100101101",
			201 => "00000000000000000000001100101101",
			202 => "11111110100011110000001100101101",
			203 => "0000000001000000000110000000011100",
			204 => "0000001100000000000100001000010000",
			205 => "0000000011000000001100110000001100",
			206 => "0000000111000000000111001000001000",
			207 => "0000001011000000001110110000000100",
			208 => "11111111100101010000001101101001",
			209 => "00000000000000000000001101101001",
			210 => "00000000000000000000001101101001",
			211 => "00000000000000000000001101101001",
			212 => "0000000010000000000011001000000100",
			213 => "00000000000000000000001101101001",
			214 => "0000000100000000000011100100000100",
			215 => "00000000101101000000001101101001",
			216 => "00000000000000000000001101101001",
			217 => "11111110101011100000001101101001",
			218 => "0000000100000000001111111100011000",
			219 => "0000000100000000000100100100001100",
			220 => "0000001001000000001100110100001000",
			221 => "0000001001000000000110000000000100",
			222 => "11111110011101110000001111001101",
			223 => "11111110110110100000001111001101",
			224 => "11111110010101010000001111001101",
			225 => "0000000101000000001000011000000100",
			226 => "11111110010101110000001111001101",
			227 => "0000000010000000000101100000000100",
			228 => "00000011011111010000001111001101",
			229 => "11111110011010110000001111001101",
			230 => "0000001111000000000000001100001100",
			231 => "0000001001000000001100100000000100",
			232 => "11111110010110100000001111001101",
			233 => "0000001100000000001110001100000100",
			234 => "11111110100111100000001111001101",
			235 => "00000011011100010000001111001101",
			236 => "0000001001000000001100100000001000",
			237 => "0000000000000000001001010000000100",
			238 => "11111111110011010000001111001101",
			239 => "11111110111010110000001111001101",
			240 => "0000000011000000000010011000000100",
			241 => "00000010100011000000001111001101",
			242 => "00000011100010010000001111001101",
			243 => "0000000100000000000101001100000100",
			244 => "11111110101100010000010000000001",
			245 => "0000000010000000001010001000000100",
			246 => "00000000000000000000010000000001",
			247 => "0000000100000000000101101000010000",
			248 => "0000001111000000001001010100001100",
			249 => "0000001001000000001100100000000100",
			250 => "00000000000000000000010000000001",
			251 => "0000000101000000001010111000000100",
			252 => "00000000000000000000010000000001",
			253 => "00000001000000100000010000000001",
			254 => "00000000000000000000010000000001",
			255 => "00000000000000000000010000000001",
			256 => "0000000100000000000010010000000100",
			257 => "11111110100000010000010001000101",
			258 => "0000001100000000000100001000001100",
			259 => "0000000000000000001011000100000100",
			260 => "00000000000000000000010001000101",
			261 => "0000000110000000000100110100000100",
			262 => "11111111011100110000010001000101",
			263 => "00000000000000000000010001000101",
			264 => "0000000110000000001101011000010000",
			265 => "0000000000000000000101001000001100",
			266 => "0000001111000000000000001100000100",
			267 => "00000000000000000000010001000101",
			268 => "0000000010000000001000101000000100",
			269 => "00000001000111100000010001000101",
			270 => "00000000000000000000010001000101",
			271 => "00000000000000000000010001000101",
			272 => "00000000000000000000010001000101",
			273 => "0000000100000000001111111100011000",
			274 => "0000000100000000000010010000000100",
			275 => "11111110011001110000010010101001",
			276 => "0000001010000000001100000100001100",
			277 => "0000001100000000000110000100000100",
			278 => "11111110111000100000010010101001",
			279 => "0000001111000000001111010000000100",
			280 => "00000001111101100000010010101001",
			281 => "11111111101101010000010010101001",
			282 => "0000000100000000001101100100000100",
			283 => "11111110100110110000010010101001",
			284 => "11111111111011100000010010101001",
			285 => "0000000000000000000111100000001100",
			286 => "0000000011000000001111000100000100",
			287 => "11111111010000100000010010101001",
			288 => "0000001111000000000000001100000100",
			289 => "00000000000000000000010010101001",
			290 => "00000001100110010000010010101001",
			291 => "0000000110000000001100011000000100",
			292 => "11111110011110110000010010101001",
			293 => "0000001010000000000010111100001000",
			294 => "0000000010000000001100010100000100",
			295 => "00000000000000000000010010101001",
			296 => "00000001011111010000010010101001",
			297 => "11111110111001110000010010101001",
			298 => "0000000100000000001111111100011000",
			299 => "0000000001000000000000011000010100",
			300 => "0000000001000000001110011100001000",
			301 => "0000001010000000001100000100000100",
			302 => "00000000000000000000010100010101",
			303 => "11111110110101010000010100010101",
			304 => "0000001010000000001001101000000100",
			305 => "11111111101101010000010100010101",
			306 => "0000000001000000001110011100000100",
			307 => "00000000000000000000010100010101",
			308 => "00000000010011000000010100010101",
			309 => "11111110011010000000010100010101",
			310 => "0000000010000000000011001000010000",
			311 => "0000000000000000001101000100001100",
			312 => "0000001010000000000001110100001000",
			313 => "0000001010000000000111000100000100",
			314 => "11111111100001100000010100010101",
			315 => "00000000000000000000010100010101",
			316 => "00000000101001110000010100010101",
			317 => "11111110011111110000010100010101",
			318 => "0000000011000000001111000100000100",
			319 => "11111111100010110000010100010101",
			320 => "0000000100000000000101101000000100",
			321 => "00000001100100100000010100010101",
			322 => "0000001111000000001010111100000100",
			323 => "11111111100101110000010100010101",
			324 => "00000000011001010000010100010101",
			325 => "0000001001000000000000011000101000",
			326 => "0000000010000000001010001000001100",
			327 => "0000001001000000001100100000001000",
			328 => "0000000001000000001110011100000100",
			329 => "11111110011110100000010101111001",
			330 => "00000000000000000000010101111001",
			331 => "00000000000000000000010101111001",
			332 => "0000000001000000001110011100010100",
			333 => "0000000110000000001100011000001000",
			334 => "0000000000000000001100100100000100",
			335 => "00000000000000000000010101111001",
			336 => "11111110110110000000010101111001",
			337 => "0000000111000000000001111100000100",
			338 => "11111111010101110000010101111001",
			339 => "0000000000000000001111010000000100",
			340 => "00000001001011010000010101111001",
			341 => "00000000000000000000010101111001",
			342 => "0000000101000000001010111000000100",
			343 => "00000000000000000000010101111001",
			344 => "00000001100000000000010101111001",
			345 => "0000000000000000000110110100001000",
			346 => "0000000001000000001100100000000100",
			347 => "00000000000000000000010101111001",
			348 => "11111110011101010000010101111001",
			349 => "00000000000000000000010101111001",
			350 => "0000000100000000000010010000000100",
			351 => "11111110011010110000010111000101",
			352 => "0000000111000000001110001100001000",
			353 => "0000000100000000001101001100000100",
			354 => "11111110011100100000010111000101",
			355 => "00000000000000000000010111000101",
			356 => "0000000110000000001101011000010100",
			357 => "0000000000000000001100100100001000",
			358 => "0000000010000000000101110000000100",
			359 => "00000000000000000000010111000101",
			360 => "00000001100101110000010111000101",
			361 => "0000000110000000001100011000000100",
			362 => "11111110101011100000010111000101",
			363 => "0000000010000000001100010100000100",
			364 => "00000000000000000000010111000101",
			365 => "00000001001011000000010111000101",
			366 => "0000000100000000001111111000000100",
			367 => "11111111000001010000010111000101",
			368 => "00000000000000000000010111000101",
			369 => "0000000100000000000010010000000100",
			370 => "11111110011101100000011000001001",
			371 => "0000001101000000000011100000000100",
			372 => "11111111000000110000011000001001",
			373 => "0000001001000000001100100000010100",
			374 => "0000000110000000001100011000001000",
			375 => "0000000000000000000010110100000100",
			376 => "00000000000000000000011000001001",
			377 => "11111110111101010000011000001001",
			378 => "0000000010000000001010001000000100",
			379 => "00000000000000000000011000001001",
			380 => "0000000000000000000010011100000100",
			381 => "00000000110100010000011000001001",
			382 => "00000000000000000000011000001001",
			383 => "0000001001000000000111100100000100",
			384 => "00000001010110010000011000001001",
			385 => "11111111110100110000011000001001",
			386 => "0000000100000000001111111100010000",
			387 => "0000000001000000000000011000001100",
			388 => "0000000101000000000100011000000100",
			389 => "11111110011001000000011001011101",
			390 => "0000000000000000001001001000000100",
			391 => "00000011111001110000011001011101",
			392 => "00000001101100010000011001011101",
			393 => "11111110011000100000011001011101",
			394 => "0000000011000000001111000100000100",
			395 => "11111110011001000000011001011101",
			396 => "0000001010000000000010111100010100",
			397 => "0000001001000000001100100000000100",
			398 => "11111110011011100000011001011101",
			399 => "0000000010000000000100101000000100",
			400 => "11111111011111100000011001011101",
			401 => "0000000100000000000011100100001000",
			402 => "0000000001000000001100100000000100",
			403 => "00000001111001110000011001011101",
			404 => "00000001001001000000011001011101",
			405 => "00000000010110110000011001011101",
			406 => "11111110011111010000011001011101",
			407 => "0000000000000000001010001100010000",
			408 => "0000000001000000000110000000001100",
			409 => "0000000101000000000100011000000100",
			410 => "11111110011010010000011011000001",
			411 => "0000001110000000001111000100000100",
			412 => "00000001011101010000011011000001",
			413 => "00000010111111000000011011000001",
			414 => "11111110011001000000011011000001",
			415 => "0000000011000000001111000100000100",
			416 => "11111110011101010000011011000001",
			417 => "0000001001000000001100100000001100",
			418 => "0000000110000000001100011000000100",
			419 => "11111110001001010000011011000001",
			420 => "0000001010000000000010011000000100",
			421 => "00000001110100100000011011000001",
			422 => "11111111111011100000011011000001",
			423 => "0000000000000000000101001000001100",
			424 => "0000000001000000001011101000001000",
			425 => "0000000010000000000111111100000100",
			426 => "00000000001000110000011011000001",
			427 => "00000001101100000000011011000001",
			428 => "11111111011000100000011011000001",
			429 => "0000000110000000001010011000000100",
			430 => "11111110101010110000011011000001",
			431 => "00000001010100000000011011000001",
			432 => "0000001001000000000000011000100100",
			433 => "0000001111000000000111001000011100",
			434 => "0000000110000000001100011000001000",
			435 => "0000001001000000001100100000000100",
			436 => "11111111001111110000011100100101",
			437 => "00000000000000000000011100100101",
			438 => "0000000110000000001101011000010000",
			439 => "0000000000000000001111010000001100",
			440 => "0000000010000000001010001000000100",
			441 => "00000000000000000000011100100101",
			442 => "0000000011000000000000111000000100",
			443 => "00000000110011100000011100100101",
			444 => "00000000000000000000011100100101",
			445 => "00000000000000000000011100100101",
			446 => "00000000000000000000011100100101",
			447 => "0000000101000000001010111000000100",
			448 => "00000000000000000000011100100101",
			449 => "00000001000111010000011100100101",
			450 => "0000000110000000001110010100000100",
			451 => "00000000000000000000011100100101",
			452 => "0000001000000000001000111000001000",
			453 => "0000000001000000001100100000000100",
			454 => "00000000000000000000011100100101",
			455 => "11111110100010100000011100100101",
			456 => "00000000000000000000011100100101",
			457 => "0000000001000000001100100000101000",
			458 => "0000001111000000001010111000100000",
			459 => "0000000110000000001100011000001100",
			460 => "0000001111000000000111001000001000",
			461 => "0000001100000000000001111100000100",
			462 => "11111111101101110000011110001001",
			463 => "00000000000000000000011110001001",
			464 => "00000000000000000000011110001001",
			465 => "0000000110000000001101011000010000",
			466 => "0000000010000000001010001000000100",
			467 => "00000000000000000000011110001001",
			468 => "0000000100000000000011100100001000",
			469 => "0000000101000000000100000100000100",
			470 => "00000000101001010000011110001001",
			471 => "00000000000000000000011110001001",
			472 => "00000000000000000000011110001001",
			473 => "00000000000000000000011110001001",
			474 => "0000000101000000001010111000000100",
			475 => "00000000000000000000011110001001",
			476 => "00000000110100110000011110001001",
			477 => "0000000100000000001101001100001000",
			478 => "0000000110000000001110010100000100",
			479 => "00000000000000000000011110001001",
			480 => "11111110100011100000011110001001",
			481 => "00000000000000000000011110001001",
			482 => "0000000100000000000010010000000100",
			483 => "11111110011010100000011111001101",
			484 => "0000001101000000000100011000000100",
			485 => "11111110011000010000011111001101",
			486 => "0000000110000000001001100100011000",
			487 => "0000000000000000001100100100001100",
			488 => "0000000010000000000101110000000100",
			489 => "00000000000000000000011111001101",
			490 => "0000000001000000000010001100000100",
			491 => "00000001101000010000011111001101",
			492 => "00000000000000000000011111001101",
			493 => "0000000110000000001100011000000100",
			494 => "11111110011111100000011111001101",
			495 => "0000000010000000001100010100000100",
			496 => "11111111010101000000011111001101",
			497 => "00000001010011100000011111001101",
			498 => "11111110110001000000011111001101",
			499 => "0000000100000000001111111100010100",
			500 => "0000000100000000000010010000000100",
			501 => "11111110011001010000100000110001",
			502 => "0000001010000000001100000100001100",
			503 => "0000001100000000000110000100000100",
			504 => "11111110101000110000100000110001",
			505 => "0000001110000000001010111000000100",
			506 => "00000010100010100000100000110001",
			507 => "11111111001001100000100000110001",
			508 => "11111110101010110000100000110001",
			509 => "0000000011000000001111000100000100",
			510 => "11111110100001110000100000110001",
			511 => "0000000110000000001011001100011000",
			512 => "0000001001000000001100100000010000",
			513 => "0000000110000000001100011000001000",
			514 => "0000000110000000001100011000000100",
			515 => "11111110000111010000100000110001",
			516 => "00000000000000000000100000110001",
			517 => "0000001010000000000010111100000100",
			518 => "00000001100110100000100000110001",
			519 => "00000000000000000000100000110001",
			520 => "0000001000000000001101111000000100",
			521 => "00000001101000100000100000110001",
			522 => "00000000001110010000100000110001",
			523 => "11111111111011000000100000110001",
			524 => "0000000000000000001010001100001100",
			525 => "0000001001000000001110100000001000",
			526 => "0000000111000000001110001100000100",
			527 => "11111110100000000000100010011101",
			528 => "00000001110010100000100010011101",
			529 => "11111110011001100000100010011101",
			530 => "0000000011000000000010011000001100",
			531 => "0000000000000000001100100100001000",
			532 => "0000000011000000001111000100000100",
			533 => "11111111101000100000100010011101",
			534 => "00000001000000000000100010011101",
			535 => "11111110100100010000100010011101",
			536 => "0000000110000000001000010000011100",
			537 => "0000001001000000001100100000001000",
			538 => "0000001010000000000010011000000100",
			539 => "11111111011000100000100010011101",
			540 => "00000000001011110000100010011101",
			541 => "0000000010000000001010001000001000",
			542 => "0000000001000000001110011100000100",
			543 => "11111111101101010000100010011101",
			544 => "00000000010110010000100010011101",
			545 => "0000000000000000000111100000000100",
			546 => "00000001100111100000100010011101",
			547 => "0000001001000000001100100000000100",
			548 => "00000000011100100000100010011101",
			549 => "00000001010000110000100010011101",
			550 => "11111110000101110000100010011101",
			551 => "0000000100000000001111111100100000",
			552 => "0000000100000000000100100100010100",
			553 => "0000000001000000000000011000010000",
			554 => "0000001001000000001110100000001100",
			555 => "0000001001000000000000011000000100",
			556 => "11111110010111010000100100010001",
			557 => "0000001001000000000000011000000100",
			558 => "11111111011001110000100100010001",
			559 => "11111110100101110000100100010001",
			560 => "00000000000000000000100100010001",
			561 => "11111110010110000000100100010001",
			562 => "0000000101000000001000011000000100",
			563 => "11111110010110100000100100010001",
			564 => "0000000001000000001011101000000100",
			565 => "00000010111101100000100100010001",
			566 => "11111110011100010000100100010001",
			567 => "0000000011000000001111000100000100",
			568 => "11111110010110110000100100010001",
			569 => "0000000000000000001111010000010100",
			570 => "0000001001000000001100100000000100",
			571 => "11111111101011010000100100010001",
			572 => "0000001111000000000000001100000100",
			573 => "00000001110000000000100100010001",
			574 => "0000000111000000001110001100000100",
			575 => "00000011111001010000100100010001",
			576 => "0000001111000000000100001000000100",
			577 => "00000011011010110000100100010001",
			578 => "00000010111110110000100100010001",
			579 => "11111110011110110000100100010001",
			580 => "0000000100000000001111111100010100",
			581 => "0000001001000000001110100000010000",
			582 => "0000001110000000001000110000001000",
			583 => "0000001110000000000111000100000100",
			584 => "11111110100000100000100110001101",
			585 => "00000000000000000000100110001101",
			586 => "0000000000000000001011000100000100",
			587 => "00000000000000000000100110001101",
			588 => "00000001110010000000100110001101",
			589 => "11111110011001100000100110001101",
			590 => "0000000011000000000010011000001100",
			591 => "0000000000000000001100100100001000",
			592 => "0000000011000000001111000100000100",
			593 => "11111111001010010000100110001101",
			594 => "00000001000101110000100110001101",
			595 => "11111110100001010000100110001101",
			596 => "0000000001000000001100100000011100",
			597 => "0000001001000000001100100000001000",
			598 => "0000001010000000000010011000000100",
			599 => "11111111010010000000100110001101",
			600 => "00000000010001100000100110001101",
			601 => "0000000010000000001010001000001000",
			602 => "0000000001000000001110011100000100",
			603 => "11111111100110010000100110001101",
			604 => "00000000011100100000100110001101",
			605 => "0000000100000000000011100100001000",
			606 => "0000000100000000000001100000000100",
			607 => "00000001101000000000100110001101",
			608 => "00000000111111000000100110001101",
			609 => "00000000000000000000100110001101",
			610 => "11111111100010110000100110001101",
			611 => "0000000100000000000010010000000100",
			612 => "11111110011101010000100111111011",
			613 => "0000001100000000000100001000011100",
			614 => "0000000011000000000011111100001100",
			615 => "0000000111000000000111001000001000",
			616 => "0000000001000000001110011100000100",
			617 => "00000000000000000000100111111011",
			618 => "11111110111111010000100111111011",
			619 => "00000000000000000000100111111011",
			620 => "0000001001000000000000011000001100",
			621 => "0000000101000000001010111000000100",
			622 => "00000000000000000000100111111011",
			623 => "0000000101000000000100000100000100",
			624 => "00000000100110010000100111111011",
			625 => "00000000000000000000100111111011",
			626 => "00000000000000000000100111111011",
			627 => "0000000001000000000010001100010100",
			628 => "0000000001000000001110011100010000",
			629 => "0000000110000000001100011000000100",
			630 => "11111111101010110000100111111011",
			631 => "0000000110000000001101011000001000",
			632 => "0000000011000000001111000100000100",
			633 => "00000000000000000000100111111011",
			634 => "00000000100101100000100111111011",
			635 => "00000000000000000000100111111011",
			636 => "00000001010011110000100111111011",
			637 => "00000000000000000000100111111011",
			638 => "00000000000000000000100111111101",
			639 => "00000000000000000000101000000001",
			640 => "00000000000000000000101000000101",
			641 => "00000000000000000000101000001001",
			642 => "00000000000000000000101000001101",
			643 => "00000000000000000000101000010001",
			644 => "00000000000000000000101000010101",
			645 => "00000000000000000000101000011001",
			646 => "00000000000000000000101000011101",
			647 => "00000000000000000000101000100001",
			648 => "00000000000000000000101000100101",
			649 => "00000000000000000000101000101001",
			650 => "00000000000000000000101000101101",
			651 => "00000000000000000000101000110001",
			652 => "00000000000000000000101000110101",
			653 => "00000000000000000000101000111001",
			654 => "00000000000000000000101000111101",
			655 => "00000000000000000000101001000001",
			656 => "00000000000000000000101001000101",
			657 => "00000000000000000000101001001001",
			658 => "00000000000000000000101001001101",
			659 => "00000000000000000000101001010001",
			660 => "00000000000000000000101001010101",
			661 => "00000000000000000000101001011001",
			662 => "00000000000000000000101001011101",
			663 => "00000000000000000000101001100001",
			664 => "00000000000000000000101001100101",
			665 => "00000000000000000000101001101001",
			666 => "00000000000000000000101001101101",
			667 => "00000000000000000000101001110001",
			668 => "00000000000000000000101001110101",
			669 => "00000000000000000000101001111001",
			670 => "00000000000000000000101001111101",
			671 => "00000000000000000000101010000001",
			672 => "00000000000000000000101010000101",
			673 => "00000000000000000000101010001001",
			674 => "00000000000000000000101010001101",
			675 => "00000000000000000000101010010001",
			676 => "0000000111000000000001111100000100",
			677 => "11111111010000010000101010011101",
			678 => "00000000000000000000101010011101",
			679 => "0000000100000000000010010000000100",
			680 => "11111111101011000000101010101001",
			681 => "00000000000000000000101010101001",
			682 => "0000000001000000000110000000000100",
			683 => "00000000000000000000101010110101",
			684 => "11111111101101010000101010110101",
			685 => "0000001001000000001110100000000100",
			686 => "00000000000000000000101011000001",
			687 => "11111111110101100000101011000001",
			688 => "0000000001000000001100100000000100",
			689 => "00000000000000000000101011001101",
			690 => "11111111111000100000101011001101",
			691 => "0000000111000000000001111100000100",
			692 => "11111111111001110000101011011001",
			693 => "00000000000000000000101011011001",
			694 => "0000000100000000000010010000000100",
			695 => "11111111010000010000101011101101",
			696 => "0000000000000000001100100100000100",
			697 => "00000000000000010000101011101101",
			698 => "00000000000000000000101011101101",
			699 => "0000000100000000000010010000000100",
			700 => "11111111100010000000101100000001",
			701 => "0000000110000000001001100100000100",
			702 => "00000000000010000000101100000001",
			703 => "00000000000000000000101100000001",
			704 => "0000001100000000000100001000001000",
			705 => "0000001101000000001010001100000100",
			706 => "11111111110111100000101100010101",
			707 => "00000000000000000000101100010101",
			708 => "00000000000000000000101100010101",
			709 => "0000001001000000001110100000001000",
			710 => "0000000000000000000111100000000100",
			711 => "00000000000111010000101100110001",
			712 => "00000000000000000000101100110001",
			713 => "0000000100000000000101001100000100",
			714 => "11111111110010000000101100110001",
			715 => "00000000000000000000101100110001",
			716 => "0000000001000000000110000000001100",
			717 => "0000000000000000001100100100001000",
			718 => "0000000000000000001011000100000100",
			719 => "00000000000000000000101101001101",
			720 => "00000000000100010000101101001101",
			721 => "00000000000000000000101101001101",
			722 => "11111111010010110000101101001101",
			723 => "0000000111000000000001111100001100",
			724 => "0000000110000000000001111000000100",
			725 => "00000000000000000000101101101001",
			726 => "0000000100000000000000100100000100",
			727 => "11111111100100110000101101101001",
			728 => "00000000000000000000101101101001",
			729 => "00000000000000000000101101101001",
			730 => "0000001101000000001010011100001100",
			731 => "0000001100000000000100001000001000",
			732 => "0000001011000000001010111000000100",
			733 => "11111111110110010000101110000101",
			734 => "00000000000000000000101110000101",
			735 => "00000000000000000000101110000101",
			736 => "00000000000000000000101110000101",
			737 => "0000000111000000000111001000001100",
			738 => "0000001110000000001001101000000100",
			739 => "00000000000000000000101110100001",
			740 => "0000000010000000001111010100000100",
			741 => "11111111111001100000101110100001",
			742 => "00000000000000000000101110100001",
			743 => "00000000000000000000101110100001",
			744 => "0000000111000000000001111100001100",
			745 => "0000000110000000000001111000000100",
			746 => "00000000000000000000101111001101",
			747 => "0000000100000000000000100100000100",
			748 => "11111111100010110000101111001101",
			749 => "00000000000000000000101111001101",
			750 => "0000000010000000001010001000000100",
			751 => "00000000000000000000101111001101",
			752 => "0000000010000000001000101000000100",
			753 => "00000000000110100000101111001101",
			754 => "00000000000000000000101111001101",
			755 => "0000000001000000000110000000010000",
			756 => "0000001111000000001101010100000100",
			757 => "00000000000000000000101111110001",
			758 => "0000001100000000000011011100000100",
			759 => "00000000000000000000101111110001",
			760 => "0000001001000000001100100000000100",
			761 => "00000000000000000000101111110001",
			762 => "00000000010110110000101111110001",
			763 => "11111111000001110000101111110001",
			764 => "0000000010000000000011001000000100",
			765 => "11111111110111000000110000010101",
			766 => "0000000001000000000110000000001100",
			767 => "0000000001000000001110011100000100",
			768 => "00000000000000000000110000010101",
			769 => "0000001110000000000001110000000100",
			770 => "00000000000000000000110000010101",
			771 => "00000000000011100000110000010101",
			772 => "00000000000000000000110000010101",
			773 => "0000000111000000000111001000010000",
			774 => "0000001110000000001001101000000100",
			775 => "00000000000000000000110000111001",
			776 => "0000000110000000000101011100000100",
			777 => "00000000000000000000110000111001",
			778 => "0000001100000000001101010100000100",
			779 => "11111111110101100000110000111001",
			780 => "00000000000000000000110000111001",
			781 => "00000000000000000000110000111001",
			782 => "0000000111000000001110001100001000",
			783 => "0000000100000000001101001100000100",
			784 => "11111110111011000000110001100101",
			785 => "00000000000000000000110001100101",
			786 => "0000000110000000001101011000001100",
			787 => "0000001001000000001100100000000100",
			788 => "00000000000000000000110001100101",
			789 => "0000001001000000000111100100000100",
			790 => "00000000011100110000110001100101",
			791 => "00000000000000000000110001100101",
			792 => "00000000000000000000110001100101",
			793 => "0000001001000000000000011000010100",
			794 => "0000001111000000000000001100000100",
			795 => "00000000000000000000110010011001",
			796 => "0000001000000000001101111000001100",
			797 => "0000001011000000001000000000001000",
			798 => "0000000101000000001010111000000100",
			799 => "00000000000000000000110010011001",
			800 => "00000000011111110000110010011001",
			801 => "00000000000000000000110010011001",
			802 => "00000000000000000000110010011001",
			803 => "0000000111000000000111001000000100",
			804 => "11111110110100110000110010011001",
			805 => "00000000000000000000110010011001",
			806 => "0000000100000000000101001100000100",
			807 => "11111110101111110000110011000101",
			808 => "0000000110000000001100011000000100",
			809 => "00000000000000000000110011000101",
			810 => "0000001010000000000010111100001100",
			811 => "0000001111000000000100010000001000",
			812 => "0000001111000000001101111000000100",
			813 => "00000000000000000000110011000101",
			814 => "00000000110010100000110011000101",
			815 => "00000000000000000000110011000101",
			816 => "00000000000000000000110011000101",
			817 => "0000000100000000001101001100001100",
			818 => "0000000001000000001100100000001000",
			819 => "0000001100000000000000001100000100",
			820 => "11111111110111100000110100001001",
			821 => "00000000000000000000110100001001",
			822 => "11111110011110110000110100001001",
			823 => "0000000010000000001110010000001000",
			824 => "0000001001000000001100100000000100",
			825 => "11111110111011010000110100001001",
			826 => "00000000000000000000110100001001",
			827 => "0000000011000000001111000100000100",
			828 => "00000000000000000000110100001001",
			829 => "0000000100000000000011100100001000",
			830 => "0000001001000000001100100000000100",
			831 => "00000000000000000000110100001001",
			832 => "00000001011010010000110100001001",
			833 => "00000000000000000000110100001001",
			834 => "0000000111000000000001111100001000",
			835 => "0000000100000000000000100100000100",
			836 => "11111110100110010000110101000101",
			837 => "00000000000000000000110101000101",
			838 => "0000000001000000000010001100010100",
			839 => "0000001001000000001100100000010000",
			840 => "0000001110000000001001101000001000",
			841 => "0000000011000000001111000100000100",
			842 => "00000000000000000000110101000101",
			843 => "00000000000000010000110101000101",
			844 => "0000000011000000000010111100000100",
			845 => "00000000000000000000110101000101",
			846 => "11111111110000000000110101000101",
			847 => "00000000110010010000110101000101",
			848 => "11111111101010100000110101000101",
			849 => "0000001100000000001100110000000100",
			850 => "11111110111000000000110110000001",
			851 => "0000000110000000001101011000010000",
			852 => "0000001111000000000000001100000100",
			853 => "00000000000000000000110110000001",
			854 => "0000000100000000000001100000001000",
			855 => "0000000001000000001100110100000100",
			856 => "00000000101111100000110110000001",
			857 => "00000000000000000000110110000001",
			858 => "00000000000000000000110110000001",
			859 => "0000000101000000000011100000000100",
			860 => "00000000000000000000110110000001",
			861 => "0000000100000000000000100100000100",
			862 => "11111111111001000000110110000001",
			863 => "00000000000000000000110110000001",
			864 => "0000000100000000001111111100001100",
			865 => "0000000001000000000110000000001000",
			866 => "0000000101000000000100011000000100",
			867 => "11111110011010110000110111001101",
			868 => "00000010011011000000110111001101",
			869 => "11111110011001000000110111001101",
			870 => "0000000011000000001111000100000100",
			871 => "11111110011101010000110111001101",
			872 => "0000001001000000001100100000001100",
			873 => "0000000110000000001100011000000100",
			874 => "11111110001111000000110111001101",
			875 => "0000001010000000000010011000000100",
			876 => "00000001101111000000110111001101",
			877 => "00000000000000000000110111001101",
			878 => "0000000100000000000011100100001000",
			879 => "0000000000000000001001010000000100",
			880 => "00000001101001110000110111001101",
			881 => "00000000000000000000110111001101",
			882 => "00000000000000000000110111001101",
			883 => "0000000100000000000010010000000100",
			884 => "11111110100000110000111000010001",
			885 => "0000001100000000000100001000010000",
			886 => "0000000000000000001011000100000100",
			887 => "00000000000000000000111000010001",
			888 => "0000000100000000000000100100001000",
			889 => "0000000111000000000111001000000100",
			890 => "11111111011101010000111000010001",
			891 => "00000000000000000000111000010001",
			892 => "00000000000000000000111000010001",
			893 => "0000000011000000000111110000001100",
			894 => "0000000010000000000011001000000100",
			895 => "00000000000000000000111000010001",
			896 => "0000000100000000000011100100000100",
			897 => "00000001000101010000111000010001",
			898 => "00000000000000000000111000010001",
			899 => "00000000000000000000111000010001",
			900 => "0000000100000000001111111100010100",
			901 => "0000000001000000000000011000001000",
			902 => "0000000101000000001000011000000100",
			903 => "11111110010111100000111001101101",
			904 => "00000011111110100000111001101101",
			905 => "0000000001000000000110000000001000",
			906 => "0000000001000000000110000000000100",
			907 => "11111110011000010000111001101101",
			908 => "11111110110011110000111001101101",
			909 => "11111110010110110000111001101101",
			910 => "0000001111000000001101111000000100",
			911 => "11111110011000100000111001101101",
			912 => "0000000100000000000011100100010000",
			913 => "0000000101000000000100011000000100",
			914 => "00000000000000000000111001101101",
			915 => "0000001001000000001100100000000100",
			916 => "00000000001100010000111001101101",
			917 => "0000000000000000001111010000000100",
			918 => "00000010011001100000111001101101",
			919 => "11111111001000010000111001101101",
			920 => "0000000110000000001100011000000100",
			921 => "11111101101001100000111001101101",
			922 => "00000000111011100000111001101101",
			923 => "0000000100000000001101001100010000",
			924 => "0000000100000000001011100100000100",
			925 => "11111110011011000000111011001001",
			926 => "0000000111000000000001111100000100",
			927 => "11111110100010110000111011001001",
			928 => "0000001001000000000111100100000100",
			929 => "00000001000110100000111011001001",
			930 => "11111111001110100000111011001001",
			931 => "0000000010000000001110010000001000",
			932 => "0000001001000000001100100000000100",
			933 => "11111110101000110000111011001001",
			934 => "00000000000000000000111011001001",
			935 => "0000000001000000001110011100010100",
			936 => "0000000110000000001100011000001000",
			937 => "0000001010000000001101010000000100",
			938 => "00000000000000000000111011001001",
			939 => "11111110111111010000111011001001",
			940 => "0000000111000000000001111100000100",
			941 => "11111111011100100000111011001001",
			942 => "0000000000000000001111010000000100",
			943 => "00000001000111100000111011001001",
			944 => "00000000000000000000111011001001",
			945 => "00000001011110010000111011001001",
			946 => "0000001001000000000000011000100100",
			947 => "0000001111000000000111001000011100",
			948 => "0000000110000000001100011000001100",
			949 => "0000000001000000001110011100001000",
			950 => "0000001001000000001100100000000100",
			951 => "11111110111101110000111100110101",
			952 => "00000000000000000000111100110101",
			953 => "00000000000000000000111100110101",
			954 => "0000001010000000000010111100001100",
			955 => "0000000010000000001010001000000100",
			956 => "00000000000000000000111100110101",
			957 => "0000000101000000000100000100000100",
			958 => "00000000110110010000111100110101",
			959 => "00000000000000000000111100110101",
			960 => "00000000000000000000111100110101",
			961 => "0000000101000000001010111000000100",
			962 => "00000000000000000000111100110101",
			963 => "00000001001100110000111100110101",
			964 => "0000000000000000000110000100001000",
			965 => "0000000001000000000000011000000100",
			966 => "00000000000000000000111100110101",
			967 => "11111110011110000000111100110101",
			968 => "0000001100000000000100001000000100",
			969 => "11111111001011110000111100110101",
			970 => "0000000001000000000010001100000100",
			971 => "00000000011111000000111100110101",
			972 => "00000000000000000000111100110101",
			973 => "0000001001000000000000011000100100",
			974 => "0000001111000000000111001000011100",
			975 => "0000000110000000001100011000001000",
			976 => "0000001001000000001100100000000100",
			977 => "11111111001010010000111110011001",
			978 => "00000000000000000000111110011001",
			979 => "0000000110000000001101011000001100",
			980 => "0000000000000000001111010000001000",
			981 => "0000000010000000001010001000000100",
			982 => "00000000000000000000111110011001",
			983 => "00000000110100110000111110011001",
			984 => "00000000000000000000111110011001",
			985 => "0000000001000000001110011100000100",
			986 => "11111111111110000000111110011001",
			987 => "00000000000000000000111110011001",
			988 => "0000000101000000001010111000000100",
			989 => "00000000000000000000111110011001",
			990 => "00000001001010000000111110011001",
			991 => "0000000110000000001110010100000100",
			992 => "00000000000000000000111110011001",
			993 => "0000001000000000001000111000001000",
			994 => "0000000001000000001100100000000100",
			995 => "00000000000000000000111110011001",
			996 => "11111110100001010000111110011001",
			997 => "00000000000000000000111110011001",
			998 => "0000000100000000001111101100000100",
			999 => "11111110100110000000111111100101",
			1000 => "0000001100000000000100001000010000",
			1001 => "0000000011000000000011111100001100",
			1002 => "0000000001000000001110011100000100",
			1003 => "00000000000000000000111111100101",
			1004 => "0000000111000000000111001000000100",
			1005 => "11111111011110000000111111100101",
			1006 => "00000000000000000000111111100101",
			1007 => "00000000000000000000111111100101",
			1008 => "0000000010000000001010001000000100",
			1009 => "00000000000000000000111111100101",
			1010 => "0000000001000000001110011100000100",
			1011 => "00000000000000000000111111100101",
			1012 => "0000000001000000000010001100001000",
			1013 => "0000000000000000000101001000000100",
			1014 => "00000000110100100000111111100101",
			1015 => "00000000000000000000111111100101",
			1016 => "00000000000000000000111111100101",
			1017 => "0000000100000000001101001100010000",
			1018 => "0000000100000000000101001100000100",
			1019 => "11111110011100100001000001000001",
			1020 => "0000000111000000000100001000000100",
			1021 => "11111110110010000001000001000001",
			1022 => "0000000001000000001001111000000100",
			1023 => "00000000101011100001000001000001",
			1024 => "00000000000000000001000001000001",
			1025 => "0000001111000000000000001100001000",
			1026 => "0000001001000000001100100000000100",
			1027 => "11111111001011100001000001000001",
			1028 => "00000000000000000001000001000001",
			1029 => "0000000100000000000011100100010100",
			1030 => "0000001011000000001100101000000100",
			1031 => "00000000000000000001000001000001",
			1032 => "0000001011000000001000000000001100",
			1033 => "0000001010000000000010111100001000",
			1034 => "0000001001000000001100100000000100",
			1035 => "00000000000000000001000001000001",
			1036 => "00000001010101110001000001000001",
			1037 => "00000000000000000001000001000001",
			1038 => "00000000000000000001000001000001",
			1039 => "00000000000000000001000001000001",
			1040 => "0000000100000000001111111100100100",
			1041 => "0000000100000000000100100100011000",
			1042 => "0000000001000000000000011000010100",
			1043 => "0000001001000000001110100000001100",
			1044 => "0000001001000000000000011000000100",
			1045 => "11111110011000010001000010101101",
			1046 => "0000001001000000000000011000000100",
			1047 => "11111111100000000001000010101101",
			1048 => "11111110101000100001000010101101",
			1049 => "0000000000000000000111111000000100",
			1050 => "11111110110101000001000010101101",
			1051 => "00000001000000100001000010101101",
			1052 => "11111110010110100001000010101101",
			1053 => "0000000101000000001000011000000100",
			1054 => "11111110010111010001000010101101",
			1055 => "0000000001000000001011101000000100",
			1056 => "00000010100111000001000010101101",
			1057 => "11111110011110000001000010101101",
			1058 => "0000001111000000001101111000000100",
			1059 => "11111110010111110001000010101101",
			1060 => "0000000000000000001111010000001100",
			1061 => "0000000011000000001111000100000100",
			1062 => "11111110011111010001000010101101",
			1063 => "0000000001000000001110011100000100",
			1064 => "00000001011100110001000010101101",
			1065 => "00000010101001000001000010101101",
			1066 => "11111110100011000001000010101101",
			1067 => "0000000100000000001111111100010100",
			1068 => "0000000100000000000010010000000100",
			1069 => "11111110011001010001000100010001",
			1070 => "0000001010000000001100000100001100",
			1071 => "0000001100000000000110000100000100",
			1072 => "11111110100100100001000100010001",
			1073 => "0000001110000000001010111000000100",
			1074 => "00000011000111110001000100010001",
			1075 => "11111110111110010001000100010001",
			1076 => "11111110101000000001000100010001",
			1077 => "0000000011000000001111000100000100",
			1078 => "11111110011110010001000100010001",
			1079 => "0000001001000000001100100000010000",
			1080 => "0000000110000000001100011000000100",
			1081 => "11111101110101100001000100010001",
			1082 => "0000000010000000000011001000001000",
			1083 => "0000000100000000001011010000000100",
			1084 => "00000000000000000001000100010001",
			1085 => "11111111110010000001000100010001",
			1086 => "00000001101100110001000100010001",
			1087 => "0000000010000000001000101000001000",
			1088 => "0000001000000000001101111000000100",
			1089 => "00000001101010000001000100010001",
			1090 => "00000000010100110001000100010001",
			1091 => "11111111111111100001000100010001",
			1092 => "0000000100000000001111111100010000",
			1093 => "0000000001000000000000011000001100",
			1094 => "0000000101000000000100011000000100",
			1095 => "11111110011001100001000101101101",
			1096 => "0000000100000000001111110100000100",
			1097 => "00000011011011000001000101101101",
			1098 => "00000001100111000001000101101101",
			1099 => "11111110011000110001000101101101",
			1100 => "0000000011000000001111000100000100",
			1101 => "11111110011001100001000101101101",
			1102 => "0000001001000000001100100000001000",
			1103 => "0000000110000000001100011000000100",
			1104 => "11111110011010000001000101101101",
			1105 => "00000001001100000001000101101101",
			1106 => "0000000100000000000011100100010000",
			1107 => "0000001010000000000011111100001100",
			1108 => "0000000010000000000100101000000100",
			1109 => "11111111101111110001000101101101",
			1110 => "0000001001000000000000011000000100",
			1111 => "00000001110110000001000101101101",
			1112 => "00000001000001010001000101101101",
			1113 => "11111110101011010001000101101101",
			1114 => "11111111100100000001000101101101",
			1115 => "0000000100000000000010010000000100",
			1116 => "11111110011010100001000110111001",
			1117 => "0000000111000000001110001100001000",
			1118 => "0000001101000000000100011000000100",
			1119 => "11111110011100100001000110111001",
			1120 => "00000000000000000001000110111001",
			1121 => "0000000110000000001011001100011000",
			1122 => "0000000000000000001100100100001100",
			1123 => "0000000010000000000101110000000100",
			1124 => "00000000000000000001000110111001",
			1125 => "0000000001000000000110101000000100",
			1126 => "00000001100111000001000110111001",
			1127 => "00000000000000000001000110111001",
			1128 => "0000000110000000001100011000000100",
			1129 => "11111110100101100001000110111001",
			1130 => "0000000010000000001100010100000100",
			1131 => "11111111011011110001000110111001",
			1132 => "00000001010000100001000110111001",
			1133 => "11111110110110010001000110111001",
			1134 => "0000000100000000000010010000000100",
			1135 => "11111110100001100001000111111101",
			1136 => "0000000010000000000101110000000100",
			1137 => "11111111110001100001000111111101",
			1138 => "0000000110000000001101011000010100",
			1139 => "0000000100000000000001100000010000",
			1140 => "0000000111000000000110000100000100",
			1141 => "00000000000000000001000111111101",
			1142 => "0000000001000000001110100000001000",
			1143 => "0000001111000000000000001100000100",
			1144 => "00000000000000000001000111111101",
			1145 => "00000001001011010001000111111101",
			1146 => "00000000000000000001000111111101",
			1147 => "00000000000000000001000111111101",
			1148 => "0000000100000000001111111000000100",
			1149 => "11111111111010000001000111111101",
			1150 => "00000000000000000001000111111101",
			1151 => "0000000000000000000111010000011100",
			1152 => "0000000000000000001111011100010000",
			1153 => "0000000001000000000000011000001100",
			1154 => "0000000101000000000100011000000100",
			1155 => "11111110010100010001001001110001",
			1156 => "0000000000000000001011000000000100",
			1157 => "00001001110011110001001001110001",
			1158 => "00000110001111000001001001110001",
			1159 => "11111110010011110001001001110001",
			1160 => "0000000011000000000000111000000100",
			1161 => "11111110010110010001001001110001",
			1162 => "0000000001000000001101101000000100",
			1163 => "00000110010100110001001001110001",
			1164 => "11111110011100100001001001110001",
			1165 => "0000000011000000001111000100000100",
			1166 => "11111110010101000001001001110001",
			1167 => "0000001010000000000010111100010100",
			1168 => "0000001111000000001101111000000100",
			1169 => "11111110100111000001001001110001",
			1170 => "0000000000000000001111010000001100",
			1171 => "0000000110000000001001100100001000",
			1172 => "0000001101000000001001001000000100",
			1173 => "00001000100111110001001001110001",
			1174 => "00000110001000100001001001110001",
			1175 => "00000000010110000001001001110001",
			1176 => "11111110110011000001001001110001",
			1177 => "0000001110000000001001101000000100",
			1178 => "00000000001111010001001001110001",
			1179 => "11111110011001110001001001110001",
			1180 => "0000000100000000000010010000000100",
			1181 => "11111110011011100001001011001101",
			1182 => "0000000010000000000101110000001000",
			1183 => "0000001100000000000001111100000100",
			1184 => "11111110101111000001001011001101",
			1185 => "00000000000000000001001011001101",
			1186 => "0000000110000000001101011000011000",
			1187 => "0000000000000000001100100100001100",
			1188 => "0000000111000000000101101100000100",
			1189 => "00000000000000000001001011001101",
			1190 => "0000001001000000000111100100000100",
			1191 => "00000001100010110001001011001101",
			1192 => "00000000000000000001001011001101",
			1193 => "0000000110000000001100011000000100",
			1194 => "11111111000011010001001011001101",
			1195 => "0000000010000000001100010100000100",
			1196 => "00000000000000000001001011001101",
			1197 => "00000001000000100001001011001101",
			1198 => "0000000110000000001001100100000100",
			1199 => "00000000000000000001001011001101",
			1200 => "0000000111000000001110001100000100",
			1201 => "00000000000000000001001011001101",
			1202 => "11111111000001000001001011001101",
			1203 => "0000000100000000001111111100100100",
			1204 => "0000000001000000000000011000100000",
			1205 => "0000001001000000000000011000001000",
			1206 => "0000001010000000001100000100000100",
			1207 => "00000000000000000001001101011001",
			1208 => "11111110111011010001001101011001",
			1209 => "0000001000000000000011111100001100",
			1210 => "0000001010000000000110011100001000",
			1211 => "0000001010000000001010110000000100",
			1212 => "11111111110101010001001101011001",
			1213 => "00000000000100010001001101011001",
			1214 => "11111111110000100001001101011001",
			1215 => "0000001000000000000100010100001000",
			1216 => "0000001010000000001001101000000100",
			1217 => "00000000000000000001001101011001",
			1218 => "00000000010101110001001101011001",
			1219 => "00000000000000000001001101011001",
			1220 => "11111110011010010001001101011001",
			1221 => "0000000010000000000011001000001100",
			1222 => "0000001001000000001100100000000100",
			1223 => "11111110101100010001001101011001",
			1224 => "0000001010000000000111000100000100",
			1225 => "00000000000000000001001101011001",
			1226 => "00000000100110010001001101011001",
			1227 => "0000000100000000000101101000001100",
			1228 => "0000000110000000001101011000001000",
			1229 => "0000001001000000001100100000000100",
			1230 => "00000000000000000001001101011001",
			1231 => "00000001100100000001001101011001",
			1232 => "00000000000000000001001101011001",
			1233 => "0000000110000000001100011000000100",
			1234 => "11111111011100000001001101011001",
			1235 => "0000000010000000000110010000000100",
			1236 => "00000000000000000001001101011001",
			1237 => "00000000100111010001001101011001",
			1238 => "0000000100000000001111101100000100",
			1239 => "11111110100111010001001110110101",
			1240 => "0000001100000000000100001000010100",
			1241 => "0000001110000000000110001000010000",
			1242 => "0000001110000000001001101000000100",
			1243 => "00000000000000000001001110110101",
			1244 => "0000001101000000001010001100001000",
			1245 => "0000000111000000001110110000000100",
			1246 => "11111111100010010001001110110101",
			1247 => "00000000000000000001001110110101",
			1248 => "00000000000000000001001110110101",
			1249 => "00000000000000000001001110110101",
			1250 => "0000000110000000001100011000000100",
			1251 => "00000000000000000001001110110101",
			1252 => "0000000110000000001101011000010000",
			1253 => "0000001001000000001100100000000100",
			1254 => "00000000000000000001001110110101",
			1255 => "0000001111000000001101111000000100",
			1256 => "00000000000000000001001110110101",
			1257 => "0000001111000000000110110100000100",
			1258 => "00000000101111100001001110110101",
			1259 => "00000000000000000001001110110101",
			1260 => "00000000000000000001001110110101",
			1261 => "0000000100000000000010010000000100",
			1262 => "11111110011100000001010000010011",
			1263 => "0000000010000000000101110000001000",
			1264 => "0000001100000000000001111100000100",
			1265 => "11111110110111110001010000010011",
			1266 => "00000000000000000001010000010011",
			1267 => "0000000001000000000110000000100000",
			1268 => "0000000001000000001110011100010100",
			1269 => "0000000000000000001100100100001000",
			1270 => "0000001110000000001001101000000100",
			1271 => "00000000000000000001010000010011",
			1272 => "00000000101010000001010000010011",
			1273 => "0000001110000000000110001000001000",
			1274 => "0000001101000000001000011000000100",
			1275 => "00000000000000000001010000010011",
			1276 => "00000000010111100001010000010011",
			1277 => "11111111010011000001010000010011",
			1278 => "0000000101000000001010111000000100",
			1279 => "00000000000000000001010000010011",
			1280 => "0000000000000000000100101000000100",
			1281 => "00000001011111100001010000010011",
			1282 => "00000000000000000001010000010011",
			1283 => "11111111001111100001010000010011",
			1284 => "00000000000000000001010000010101",
			1285 => "00000000000000000001010000011001",
			1286 => "00000000000000000001010000011101",
			1287 => "00000000000000000001010000100001",
			1288 => "00000000000000000001010000100101",
			1289 => "00000000000000000001010000101001",
			1290 => "00000000000000000001010000101101",
			1291 => "00000000000000000001010000110001",
			1292 => "00000000000000000001010000110101",
			1293 => "00000000000000000001010000111001",
			1294 => "00000000000000000001010000111101",
			1295 => "00000000000000000001010001000001",
			1296 => "00000000000000000001010001000101",
			1297 => "00000000000000000001010001001001",
			1298 => "00000000000000000001010001001101",
			1299 => "00000000000000000001010001010001",
			1300 => "00000000000000000001010001010101",
			1301 => "00000000000000000001010001011001",
			1302 => "00000000000000000001010001011101",
			1303 => "00000000000000000001010001100001",
			1304 => "00000000000000000001010001100101",
			1305 => "00000000000000000001010001101001",
			1306 => "00000000000000000001010001101101",
			1307 => "00000000000000000001010001110001",
			1308 => "00000000000000000001010001110101",
			1309 => "00000000000000000001010001111001",
			1310 => "00000000000000000001010001111101",
			1311 => "00000000000000000001010010000001",
			1312 => "00000000000000000001010010000101",
			1313 => "00000000000000000001010010001001",
			1314 => "00000000000000000001010010001101",
			1315 => "00000000000000000001010010010001",
			1316 => "00000000000000000001010010010101",
			1317 => "00000000000000000001010010011001",
			1318 => "00000000000000000001010010011101",
			1319 => "00000000000000000001010010100001",
			1320 => "00000000000000000001010010100101",
			1321 => "00000000000000000001010010101001",
			1322 => "0000000100000000000010010000000100",
			1323 => "11111111010101000001010010110101",
			1324 => "00000000000000000001010010110101",
			1325 => "0000000111000000000110000100000100",
			1326 => "11111111101100100001010011000001",
			1327 => "00000000000000000001010011000001",
			1328 => "0000000111000000000001111100000100",
			1329 => "11111111101001100001010011001101",
			1330 => "00000000000000000001010011001101",
			1331 => "0000001001000000001110100000000100",
			1332 => "00000000000000000001010011011001",
			1333 => "11111111110110010001010011011001",
			1334 => "0000001001000000000000011000000100",
			1335 => "00000000000000000001010011100101",
			1336 => "11111111111001010001010011100101",
			1337 => "0000000111000000000001111100000100",
			1338 => "11111111111010010001010011110001",
			1339 => "00000000000000000001010011110001",
			1340 => "0000000001000000000000011000001000",
			1341 => "0000000010000000001010001000000100",
			1342 => "00000000000000000001010100000101",
			1343 => "00000000000010000001010100000101",
			1344 => "11111111010100000001010100000101",
			1345 => "0000001001000000001110100000000100",
			1346 => "00000000000000000001010100011001",
			1347 => "0000000100000000000101001100000100",
			1348 => "11111111101010100001010100011001",
			1349 => "00000000000000000001010100011001",
			1350 => "0000001011000000001110001100001000",
			1351 => "0000001110000000001001101000000100",
			1352 => "00000000000000000001010100110101",
			1353 => "11111111011110000001010100110101",
			1354 => "0000000110000000001101011000000100",
			1355 => "00000000000010000001010100110101",
			1356 => "00000000000000000001010100110101",
			1357 => "0000001001000000001110100000001000",
			1358 => "0000000000000000000111100000000100",
			1359 => "00000000000101100001010101010001",
			1360 => "00000000000000000001010101010001",
			1361 => "0000000100000000000101001100000100",
			1362 => "11111111110011010001010101010001",
			1363 => "00000000000000000001010101010001",
			1364 => "0000000001000000000000011000001100",
			1365 => "0000000110000000001100011000000100",
			1366 => "00000000000000000001010101101101",
			1367 => "0000000010000000001010001000000100",
			1368 => "00000000000000000001010101101101",
			1369 => "00000000001101000001010101101101",
			1370 => "11111111011000100001010101101101",
			1371 => "0000000111000000000001111100000100",
			1372 => "11111111100101100001010110001001",
			1373 => "0000000010000000001010001000000100",
			1374 => "00000000000000000001010110001001",
			1375 => "0000000010000000001100111000000100",
			1376 => "00000000001011010001010110001001",
			1377 => "00000000000000000001010110001001",
			1378 => "0000001101000000001010011100001100",
			1379 => "0000001100000000000100001000001000",
			1380 => "0000001011000000001010111000000100",
			1381 => "11111111110111000001010110100101",
			1382 => "00000000000000000001010110100101",
			1383 => "00000000000000000001010110100101",
			1384 => "00000000000000000001010110100101",
			1385 => "0000001100000000000100001000001100",
			1386 => "0000001101000000001010001100001000",
			1387 => "0000000111000000000111001000000100",
			1388 => "11111111110111100001010111000001",
			1389 => "00000000000000000001010111000001",
			1390 => "00000000000000000001010111000001",
			1391 => "00000000000000000001010111000001",
			1392 => "0000000111000000000110000100000100",
			1393 => "11111110110011010001010111100101",
			1394 => "0000000001000000001100110100001100",
			1395 => "0000001111000000000000001100000100",
			1396 => "00000000000000000001010111100101",
			1397 => "0000000000000000001100100100000100",
			1398 => "00000000101010000001010111100101",
			1399 => "00000000000000000001010111100101",
			1400 => "00000000000000000001010111100101",
			1401 => "0000000010000000000011001000000100",
			1402 => "11111111110101100001011000001001",
			1403 => "0000000001000000000110000000001100",
			1404 => "0000001001000000001100100000000100",
			1405 => "00000000000000000001011000001001",
			1406 => "0000001110000000000001110000000100",
			1407 => "00000000000000000001011000001001",
			1408 => "00000000000111000001011000001001",
			1409 => "00000000000000000001011000001001",
			1410 => "0000000111000000000001111100000100",
			1411 => "11111111110001110001011000101101",
			1412 => "0000000001000000001001111000001100",
			1413 => "0000001001000000001100100000000100",
			1414 => "00000000000000000001011000101101",
			1415 => "0000001101000000000001101000000100",
			1416 => "00000000000000000001011000101101",
			1417 => "00000000000110100001011000101101",
			1418 => "00000000000000000001011000101101",
			1419 => "0000001100000000000100001000010000",
			1420 => "0000001110000000001100000100000100",
			1421 => "00000000000000000001011001010001",
			1422 => "0000001101000000001010001100001000",
			1423 => "0000000111000000000111001000000100",
			1424 => "11111111110001100001011001010001",
			1425 => "00000000000000000001011001010001",
			1426 => "00000000000000000001011001010001",
			1427 => "00000000000000000001011001010001",
			1428 => "0000000111000000001110001100001000",
			1429 => "0000000100000000001111111000000100",
			1430 => "11111111000101010001011001111101",
			1431 => "00000000000000000001011001111101",
			1432 => "0000000110000000001101011000001100",
			1433 => "0000000110000000001100011000000100",
			1434 => "00000000000000000001011001111101",
			1435 => "0000000110000000001101011000000100",
			1436 => "00000000001110000001011001111101",
			1437 => "00000000000000000001011001111101",
			1438 => "00000000000000000001011001111101",
			1439 => "0000000111000000001110001100001000",
			1440 => "0000000100000000001111111000000100",
			1441 => "11111111000010100001011010110001",
			1442 => "00000000000000000001011010110001",
			1443 => "0000000110000000001101011000010000",
			1444 => "0000001001000000001100100000000100",
			1445 => "00000000000000000001011010110001",
			1446 => "0000000001000000000010001100001000",
			1447 => "0000001110000000001100000100000100",
			1448 => "00000000000000000001011010110001",
			1449 => "00000000011000110001011010110001",
			1450 => "00000000000000000001011010110001",
			1451 => "00000000000000000001011010110001",
			1452 => "0000000111000000000001111100000100",
			1453 => "11111111110000010001011011011101",
			1454 => "0000000001000000001001111000010000",
			1455 => "0000000010000000001010001000000100",
			1456 => "00000000000000000001011011011101",
			1457 => "0000000100000000000101101000001000",
			1458 => "0000001001000000001100100000000100",
			1459 => "00000000000000000001011011011101",
			1460 => "00000000010101010001011011011101",
			1461 => "00000000000000000001011011011101",
			1462 => "00000000000000000001011011011101",
			1463 => "0000000001000000000000011000011100",
			1464 => "0000001101000000000110100100001100",
			1465 => "0000000011000000000011111100001000",
			1466 => "0000001011000000001010111100000100",
			1467 => "11111111010101000001011100100001",
			1468 => "00000000000000000001011100100001",
			1469 => "00000000000000000001011100100001",
			1470 => "0000000010000000001010001000001000",
			1471 => "0000001001000000001100100000000100",
			1472 => "11111111111111110001011100100001",
			1473 => "00000000000000000001011100100001",
			1474 => "0000000000000000000001000000000100",
			1475 => "00000000111111100001011100100001",
			1476 => "00000000000000000001011100100001",
			1477 => "0000000000000000001010001100000100",
			1478 => "11111110100011000001011100100001",
			1479 => "00000000000000000001011100100001",
			1480 => "0000000100000000000010010000000100",
			1481 => "11111110101010000001011101011101",
			1482 => "0000001100000000000100001000001100",
			1483 => "0000000011000000000011111100001000",
			1484 => "0000000111000000001110110000000100",
			1485 => "11111111100110010001011101011101",
			1486 => "00000000000000000001011101011101",
			1487 => "00000000000000000001011101011101",
			1488 => "0000000001000000000010001100001100",
			1489 => "0000000010000000000011001000000100",
			1490 => "00000000000000000001011101011101",
			1491 => "0000000100000000000011100100000100",
			1492 => "00000000110000010001011101011101",
			1493 => "00000000000000000001011101011101",
			1494 => "00000000000000000001011101011101",
			1495 => "0000000111000000001110001100001000",
			1496 => "0000001100000000000110000100000100",
			1497 => "11111110101001110001011110011001",
			1498 => "00000000000000000001011110011001",
			1499 => "0000000001000000000010001100010100",
			1500 => "0000000000000000000110100000000100",
			1501 => "00000000110011110001011110011001",
			1502 => "0000000110000000001100011000000100",
			1503 => "11111111110101010001011110011001",
			1504 => "0000000110000000001011001100001000",
			1505 => "0000001100000000001110001100000100",
			1506 => "00000000000000000001011110011001",
			1507 => "00000000001111100001011110011001",
			1508 => "00000000000000000001011110011001",
			1509 => "11111111101110100001011110011001",
			1510 => "0000000100000000000010010000000100",
			1511 => "11111110011111100001011111001101",
			1512 => "0000000110000000001001100100010100",
			1513 => "0000000010000000000101110000000100",
			1514 => "11111111100010010001011111001101",
			1515 => "0000000000000000000111100000001100",
			1516 => "0000000111000000000110000100000100",
			1517 => "00000000000000000001011111001101",
			1518 => "0000000001000000001110100000000100",
			1519 => "00000001001111110001011111001101",
			1520 => "00000000000000000001011111001101",
			1521 => "00000000000000000001011111001101",
			1522 => "11111111001100110001011111001101",
			1523 => "0000000100000000001101001100010000",
			1524 => "0000000100000000001011100100000100",
			1525 => "11111110011011010001100000101001",
			1526 => "0000000111000000000001111100000100",
			1527 => "11111110100111000001100000101001",
			1528 => "0000001001000000000111100100000100",
			1529 => "00000001000001010001100000101001",
			1530 => "11111111010100100001100000101001",
			1531 => "0000001111000000000111001000011000",
			1532 => "0000000110000000001100011000001000",
			1533 => "0000001001000000001100100000000100",
			1534 => "11111110100011000001100000101001",
			1535 => "00000000000000000001100000101001",
			1536 => "0000000110000000001101011000001000",
			1537 => "0000001111000000000000001100000100",
			1538 => "00000000000000000001100000101001",
			1539 => "00000001001011100001100000101001",
			1540 => "0000000111000000000111001000000100",
			1541 => "11111111010110010001100000101001",
			1542 => "00000000000000000001100000101001",
			1543 => "0000001001000000001100100000000100",
			1544 => "00000000000000000001100000101001",
			1545 => "00000001011011110001100000101001",
			1546 => "0000000100000000001111111100011000",
			1547 => "0000000100000000000010010000000100",
			1548 => "11111110011001110001100010000101",
			1549 => "0000001010000000001100000100001100",
			1550 => "0000001100000000000110000100000100",
			1551 => "11111110110100110001100010000101",
			1552 => "0000001111000000001111010000000100",
			1553 => "00000010001001100001100010000101",
			1554 => "11111111100111110001100010000101",
			1555 => "0000000100000000001101100100000100",
			1556 => "11111110100110000001100010000101",
			1557 => "11111111111110010001100010000101",
			1558 => "0000001111000000001101111000000100",
			1559 => "11111110101111100001100010000101",
			1560 => "0000000000000000000111100000001000",
			1561 => "0000001011000000001110001100000100",
			1562 => "00000000000000000001100010000101",
			1563 => "00000001100110000001100010000101",
			1564 => "0000000110000000001100011000000100",
			1565 => "11111110011001100001100010000101",
			1566 => "0000001010000000000010111100000100",
			1567 => "00000001011110110001100010000101",
			1568 => "11111111010010100001100010000101",
			1569 => "0000000100000000000010100000011100",
			1570 => "0000000100000000001111111100010100",
			1571 => "0000000100000000000100100100001000",
			1572 => "0000000001000000000110000000000100",
			1573 => "11010011100100010001100011111001",
			1574 => "11010011011101110001100011111001",
			1575 => "0000000101000000001000011000000100",
			1576 => "11010011011110000001100011111001",
			1577 => "0000000001000000001101101000000100",
			1578 => "11101011011011110001100011111001",
			1579 => "11010011100001010001100011111001",
			1580 => "0000000010000000000011001000000100",
			1581 => "11010011100010110001100011111001",
			1582 => "11101010110100000001100011111001",
			1583 => "0000001111000000000000001100001100",
			1584 => "0000000000000000001101000100001000",
			1585 => "0000000010000000000101110000000100",
			1586 => "11010011101010010001100011111001",
			1587 => "11100101111000100001100011111001",
			1588 => "11010011011110010001100011111001",
			1589 => "0000000000000000001111010000010000",
			1590 => "0000001111000000000100001000001000",
			1591 => "0000000000000000000111100000000100",
			1592 => "11101010001101010001100011111001",
			1593 => "11010101101011000001100011111001",
			1594 => "0000000101000000001001001000000100",
			1595 => "11100010100101100001100011111001",
			1596 => "11101100010011100001100011111001",
			1597 => "11010011101011100001100011111001",
			1598 => "0000000000000000001010001100010000",
			1599 => "0000000100000000000010010000000100",
			1600 => "11111110011010000001100101011101",
			1601 => "0000000111000000001110001100000100",
			1602 => "11111110100100010001100101011101",
			1603 => "0000000001000000000010001100000100",
			1604 => "00000001110000110001100101011101",
			1605 => "11111110101001010001100101011101",
			1606 => "0000001001000000001100100000010000",
			1607 => "0000000110000000001100011000000100",
			1608 => "11111110100011100001100101011101",
			1609 => "0000000000000000001111010000001000",
			1610 => "0000000011000000001111000100000100",
			1611 => "00000000000000000001100101011101",
			1612 => "00000001010111010001100101011101",
			1613 => "11111111010001110001100101011101",
			1614 => "0000001010000000000010111100010000",
			1615 => "0000000100000000001111111100000100",
			1616 => "00000000000000000001100101011101",
			1617 => "0000000000000000000101001000001000",
			1618 => "0000000011000000001111000100000100",
			1619 => "00000000000000000001100101011101",
			1620 => "00000001100101110001100101011101",
			1621 => "00000000000000000001100101011101",
			1622 => "11111111011001100001100101011101",
			1623 => "0000000100000000001111111100010000",
			1624 => "0000000001000000000110000000001100",
			1625 => "0000000111000000000001111100000100",
			1626 => "11111110011000000001100110111001",
			1627 => "0000000000000000001000000000000100",
			1628 => "00000110011001100001100110111001",
			1629 => "00000001110111010001100110111001",
			1630 => "11111110010111100001100110111001",
			1631 => "0000000011000000001111000100000100",
			1632 => "11111110011001010001100110111001",
			1633 => "0000000100000000000011100100010100",
			1634 => "0000001111000000000000001100001000",
			1635 => "0000000100000000001111111000000100",
			1636 => "00000001011101110001100110111001",
			1637 => "11111110100101010001100110111001",
			1638 => "0000000001000000001110011100000100",
			1639 => "00000001010110010001100110111001",
			1640 => "0000000010000000001000101000000100",
			1641 => "00000010000101110001100110111001",
			1642 => "00000001011001110001100110111001",
			1643 => "0000000110000000001100011000000100",
			1644 => "11111101110101010001100110111001",
			1645 => "00000000011110010001100110111001",
			1646 => "0000000100000000001111111100011000",
			1647 => "0000000001000000000000011000010100",
			1648 => "0000000001000000001100100000001000",
			1649 => "0000001010000000001111001000000100",
			1650 => "11111111010001010001101000101101",
			1651 => "00000000000000000001101000101101",
			1652 => "0000001000000000000001110100000100",
			1653 => "00000000000000000001101000101101",
			1654 => "0000001010000000000110011100000100",
			1655 => "00000000010001010001101000101101",
			1656 => "00000000000000000001101000101101",
			1657 => "11111110011010000001101000101101",
			1658 => "0000000010000000000011001000010000",
			1659 => "0000000000000000001101000100001100",
			1660 => "0000001010000000000001110100001000",
			1661 => "0000001010000000000111000100000100",
			1662 => "11111111100110010001101000101101",
			1663 => "00000000000000000001101000101101",
			1664 => "00000000100100010001101000101101",
			1665 => "11111110100100100001101000101101",
			1666 => "0000000100000000000101101000001000",
			1667 => "0000000110000000001101011000000100",
			1668 => "00000001100011110001101000101101",
			1669 => "00000000000000000001101000101101",
			1670 => "0000000110000000001100011000000100",
			1671 => "11111111011000000001101000101101",
			1672 => "0000000010000000000110010000000100",
			1673 => "00000000000000000001101000101101",
			1674 => "00000000101101110001101000101101",
			1675 => "0000001001000000000000011000100000",
			1676 => "0000001111000000000000001100001000",
			1677 => "0000000001000000001110011100000100",
			1678 => "11111111001011000001101010001001",
			1679 => "00000000000000000001101010001001",
			1680 => "0000000011000000001111000100000100",
			1681 => "00000000000000000001101010001001",
			1682 => "0000001001000000001100100000000100",
			1683 => "00000000000000000001101010001001",
			1684 => "0000001011000000001000000000001100",
			1685 => "0000000000000000000101001000001000",
			1686 => "0000001010000000000010111100000100",
			1687 => "00000001010010110001101010001001",
			1688 => "00000000000000000001101010001001",
			1689 => "00000000000000000001101010001001",
			1690 => "00000000000000000001101010001001",
			1691 => "0000000000000000000110110100001100",
			1692 => "0000000110000000001110010100000100",
			1693 => "00000000000000000001101010001001",
			1694 => "0000000001000000001100100000000100",
			1695 => "00000000000000000001101010001001",
			1696 => "11111110011111000001101010001001",
			1697 => "00000000000000000001101010001001",
			1698 => "0000000100000000001111111100010100",
			1699 => "0000000001000000000000011000001000",
			1700 => "0000000101000000001000011000000100",
			1701 => "11111110011000000001101011101101",
			1702 => "00000011101011000001101011101101",
			1703 => "0000000001000000000110000000001000",
			1704 => "0000000001000000000110000000000100",
			1705 => "11111110011001000001101011101101",
			1706 => "11111110110111100001101011101101",
			1707 => "11111110010111000001101011101101",
			1708 => "0000000011000000001111000100000100",
			1709 => "11111110011000100001101011101101",
			1710 => "0000000100000000000011100100010100",
			1711 => "0000001111000000001101111000000100",
			1712 => "11111110101101100001101011101101",
			1713 => "0000001001000000001100100000000100",
			1714 => "00000000011101000001101011101101",
			1715 => "0000001111000000000000001100000100",
			1716 => "00000001010101100001101011101101",
			1717 => "0000001111000000000100001000000100",
			1718 => "00000010100101010001101011101101",
			1719 => "00000010001101010001101011101101",
			1720 => "0000000110000000001100011000000100",
			1721 => "11111101101011010001101011101101",
			1722 => "00000000100011000001101011101101",
			1723 => "0000000000000000001010001100010100",
			1724 => "0000001001000000001100110100001000",
			1725 => "0000000101000000000100011000000100",
			1726 => "11111110011100100001101101010001",
			1727 => "00000010000001000001101101010001",
			1728 => "0000000000000000000110000100000100",
			1729 => "11111110011001010001101101010001",
			1730 => "0000001111000000000100010000000100",
			1731 => "00000010010101010001101101010001",
			1732 => "11111110011110000001101101010001",
			1733 => "0000000011000000001111000100000100",
			1734 => "11111110100001100001101101010001",
			1735 => "0000000110000000001000010000011000",
			1736 => "0000001001000000001100100000010000",
			1737 => "0000000110000000001100011000001000",
			1738 => "0000000110000000001100011000000100",
			1739 => "11111101111110100001101101010001",
			1740 => "00000000000000000001101101010001",
			1741 => "0000001010000000000010111100000100",
			1742 => "00000001101001100001101101010001",
			1743 => "00000000000000000001101101010001",
			1744 => "0000001000000000001101111000000100",
			1745 => "00000001101001010001101101010001",
			1746 => "00000000010001000001101101010001",
			1747 => "11111101110001010001101101010001",
			1748 => "0000000100000000001111111100010000",
			1749 => "0000000001000000000110000000001100",
			1750 => "0000000101000000000100011000000100",
			1751 => "11111110011010010001101110101101",
			1752 => "0000001110000000001111000100000100",
			1753 => "00000001011101010001101110101101",
			1754 => "00000011001101000001101110101101",
			1755 => "11111110011000110001101110101101",
			1756 => "0000000011000000001111000100000100",
			1757 => "11111110011011010001101110101101",
			1758 => "0000001001000000001100100000001000",
			1759 => "0000000110000000001100011000000100",
			1760 => "11111110100101110001101110101101",
			1761 => "00000000111110010001101110101101",
			1762 => "0000000100000000000011100100010000",
			1763 => "0000001111000000001101111000000100",
			1764 => "11111111001110100001101110101101",
			1765 => "0000000100000000000101101000000100",
			1766 => "00000001101100110001101110101101",
			1767 => "0000001111000000001010111000000100",
			1768 => "11111111110101110001101110101101",
			1769 => "00000001100100100001101110101101",
			1770 => "11111111111111110001101110101101",
			1771 => "0000000100000000001111111100100000",
			1772 => "0000001001000000001110100000011100",
			1773 => "0000001001000000000000011000001000",
			1774 => "0000001001000000000000011000000100",
			1775 => "11111110101110110001110000101001",
			1776 => "00000000000000000001110000101001",
			1777 => "0000000001000000001100100000001000",
			1778 => "0000000000000000001100001000000100",
			1779 => "00000001100110010001110000101001",
			1780 => "00000000000000000001110000101001",
			1781 => "0000000100000000001110001000001000",
			1782 => "0000000001000000000000011000000100",
			1783 => "11111111001111010001110000101001",
			1784 => "00000000000000000001110000101001",
			1785 => "00000000100101010001110000101001",
			1786 => "11111110011001100001110000101001",
			1787 => "0000000011000000000010011000001100",
			1788 => "0000000000000000001100100100001000",
			1789 => "0000000011000000001111000100000100",
			1790 => "11111111010101010001110000101001",
			1791 => "00000000111010000001110000101001",
			1792 => "11111110100111010001110000101001",
			1793 => "0000000010000000001000101000010000",
			1794 => "0000000100000000000001100000001000",
			1795 => "0000000010000000001010001000000100",
			1796 => "00000000000000000001110000101001",
			1797 => "00000001100110010001110000101001",
			1798 => "0000000110000000001100011000000100",
			1799 => "11111110011011100001110000101001",
			1800 => "00000001011000100001110000101001",
			1801 => "11111111100101110001110000101001",
			1802 => "0000000000000000001010001100010000",
			1803 => "0000000001000000000000011000001100",
			1804 => "0000000101000000000100011000000100",
			1805 => "11111110011000110001110010001101",
			1806 => "0000000000000000001001001000000100",
			1807 => "00000100100000000001110010001101",
			1808 => "00000001110110110001110010001101",
			1809 => "11111110011000000001110010001101",
			1810 => "0000000011000000001111000100000100",
			1811 => "11111110011000100001110010001101",
			1812 => "0000000110000000001001100100011000",
			1813 => "0000001001000000001100100000001000",
			1814 => "0000000110000000001100011000000100",
			1815 => "11111110010100010001110010001101",
			1816 => "00000001011111000001110010001101",
			1817 => "0000000000000000001111010000001100",
			1818 => "0000000010000000000100101000000100",
			1819 => "11111111101001000001110010001101",
			1820 => "0000000000000000000101001000000100",
			1821 => "00000001111111010001110010001101",
			1822 => "00000001011010100001110010001101",
			1823 => "11111110110101010001110010001101",
			1824 => "0000001000000000001100110000000100",
			1825 => "11111110010101010001110010001101",
			1826 => "00000000000000000001110010001101",
			1827 => "0000000100000000001111111100010000",
			1828 => "0000000001000000000110000000001100",
			1829 => "0000000101000000001000011000000100",
			1830 => "11111110011001010001110011110001",
			1831 => "0000000100000000001111110000000100",
			1832 => "00000011111000000001110011110001",
			1833 => "00000001100111000001110011110001",
			1834 => "11111110011000100001110011110001",
			1835 => "0000000011000000001111000100000100",
			1836 => "11111110011010010001110011110001",
			1837 => "0000001001000000001100100000001000",
			1838 => "0000001100000000001010111100000100",
			1839 => "11111110010111110001110011110001",
			1840 => "00000000000000000001110011110001",
			1841 => "0000001010000000000010111100010100",
			1842 => "0000000100000000000001100000001100",
			1843 => "0000000010000000000111111100000100",
			1844 => "00000000101011110001110011110001",
			1845 => "0000000010000000001000101000000100",
			1846 => "00000001110011110001110011110001",
			1847 => "00000000101100010001110011110001",
			1848 => "0000000110000000001100011000000100",
			1849 => "11111110000000010001110011110001",
			1850 => "00000001110101000001110011110001",
			1851 => "11111110101010010001110011110001",
			1852 => "0000000100000000000010010000000100",
			1853 => "11111110011011110001110101001101",
			1854 => "0000000010000000000101110000001000",
			1855 => "0000000011000000000000111000000100",
			1856 => "11111110110011100001110101001101",
			1857 => "00000000000000000001110101001101",
			1858 => "0000000110000000001101011000011000",
			1859 => "0000000000000000001100100100001100",
			1860 => "0000000111000000000101101100000100",
			1861 => "00000000000000000001110101001101",
			1862 => "0000000001000000000010001100000100",
			1863 => "00000001100001010001110101001101",
			1864 => "00000000000000000001110101001101",
			1865 => "0000000110000000001100011000000100",
			1866 => "11111111001001010001110101001101",
			1867 => "0000000010000000001100010100000100",
			1868 => "00000000000000000001110101001101",
			1869 => "00000000111100010001110101001101",
			1870 => "0000000110000000001001100100000100",
			1871 => "00000000000000000001110101001101",
			1872 => "0000000111000000001110001100000100",
			1873 => "00000000000000000001110101001101",
			1874 => "11111111000110110001110101001101",
			1875 => "0000000100000000001111111100010000",
			1876 => "0000000001000000000110000000001100",
			1877 => "0000000101000000001000011000000100",
			1878 => "11111110011001110001110110110001",
			1879 => "0000001011000000001000000000000100",
			1880 => "00000001101010110001110110110001",
			1881 => "00000011010011100001110110110001",
			1882 => "11111110011000110001110110110001",
			1883 => "0000000011000000001111000100000100",
			1884 => "11111110011011110001110110110001",
			1885 => "0000001001000000001100100000001000",
			1886 => "0000001100000000001010111100000100",
			1887 => "11111110100010110001110110110001",
			1888 => "00000000000000000001110110110001",
			1889 => "0000001010000000000010111100010100",
			1890 => "0000001111000000001101111000000100",
			1891 => "11111111010001010001110110110001",
			1892 => "0000000100000000000001100000001000",
			1893 => "0000000010000000001000101000000100",
			1894 => "00000001101110100001110110110001",
			1895 => "00000000011100000001110110110001",
			1896 => "0000000110000000001100011000000100",
			1897 => "11111110010111010001110110110001",
			1898 => "00000001101111100001110110110001",
			1899 => "11111110110110100001110110110001",
			1900 => "0000000100000000001111111100101000",
			1901 => "0000000100000000000100100100011100",
			1902 => "0000000001000000000110000000011000",
			1903 => "0000001001000000001001111000010100",
			1904 => "0000000100000000000010010000000100",
			1905 => "11111110010101000001111000110101",
			1906 => "0000001001000000000110000000001000",
			1907 => "0000000100000000000110110000000100",
			1908 => "00000000001100010001111000110101",
			1909 => "11111110011001000001111000110101",
			1910 => "0000000100000000001011100100000100",
			1911 => "11111110100011010001111000110101",
			1912 => "00000011100111100001111000110101",
			1913 => "00000001000011010001111000110101",
			1914 => "11111110010100100001111000110101",
			1915 => "0000000101000000001000011000000100",
			1916 => "11111110010101000001111000110101",
			1917 => "0000000001000000001101101000000100",
			1918 => "00000100010111100001111000110101",
			1919 => "11111110011001000001111000110101",
			1920 => "0000001111000000001101111000000100",
			1921 => "11111110010110000001111000110101",
			1922 => "0000001001000000001100100000001000",
			1923 => "0000000110000000001100011000000100",
			1924 => "11111110001111110001111000110101",
			1925 => "00000000000000000001111000110101",
			1926 => "0000000000000000001111010000001100",
			1927 => "0000000000000000000101001000001000",
			1928 => "0000001011000000001110001100000100",
			1929 => "00000010111011100001111000110101",
			1930 => "00000100011001110001111000110101",
			1931 => "00000010111001000001111000110101",
			1932 => "11111110100111010001111000110101",
			1933 => "0000000100000000001111111100100100",
			1934 => "0000000100000000000101001100000100",
			1935 => "11111110011001000001111010111011",
			1936 => "0000001010000000001100000100001000",
			1937 => "0000000111000000001101111000000100",
			1938 => "11111110100110010001111010111011",
			1939 => "00000011011101110001111010111011",
			1940 => "0000000100000000001101100100010000",
			1941 => "0000001000000000000011010000001100",
			1942 => "0000001010000000001001101000000100",
			1943 => "11111110101110110001111010111011",
			1944 => "0000001010000000001001101000000100",
			1945 => "00000001010000010001111010111011",
			1946 => "00000000000000000001111010111011",
			1947 => "11111110011111110001111010111011",
			1948 => "0000000011000000001010000000000100",
			1949 => "11111110011111100001111010111011",
			1950 => "00000001011011000001111010111011",
			1951 => "0000000011000000001111000100000100",
			1952 => "11111110011010110001111010111011",
			1953 => "0000001010000000000010111100011000",
			1954 => "0000001111000000001101111000000100",
			1955 => "11111111000011100001111010111011",
			1956 => "0000000100000000000001100000001100",
			1957 => "0000000010000000001000101000001000",
			1958 => "0000000010000000001110010000000100",
			1959 => "00000001010000000001111010111011",
			1960 => "00000001110001000001111010111011",
			1961 => "00000000100011100001111010111011",
			1962 => "0000000110000000001100011000000100",
			1963 => "11111101010001110001111010111011",
			1964 => "00000001110000110001111010111011",
			1965 => "11111110101011010001111010111011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(638, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(1284, initial_addr_3'length));
	end generate gen_rom_1;

	gen_rom_2: if SELECT_ROM = 2 generate
		bank <= (
			0 => "00000000000000000000000000000101",
			1 => "00000000000000000000000000001001",
			2 => "00000000000000000000000000001101",
			3 => "0000001100000000001011000000000100",
			4 => "00000000000000000000000000100001",
			5 => "0000001100000000000110100100000100",
			6 => "00000000000001110000000000100001",
			7 => "00000000000000000000000000100001",
			8 => "0000001011000000000100010000001000",
			9 => "0000001011000000000000011100000100",
			10 => "00000000000000000000000000110101",
			11 => "11111111111100110000000000110101",
			12 => "00000000000000000000000000110101",
			13 => "0000001011000000001011011100000100",
			14 => "00000000000000000000000001001001",
			15 => "0000001011000000000001001000000100",
			16 => "00000000000010100000000001001001",
			17 => "00000000000000000000000001001001",
			18 => "0000000000000000001001101000001000",
			19 => "0000001100000000001010111000000100",
			20 => "00000000000000000000000001100101",
			21 => "00000000000111010000000001100101",
			22 => "0000001100000000001001110100000100",
			23 => "11111111110101000000000001100101",
			24 => "00000000000000000000000001100101",
			25 => "0000000101000000001100100100001000",
			26 => "0000000101000000000110110100000100",
			27 => "00000000000000000000000010000001",
			28 => "00000000000100100000000010000001",
			29 => "0000000101000000001111010000000100",
			30 => "11111111111101000000000010000001",
			31 => "00000000000000000000000010000001",
			32 => "0000001011000000001011011100000100",
			33 => "00000000000000000000000010011101",
			34 => "0000000010000000001100000000001000",
			35 => "0000000010000000000010000000000100",
			36 => "00000000000000000000000010011101",
			37 => "00000000001010110000000010011101",
			38 => "00000000000000000000000010011101",
			39 => "0000000010000000001100010000001100",
			40 => "0000000000000000001100000100001000",
			41 => "0000000010000000001101000100000100",
			42 => "00000000000000000000000011000001",
			43 => "00000000001010000000000011000001",
			44 => "00000000000000000000000011000001",
			45 => "0000000010000000001010000100000100",
			46 => "11111111111100010000000011000001",
			47 => "00000000000000000000000011000001",
			48 => "0000000000000000001001101000001100",
			49 => "0000000010000000001101000100000100",
			50 => "00000000000000000000000011100101",
			51 => "0000000010000000001010000100000100",
			52 => "00000000000011000000000011100101",
			53 => "00000000000000000000000011100101",
			54 => "0000000010000000001000101000000100",
			55 => "11111111111110000000000011100101",
			56 => "00000000000000000000000011100101",
			57 => "0000000000000000001100000100001100",
			58 => "0000000010000000001100000000001000",
			59 => "0000000010000000001101000100000100",
			60 => "00000000000000000000000100010001",
			61 => "00000000000110110000000100010001",
			62 => "00000000000000000000000100010001",
			63 => "0000000010000000001000001100000100",
			64 => "11111111110111100000000100010001",
			65 => "0000000010000000001101101100000100",
			66 => "00000000000001010000000100010001",
			67 => "00000000000000000000000100010001",
			68 => "0000000000000000000001110100010000",
			69 => "0000001001000000001111000000000100",
			70 => "00000000000000000000000100110101",
			71 => "0000000100000000001110000000001000",
			72 => "0000000100000000000111011000000100",
			73 => "00000000000000000000000100110101",
			74 => "00000000000100000000000100110101",
			75 => "00000000000000000000000100110101",
			76 => "00000000000000000000000100110101",
			77 => "0000000100000000001101101100010000",
			78 => "0000000111000000000110100100000100",
			79 => "00000000000000000000000101100001",
			80 => "0000000100000000000111011000000100",
			81 => "00000000000000000000000101100001",
			82 => "0000001100000000000100011000000100",
			83 => "00000000000000000000000101100001",
			84 => "00000000001111100000000101100001",
			85 => "0000001100000000001001110100000100",
			86 => "11111111110101110000000101100001",
			87 => "00000000000000000000000101100001",
			88 => "0000000110000000001101111100001000",
			89 => "0000001100000000000100011000000100",
			90 => "00000000000000000000000110001101",
			91 => "00000000010011100000000110001101",
			92 => "0000001100000000001001110100001100",
			93 => "0000000100000000001010000100000100",
			94 => "00000000000000000000000110001101",
			95 => "0000000110000000001011001100000100",
			96 => "11111111110100010000000110001101",
			97 => "00000000000000000000000110001101",
			98 => "00000000000000000000000110001101",
			99 => "0000000000000000001100000100001000",
			100 => "0000001011000000001001110100000100",
			101 => "00000000000000000000000111000001",
			102 => "00000000000010010000000111000001",
			103 => "0000001011000000000101100100001000",
			104 => "0000001011000000000000011100000100",
			105 => "00000000000000000000000111000001",
			106 => "11111111110001100000000111000001",
			107 => "0000001011000000000101110100001000",
			108 => "0000001011000000001011011100000100",
			109 => "00000000000000000000000111000001",
			110 => "00000000000111110000000111000001",
			111 => "00000000000000000000000111000001",
			112 => "0000000000000000001100000100001000",
			113 => "0000001011000000001001110100000100",
			114 => "00000000000000000000000111111101",
			115 => "00000000000010010000000111111101",
			116 => "0000001011000000000101100100001000",
			117 => "0000001011000000000000011100000100",
			118 => "00000000000000000000000111111101",
			119 => "11111111101111010000000111111101",
			120 => "0000001011000000000101110100001000",
			121 => "0000001011000000001011011100000100",
			122 => "00000000000000000000000111111101",
			123 => "00000000001000100000000111111101",
			124 => "0000001011000000001011110100000100",
			125 => "11111111111111010000000111111101",
			126 => "00000000000000000000000111111101",
			127 => "0000001011000000001011011100001000",
			128 => "0000001001000000000111101100000100",
			129 => "11111111111010000000001000110001",
			130 => "00000000000000000000001000110001",
			131 => "0000000111000000000110100100000100",
			132 => "00000000000000000000001000110001",
			133 => "0000000111000000001000011000001100",
			134 => "0000001001000000001111000000000100",
			135 => "00000000000000000000001000110001",
			136 => "0000001001000000000010101100000100",
			137 => "00000000010111000000001000110001",
			138 => "00000000000000000000001000110001",
			139 => "00000000000000000000001000110001",
			140 => "0000001110000000000111010100010100",
			141 => "0000001011000000000101110100010000",
			142 => "0000000100000000000110010000000100",
			143 => "00000000000000000000001001011101",
			144 => "0000000110000000001101011000001000",
			145 => "0000000111000000001111011100000100",
			146 => "11111111110110010000001001011101",
			147 => "00000000000000000000001001011101",
			148 => "00000000000000000000001001011101",
			149 => "00000000000000000000001001011101",
			150 => "00000000000000000000001001011101",
			151 => "0000000100000000000001011100010100",
			152 => "0000001000000000001000100100000100",
			153 => "00000000000000000000001010011001",
			154 => "0000001100000000000100011000000100",
			155 => "00000000000000000000001010011001",
			156 => "0000001100000000000001101000001000",
			157 => "0000000000000000001111001000000100",
			158 => "00000000010011010000001010011001",
			159 => "00000000000000000000001010011001",
			160 => "00000000000000000000001010011001",
			161 => "0000000001000000001100011000001000",
			162 => "0000001100000000001011011100000100",
			163 => "11111111110111000000001010011001",
			164 => "00000000000000000000001010011001",
			165 => "00000000000000000000001010011001",
			166 => "0000001110000000001100000000010000",
			167 => "0000000100000000001100010000000100",
			168 => "00000000000000000000001011011101",
			169 => "0000001010000000000000001000000100",
			170 => "11111111110000010000001011011101",
			171 => "0000001010000000001010100000000100",
			172 => "00000000000001000000001011011101",
			173 => "11111111111011110000001011011101",
			174 => "0000000100000000000001011100010000",
			175 => "0000000001000000001101111100001100",
			176 => "0000000011000000001000100000001000",
			177 => "0000000011000000001010000100000100",
			178 => "00000000000000000000001011011101",
			179 => "00000000100101000000001011011101",
			180 => "00000000000000000000001011011101",
			181 => "00000000000000000000001011011101",
			182 => "00000000000000000000001011011101",
			183 => "0000000100000000001101101100011100",
			184 => "0000001110000000000111011000010100",
			185 => "0000000000000000001100000100001100",
			186 => "0000000000000000000001010100000100",
			187 => "00000000000000000000001100110001",
			188 => "0000000001000000001001011000000100",
			189 => "00000000000000000000001100110001",
			190 => "00000000010000010000001100110001",
			191 => "0000001011000000000101100100000100",
			192 => "11111111101011010000001100110001",
			193 => "00000000000000000000001100110001",
			194 => "0000000011000000001010000100000100",
			195 => "00000000000000000000001100110001",
			196 => "00000000110001100000001100110001",
			197 => "0000001001000000001010100000001100",
			198 => "0000000111000000000101110100001000",
			199 => "0000001000000000000001010000000100",
			200 => "00000000000000000000001100110001",
			201 => "11111111101010100000001100110001",
			202 => "00000000000000000000001100110001",
			203 => "00000000000000000000001100110001",
			204 => "0000000100000000000001011100011000",
			205 => "0000001001000000000100111100000100",
			206 => "00000000000000000000001101101101",
			207 => "0000000001000000001101111100010000",
			208 => "0000000111000000000110100100000100",
			209 => "00000000000000000000001101101101",
			210 => "0000000000000000001111001000001000",
			211 => "0000001011000000000100000100000100",
			212 => "00000000000000000000001101101101",
			213 => "00000000100010100000001101101101",
			214 => "00000000000000000000001101101101",
			215 => "00000000000000000000001101101101",
			216 => "0000000110000000000100111100000100",
			217 => "11111111111101000000001101101101",
			218 => "00000000000000000000001101101101",
			219 => "0000001110000000001100000000001000",
			220 => "0000001101000000001001010100000100",
			221 => "00000000000000000000001110101001",
			222 => "11111111111110100000001110101001",
			223 => "0000001101000000000011001000010100",
			224 => "0000001001000000000100111100000100",
			225 => "00000000000000000000001110101001",
			226 => "0000001110000000000010010100001100",
			227 => "0000001101000000001110000100000100",
			228 => "00000000000000000000001110101001",
			229 => "0000001001000000000010101100000100",
			230 => "00000000001100000000001110101001",
			231 => "00000000000000000000001110101001",
			232 => "00000000000000000000001110101001",
			233 => "00000000000000000000001110101001",
			234 => "0000000001000000000000111100001000",
			235 => "0000001000000000000100101100000100",
			236 => "00000000000000000000001111100101",
			237 => "11111111111000010000001111100101",
			238 => "0000001111000000001011110000010100",
			239 => "0000001110000000001100010000000100",
			240 => "00000000000000000000001111100101",
			241 => "0000001001000000000100111100000100",
			242 => "00000000000000000000001111100101",
			243 => "0000000001000000001100011000001000",
			244 => "0000001000000000000001110000000100",
			245 => "00000000001110110000001111100101",
			246 => "00000000000000000000001111100101",
			247 => "00000000000000000000001111100101",
			248 => "00000000000000000000001111100101",
			249 => "0000000100000000001101101100011000",
			250 => "0000000001000000001001011000000100",
			251 => "00000000000000000000010000101001",
			252 => "0000000011000000001000100000010000",
			253 => "0000000000000000001111001000001100",
			254 => "0000001111000000000010000100000100",
			255 => "00000000000000000000010000101001",
			256 => "0000000011000000000010000100000100",
			257 => "00000000000000000000010000101001",
			258 => "00000000001100100000010000101001",
			259 => "00000000000000000000010000101001",
			260 => "00000000000000000000010000101001",
			261 => "0000000001000000000001111000001000",
			262 => "0000000011000000001111101000000100",
			263 => "11111111111101110000010000101001",
			264 => "00000000000000000000010000101001",
			265 => "00000000000000000000010000101001",
			266 => "0000001100000000001010111000000100",
			267 => "00000000000000000000010001011101",
			268 => "0000000101000000001111010000010100",
			269 => "0000000000000000000001110100010000",
			270 => "0000001101000000001010001000001100",
			271 => "0000001101000000001110000100000100",
			272 => "00000000000000000000010001011101",
			273 => "0000000111000000001111011100000100",
			274 => "00000000010010110000010001011101",
			275 => "00000000000000000000010001011101",
			276 => "00000000000000000000010001011101",
			277 => "00000000000000000000010001011101",
			278 => "00000000000000000000010001011101",
			279 => "0000001100000000001001110100011000",
			280 => "0000000100000000001100010000000100",
			281 => "00000000000000000000010010010001",
			282 => "0000001001000000000111101100010000",
			283 => "0000001100000000001010111000000100",
			284 => "00000000000000000000010010010001",
			285 => "0000000111000000001001001000000100",
			286 => "00000000000000000000010010010001",
			287 => "0000000001000000000001111000000100",
			288 => "11111111101001100000010010010001",
			289 => "00000000000000000000010010010001",
			290 => "00000000000000000000010010010001",
			291 => "00000000000000000000010010010001",
			292 => "0000000100000000001011101100010000",
			293 => "0000001010000000000000001000000100",
			294 => "00000000000000000000010011100101",
			295 => "0000001101000000000101001000000100",
			296 => "00000000000000000000010011100101",
			297 => "0000000011000000001111100100000100",
			298 => "00000000010001010000010011100101",
			299 => "00000000000000000000010011100101",
			300 => "0000001001000000000111101100001000",
			301 => "0000001100000000001001110100000100",
			302 => "11111111100001010000010011100101",
			303 => "00000000000000000000010011100101",
			304 => "0000001100000000000110100100010000",
			305 => "0000001110000000000111010100000100",
			306 => "00000000000000000000010011100101",
			307 => "0000000001000000001010011000001000",
			308 => "0000000000000000001010101100000100",
			309 => "00000000010100110000010011100101",
			310 => "00000000000000000000010011100101",
			311 => "00000000000000000000010011100101",
			312 => "00000000000000000000010011100101",
			313 => "0000000000000000001100000100001100",
			314 => "0000001000000000001000100100000100",
			315 => "00000000000000000000010101000001",
			316 => "0000001001000000001111000000000100",
			317 => "00000000000000000000010101000001",
			318 => "00000000000101000000010101000001",
			319 => "0000000110000000000100111100010000",
			320 => "0000001011000000001011110100001100",
			321 => "0000000010000000000111011000000100",
			322 => "00000000000000000000010101000001",
			323 => "0000001000000000001000010100000100",
			324 => "00000000000000000000010101000001",
			325 => "11111111011011010000010101000001",
			326 => "00000000000000000000010101000001",
			327 => "0000000000000000001010101100010000",
			328 => "0000001001000000001010100000000100",
			329 => "00000000000000000000010101000001",
			330 => "0000001001000000000011101000001000",
			331 => "0000001011000000000001001000000100",
			332 => "00000000001110110000010101000001",
			333 => "00000000000000000000010101000001",
			334 => "00000000000000000000010101000001",
			335 => "00000000000000000000010101000001",
			336 => "0000000110000000001001100100011000",
			337 => "0000001011000000001011110100010100",
			338 => "0000000010000000001010000100001100",
			339 => "0000001110000000001100000000001000",
			340 => "0000001110000000001110010000000100",
			341 => "00000000000000000000010110011101",
			342 => "11111111111011000000010110011101",
			343 => "00000000000000000000010110011101",
			344 => "0000001011000000000000011100000100",
			345 => "00000000000000000000010110011101",
			346 => "11111111100011000000010110011101",
			347 => "00000000000000000000010110011101",
			348 => "0000001011000000001010010100010100",
			349 => "0000001001000000000111101100000100",
			350 => "00000000000000000000010110011101",
			351 => "0000001010000000001001000100001100",
			352 => "0000001110000000001000001100000100",
			353 => "00000000000000000000010110011101",
			354 => "0000001111000000001110000000000100",
			355 => "00000000011001010000010110011101",
			356 => "00000000000000000000010110011101",
			357 => "00000000000000000000010110011101",
			358 => "00000000000000000000010110011101",
			359 => "0000001011000000001011011100010000",
			360 => "0000001110000000000111011000001000",
			361 => "0000000011000000001010000100000100",
			362 => "11111111110001000000010111110001",
			363 => "00000000000000000000010111110001",
			364 => "0000001001000000000000001000000100",
			365 => "00000000000001000000010111110001",
			366 => "00000000000000000000010111110001",
			367 => "0000000111000000000110100100000100",
			368 => "00000000000000000000010111110001",
			369 => "0000000100000000001101101100010100",
			370 => "0000000000000000000101000100000100",
			371 => "00000000000000000000010111110001",
			372 => "0000000100000000000111011000000100",
			373 => "00000000000000000000010111110001",
			374 => "0000000001000000001001011000000100",
			375 => "00000000000000000000010111110001",
			376 => "0000001111000000001100010000000100",
			377 => "00000000000000000000010111110001",
			378 => "00000000100000000000010111110001",
			379 => "00000000000000000000010111110001",
			380 => "0000000000000000000111000100011100",
			381 => "0000001100000000001010111000000100",
			382 => "00000000000000000000011000110101",
			383 => "0000001101000000001010001000010100",
			384 => "0000001101000000001110000100000100",
			385 => "00000000000000000000011000110101",
			386 => "0000001010000000000000001000000100",
			387 => "00000000000000000000011000110101",
			388 => "0000001011000000000001011000000100",
			389 => "00000000000000000000011000110101",
			390 => "0000001011000000000101110100000100",
			391 => "00000000010111010000011000110101",
			392 => "00000000000000000000011000110101",
			393 => "00000000000000000000011000110101",
			394 => "0000000110000000001000010000000100",
			395 => "11111111111101100000011000110101",
			396 => "00000000000000000000011000110101",
			397 => "0000000100000000001101101100100100",
			398 => "0000001110000000000111011000011100",
			399 => "0000000000000000001100000100010100",
			400 => "0000001000000000001000100100010000",
			401 => "0000001101000000000111111100001100",
			402 => "0000001111000000000010000000000100",
			403 => "00000000000000000000011010010001",
			404 => "0000001101000000001110000100000100",
			405 => "00000000000000000000011010010001",
			406 => "11111111110000110000011010010001",
			407 => "00000000000000000000011010010001",
			408 => "00000000010100100000011010010001",
			409 => "0000001011000000000101100100000100",
			410 => "11111111100111110000011010010001",
			411 => "00000000000000000000011010010001",
			412 => "0000000011000000001010000100000100",
			413 => "00000000000000000000011010010001",
			414 => "00000000110111110000011010010001",
			415 => "0000000110000000000100111100001000",
			416 => "0000001100000000001111011100000100",
			417 => "11111111100111100000011010010001",
			418 => "00000000000000000000011010010001",
			419 => "00000000000000000000011010010001",
			420 => "0000000101000000001111010000100100",
			421 => "0000000101000000001101000100001100",
			422 => "0000000000000000000001010100000100",
			423 => "00000000000000000000011011110101",
			424 => "0000000010000000001000001100000100",
			425 => "11111111101011100000011011110101",
			426 => "00000000000000000000011011110101",
			427 => "0000001100000000001001001000010100",
			428 => "0000000110000000000100110100000100",
			429 => "00000000000000000000011011110101",
			430 => "0000000010000000001101101100001100",
			431 => "0000000001000000000100110100001000",
			432 => "0000000000000000000001110100000100",
			433 => "00000000101101110000011011110101",
			434 => "00000000000000000000011011110101",
			435 => "00000000000000000000011011110101",
			436 => "00000000000000000000011011110101",
			437 => "00000000000000000000011011110101",
			438 => "0000001011000000001011110100001100",
			439 => "0000001110000000000001011100001000",
			440 => "0000001011000000000010001000000100",
			441 => "00000000000000000000011011110101",
			442 => "11111111101110100000011011110101",
			443 => "00000000000000000000011011110101",
			444 => "00000000000000000000011011110101",
			445 => "0000000100000000000111010100010000",
			446 => "0000001000000000001000100100000100",
			447 => "00000000000000000000011101011001",
			448 => "0000001111000000001111010100001000",
			449 => "0000001110000000000011001000000100",
			450 => "00000000000000000000011101011001",
			451 => "00000000001100110000011101011001",
			452 => "00000000000000000000011101011001",
			453 => "0000000110000000000100111100011000",
			454 => "0000001011000000001011110100010100",
			455 => "0000000000000000001100000100000100",
			456 => "00000000000000000000011101011001",
			457 => "0000000110000000001111000000001100",
			458 => "0000001011000000000000011100000100",
			459 => "00000000000000000000011101011001",
			460 => "0000001000000000001000010100000100",
			461 => "00000000000000000000011101011001",
			462 => "11111111011010100000011101011001",
			463 => "00000000000000000000011101011001",
			464 => "00000000000000000000011101011001",
			465 => "0000000000000000001010101100001000",
			466 => "0000000001000000001010011000000100",
			467 => "00000000001000100000011101011001",
			468 => "00000000000000000000011101011001",
			469 => "00000000000000000000011101011001",
			470 => "0000000100000000001100010000000100",
			471 => "00000000000000000000011110010101",
			472 => "0000000101000000001111010000011000",
			473 => "0000001110000000000111010100010100",
			474 => "0000001011000000000100010000010000",
			475 => "0000001100000000001010111000000100",
			476 => "00000000000000000000011110010101",
			477 => "0000001011000000000000011100000100",
			478 => "00000000000000000000011110010101",
			479 => "0000000011000000000000010000000100",
			480 => "11111111011111000000011110010101",
			481 => "00000000000000000000011110010101",
			482 => "00000000000000000000011110010101",
			483 => "00000000000000000000011110010101",
			484 => "00000000000000000000011110010101",
			485 => "0000001110000000000111010100011100",
			486 => "0000001011000000000101110100011000",
			487 => "0000000101000000001100100100000100",
			488 => "00000000000000000000011111010001",
			489 => "0000000001000000001001011000000100",
			490 => "00000000000000000000011111010001",
			491 => "0000000101000000001111010000001100",
			492 => "0000001010000000000010101100001000",
			493 => "0000000111000000001111011100000100",
			494 => "11111111100111010000011111010001",
			495 => "00000000000000000000011111010001",
			496 => "00000000000000000000011111010001",
			497 => "00000000000000000000011111010001",
			498 => "00000000000000000000011111010001",
			499 => "00000000000000000000011111010001",
			500 => "0000001001000000001111000000000100",
			501 => "00000000000000000000100000001101",
			502 => "0000000000000000000111000100011000",
			503 => "0000001101000000001010001000010100",
			504 => "0000001101000000001110000100000100",
			505 => "00000000000000000000100000001101",
			506 => "0000001011000000000000011100000100",
			507 => "00000000000000000000100000001101",
			508 => "0000001010000000000000001000000100",
			509 => "00000000000000000000100000001101",
			510 => "0000001100000000001010111000000100",
			511 => "00000000000000000000100000001101",
			512 => "00000000010011100000100000001101",
			513 => "00000000000000000000100000001101",
			514 => "00000000000000000000100000001101",
			515 => "0000000000000000000010101000011100",
			516 => "0000001001000000001111000000000100",
			517 => "00000000000000000000100001001001",
			518 => "0000000111000000000110100100000100",
			519 => "00000000000000000000100001001001",
			520 => "0000000000000000000001010100000100",
			521 => "00000000000000000000100001001001",
			522 => "0000000001000000001010011000001100",
			523 => "0000001100000000001010111000000100",
			524 => "00000000000000000000100001001001",
			525 => "0000000100000000000111011000000100",
			526 => "00000000000000000000100001001001",
			527 => "00000000011000110000100001001001",
			528 => "00000000000000000000100001001001",
			529 => "00000000000000000000100001001001",
			530 => "0000000001000000000000111100010100",
			531 => "0000000010000000001100010000000100",
			532 => "00000000000000000000100010100101",
			533 => "0000001101000000000111111100000100",
			534 => "00000000000000000000100010100101",
			535 => "0000000101000000000101110000001000",
			536 => "0000001110000000001100010000000100",
			537 => "00000000000000000000100010100101",
			538 => "11111111101000010000100010100101",
			539 => "00000000000000000000100010100101",
			540 => "0000000000000000000001110100011000",
			541 => "0000001100000000000100011000000100",
			542 => "00000000000000000000100010100101",
			543 => "0000001110000000001100000000000100",
			544 => "00000000000000000000100010100101",
			545 => "0000000001000000001101111100001100",
			546 => "0000000010000000001101101100001000",
			547 => "0000000101000000000110100000000100",
			548 => "00000000000000000000100010100101",
			549 => "00000000100011110000100010100101",
			550 => "00000000000000000000100010100101",
			551 => "00000000000000000000100010100101",
			552 => "00000000000000000000100010100101",
			553 => "0000000100000000001111100100011000",
			554 => "0000001111000000001110110100000100",
			555 => "00000000000000000000100100011001",
			556 => "0000000011000000000000010000010000",
			557 => "0000001010000000001010100000000100",
			558 => "00000000000000000000100100011001",
			559 => "0000000111000000000110100100000100",
			560 => "00000000000000000000100100011001",
			561 => "0000001010000000000011101000000100",
			562 => "00000000101010010000100100011001",
			563 => "00000000000000000000100100011001",
			564 => "00000000000000000000100100011001",
			565 => "0000000011000000001111100100010000",
			566 => "0000001100000000001010111000000100",
			567 => "00000000000000000000100100011001",
			568 => "0000000101000000000010110100000100",
			569 => "00000000000000000000100100011001",
			570 => "0000000101000000000111100000000100",
			571 => "11111111100010010000100100011001",
			572 => "00000000000000000000100100011001",
			573 => "0000000001000000001110010100000100",
			574 => "00000000000000000000100100011001",
			575 => "0000000010000000001011110000001100",
			576 => "0000000001000000001010011000001000",
			577 => "0000001111000000001011110000000100",
			578 => "00000000001000110000100100011001",
			579 => "00000000000000000000100100011001",
			580 => "00000000000000000000100100011001",
			581 => "00000000000000000000100100011001",
			582 => "0000001011000000001011011100010000",
			583 => "0000000100000000001010000100000100",
			584 => "00000000000000000000100110010101",
			585 => "0000001110000000000111010100001000",
			586 => "0000000101000000000111100000000100",
			587 => "11111111011011000000100110010101",
			588 => "00000000000000000000100110010101",
			589 => "00000000000000000000100110010101",
			590 => "0000000110000000000100110100010000",
			591 => "0000001011000000000010001000000100",
			592 => "00000000000000000000100110010101",
			593 => "0000000101000000001001010000001000",
			594 => "0000001100000000001011000000000100",
			595 => "00000000000000000000100110010101",
			596 => "11111111011010000000100110010101",
			597 => "00000000000000000000100110010101",
			598 => "0000000100000000000001011100001000",
			599 => "0000000111000000000110100100000100",
			600 => "00000000000000000000100110010101",
			601 => "00000000110000010000100110010101",
			602 => "0000001001000000001010100000001000",
			603 => "0000001011000000000001001000000100",
			604 => "11111111011101110000100110010101",
			605 => "00000000000000000000100110010101",
			606 => "0000000001000000001010011000001100",
			607 => "0000001101000000001100010100001000",
			608 => "0000000011000000001000100000000100",
			609 => "00000000000000000000100110010101",
			610 => "00000000100000100000100110010101",
			611 => "00000000000000000000100110010101",
			612 => "00000000000000000000100110010101",
			613 => "0000001100000000001011000000101100",
			614 => "0000000100000000000110111100010000",
			615 => "0000001100000000001010111000000100",
			616 => "00000000000000000000101000011001",
			617 => "0000000111000000001000011000001000",
			618 => "0000000111000000001011000000000100",
			619 => "00000000000000000000101000011001",
			620 => "00000000001100010000101000011001",
			621 => "00000000000000000000101000011001",
			622 => "0000001001000000000111101100001100",
			623 => "0000000101000000001110101000000100",
			624 => "00000000000000000000101000011001",
			625 => "0000001110000000001100010000000100",
			626 => "00000000000000000000101000011001",
			627 => "11111111011001100000101000011001",
			628 => "0000000001000000001101111100001100",
			629 => "0000001110000000001111010100000100",
			630 => "00000000000000000000101000011001",
			631 => "0000001010000000001000100100000100",
			632 => "00000000001111110000101000011001",
			633 => "00000000000000000000101000011001",
			634 => "00000000000000000000101000011001",
			635 => "0000001011000000000100010000000100",
			636 => "00000000000000000000101000011001",
			637 => "0000000001000000001100011000010000",
			638 => "0000000111000000001000011000000100",
			639 => "00000000000000000000101000011001",
			640 => "0000001111000000001011110000001000",
			641 => "0000000000000000000111000000000100",
			642 => "00000000101110000000101000011001",
			643 => "00000000000000000000101000011001",
			644 => "00000000000000000000101000011001",
			645 => "00000000000000000000101000011001",
			646 => "0000000110000000001101111100010000",
			647 => "0000000111000000001011000000000100",
			648 => "00000000000000000000101010010101",
			649 => "0000000111000000001111011100001000",
			650 => "0000000010000000001100000000000100",
			651 => "00000000010110000000101010010101",
			652 => "00000000000000000000101010010101",
			653 => "00000000000000000000101010010101",
			654 => "0000000111000000001000011000100100",
			655 => "0000001001000000000100101100010000",
			656 => "0000000101000000001100100100000100",
			657 => "00000000000000000000101010010101",
			658 => "0000001101000000001001011100001000",
			659 => "0000001101000000000010011100000100",
			660 => "00000000000000000000101010010101",
			661 => "11111111011010000000101010010101",
			662 => "00000000000000000000101010010101",
			663 => "0000001010000000001000100100010000",
			664 => "0000001010000000000010101100000100",
			665 => "00000000000000000000101010010101",
			666 => "0000000010000000001101101100001000",
			667 => "0000000010000000000010000100000100",
			668 => "00000000000000000000101010010101",
			669 => "00000000001010010000101010010101",
			670 => "00000000000000000000101010010101",
			671 => "00000000000000000000101010010101",
			672 => "0000000011000000001000100000001000",
			673 => "0000001000000000000110011100000100",
			674 => "00000000011000000000101010010101",
			675 => "00000000000000000000101010010101",
			676 => "00000000000000000000101010010101",
			677 => "0000001100000000001001110100110000",
			678 => "0000000110000000000100111100100100",
			679 => "0000000100000000001111100100011000",
			680 => "0000000010000000000110111100010000",
			681 => "0000000010000000001110110100000100",
			682 => "00000000000000000000101100011001",
			683 => "0000001010000000000010101100001000",
			684 => "0000001111000000000010000100000100",
			685 => "00000000000000000000101100011001",
			686 => "11111111110000000000101100011001",
			687 => "00000000000000000000101100011001",
			688 => "0000000110000000001100011000000100",
			689 => "00000000000000000000101100011001",
			690 => "00000000010011100000101100011001",
			691 => "0000000111000000000110100100000100",
			692 => "00000000000000000000101100011001",
			693 => "0000000110000000001101011000000100",
			694 => "00000000000000000000101100011001",
			695 => "11111111010111010000101100011001",
			696 => "0000000000000000000010101000001000",
			697 => "0000000011000000001100111000000100",
			698 => "00000000000000000000101100011001",
			699 => "00000000010010000000101100011001",
			700 => "00000000000000000000101100011001",
			701 => "0000000010000000000010010100010000",
			702 => "0000001000000000001000100100000100",
			703 => "00000000000000000000101100011001",
			704 => "0000000111000000000101100100001000",
			705 => "0000000001000000001100011000000100",
			706 => "00000000100010110000101100011001",
			707 => "00000000000000000000101100011001",
			708 => "00000000000000000000101100011001",
			709 => "00000000000000000000101100011001",
			710 => "0000000100000000001011101100111000",
			711 => "0000001100000000001011000000100100",
			712 => "0000000111000000000110100100010000",
			713 => "0000000111000000001001001000000100",
			714 => "00000000000000000000101110110101",
			715 => "0000001010000000000010101100001000",
			716 => "0000000100000000001001100000000100",
			717 => "00000000000000000000101110110101",
			718 => "11111111100110110000101110110101",
			719 => "00000000000000000000101110110101",
			720 => "0000000110000000001101111100000100",
			721 => "00000000000000000000101110110101",
			722 => "0000000100000000001000100000001100",
			723 => "0000000101000000001111010000001000",
			724 => "0000001010000000000000001000000100",
			725 => "00000000000000000000101110110101",
			726 => "00000000110010110000101110110101",
			727 => "00000000000000000000101110110101",
			728 => "00000000000000000000101110110101",
			729 => "0000000101000000000111100000001100",
			730 => "0000001001000000000100101100001000",
			731 => "0000000100000000000010000100000100",
			732 => "00000000000000000000101110110101",
			733 => "11111111011010100000101110110101",
			734 => "00000000000000000000101110110101",
			735 => "0000000010000000001110110100000100",
			736 => "00000000000000000000101110110101",
			737 => "00000000001111110000101110110101",
			738 => "0000000110000000001001100100001100",
			739 => "0000001100000000001001110100001000",
			740 => "0000000000000000001011010100000100",
			741 => "00000000000000000000101110110101",
			742 => "11111111010101110000101110110101",
			743 => "00000000000000000000101110110101",
			744 => "0000000000000000000111000100001000",
			745 => "0000000111000000000111010000000100",
			746 => "00000000011000000000101110110101",
			747 => "00000000000000000000101110110101",
			748 => "00000000000000000000101110110101",
			749 => "0000000100000000000001011100110000",
			750 => "0000001011000000000100010000101000",
			751 => "0000001101000000000101110000010100",
			752 => "0000001101000000001110000100000100",
			753 => "00000000000000000000110000101001",
			754 => "0000001001000000001111000000000100",
			755 => "00000000000000000000110000101001",
			756 => "0000001001000000000111101100001000",
			757 => "0000001010000000000000001000000100",
			758 => "00000000000000000000110000101001",
			759 => "00000000100010000000110000101001",
			760 => "00000000000000000000110000101001",
			761 => "0000001000000000000001010000010000",
			762 => "0000001101000000000111111100001100",
			763 => "0000001001000000001111000000000100",
			764 => "00000000000000000000110000101001",
			765 => "0000000010000000000110010000000100",
			766 => "00000000000000000000110000101001",
			767 => "11111111101010010000110000101001",
			768 => "00000000000000000000110000101001",
			769 => "00000000000000000000110000101001",
			770 => "0000000011000000001000100000000100",
			771 => "00000000010111110000110000101001",
			772 => "00000000000000000000110000101001",
			773 => "0000001100000000001001110100001000",
			774 => "0000000011000000000010010100000100",
			775 => "11111111101011100000110000101001",
			776 => "00000000000000000000110000101001",
			777 => "00000000000000000000110000101001",
			778 => "0000001011000000001011011100010100",
			779 => "0000000000000000001100000100001100",
			780 => "0000001100000000001011000000001000",
			781 => "0000001100000000001101010100000100",
			782 => "00000000000000000000110011000101",
			783 => "00000000000111000000110011000101",
			784 => "00000000000000000000110011000101",
			785 => "0000001110000000000111010100000100",
			786 => "11111111100001100000110011000101",
			787 => "00000000000000000000110011000101",
			788 => "0000000110000000000100110100010100",
			789 => "0000001110000000001100010000010000",
			790 => "0000001101000000000010011100000100",
			791 => "00000000000000000000110011000101",
			792 => "0000001100000000000100011000000100",
			793 => "00000000000000000000110011000101",
			794 => "0000001110000000000010000000000100",
			795 => "00000000000000000000110011000101",
			796 => "11111111011001000000110011000101",
			797 => "00000000000000000000110011000101",
			798 => "0000000100000000000001011100001100",
			799 => "0000001001000000001111000000000100",
			800 => "00000000000000000000110011000101",
			801 => "0000000111000000000110100100000100",
			802 => "00000000000000000000110011000101",
			803 => "00000000101110000000110011000101",
			804 => "0000001001000000001010100000001100",
			805 => "0000001011000000000001001000001000",
			806 => "0000001001000000001010100000000100",
			807 => "11111111100100000000110011000101",
			808 => "00000000000000000000110011000101",
			809 => "00000000000000000000110011000101",
			810 => "0000000001000000001010011000001100",
			811 => "0000001101000000001100010100001000",
			812 => "0000000000000000001010101100000100",
			813 => "00000000011110110000110011000101",
			814 => "00000000000000000000110011000101",
			815 => "00000000000000000000110011000101",
			816 => "00000000000000000000110011000101",
			817 => "0000000000000000001001101000101100",
			818 => "0000001110000000001010000100100100",
			819 => "0000001100000000001010111000000100",
			820 => "00000000000000000000110101100001",
			821 => "0000001010000000001010100000010000",
			822 => "0000001001000000001111000000001000",
			823 => "0000000011000000001111010100000100",
			824 => "00000000010110100000110101100001",
			825 => "00000000000000000000110101100001",
			826 => "0000000010000000000010000000000100",
			827 => "00000000000000000000110101100001",
			828 => "11111111111000110000110101100001",
			829 => "0000000101000000000110100000000100",
			830 => "00000000000000000000110101100001",
			831 => "0000000111000000000110100100000100",
			832 => "00000000000000000000110101100001",
			833 => "0000000011000000001011111000000100",
			834 => "00000000111011010000110101100001",
			835 => "00000000000000000000110101100001",
			836 => "0000001100000000001001001000000100",
			837 => "11111111111001100000110101100001",
			838 => "00000000000000000000110101100001",
			839 => "0000000110000000001001100100010000",
			840 => "0000000100000000001011101100001000",
			841 => "0000000100000000000110101100000100",
			842 => "11111111111100000000110101100001",
			843 => "00000000000000000000110101100001",
			844 => "0000001100000000001001110100000100",
			845 => "11111111000010110000110101100001",
			846 => "00000000000000000000110101100001",
			847 => "0000001100000000001001110100010000",
			848 => "0000000100000000000101000000001100",
			849 => "0000001100000000000100011000000100",
			850 => "00000000000000000000110101100001",
			851 => "0000001010000000001001000100000100",
			852 => "00000000001101100000110101100001",
			853 => "00000000000000000000110101100001",
			854 => "00000000000000000000110101100001",
			855 => "00000000000000000000110101100001",
			856 => "0000000000000000001010101100101000",
			857 => "0000001100000000001101010100000100",
			858 => "11111110001011010000110110110101",
			859 => "0000000101000000001110010000100000",
			860 => "0000001110000000001101101100010100",
			861 => "0000001001000000001111000000001000",
			862 => "0000000010000000000001000000000100",
			863 => "00000001101110010000110110110101",
			864 => "11111110011000100000110110110101",
			865 => "0000000000000000000001110100001000",
			866 => "0000001100000000001001110100000100",
			867 => "00000000101000010000110110110101",
			868 => "00000001101011110000110110110101",
			869 => "11111110100000100000110110110101",
			870 => "0000000000000000001010101100001000",
			871 => "0000001000000000000001010100000100",
			872 => "00000000011000000000110110110101",
			873 => "00000010011110000000110110110101",
			874 => "00000100100010010000110110110101",
			875 => "11111110100011100000110110110101",
			876 => "11111110011001100000110110110101",
			877 => "0000000100000000001000001100100000",
			878 => "0000001100000000001010111000000100",
			879 => "00000000000000000000111001100001",
			880 => "0000000111000000001000011000001100",
			881 => "0000000001000000001011111100001000",
			882 => "0000000001000000001001011000000100",
			883 => "00000000000000000000111001100001",
			884 => "00000000111100000000111001100001",
			885 => "00000000000000000000111001100001",
			886 => "0000000000000000000001010100001000",
			887 => "0000000000000000000101000100000100",
			888 => "00000000000000000000111001100001",
			889 => "11111111101101110000111001100001",
			890 => "0000000000000000000001010100000100",
			891 => "00000000000000000000111001100001",
			892 => "00000000010001100000111001100001",
			893 => "0000000011000000001010000100010000",
			894 => "0000001100000000001011000000001100",
			895 => "0000000111000000000001101000001000",
			896 => "0000001110000000001111010100000100",
			897 => "11111110111001110000111001100001",
			898 => "00000000000000000000111001100001",
			899 => "00000000000000000000111001100001",
			900 => "00000000000000000000111001100001",
			901 => "0000000010000000001000001100001000",
			902 => "0000000001000000000000111100000100",
			903 => "00000000000000000000111001100001",
			904 => "00000000111001000000111001100001",
			905 => "0000001110000000000111010100001100",
			906 => "0000001100000000001011000000001000",
			907 => "0000000111000000000110100100000100",
			908 => "00000000000000000000111001100001",
			909 => "11111111000100000000111001100001",
			910 => "00000000000000000000111001100001",
			911 => "0000000010000000001011111000000100",
			912 => "00000000100110110000111001100001",
			913 => "0000000001000000000001111000001000",
			914 => "0000000111000000000001011000000100",
			915 => "11111111010110110000111001100001",
			916 => "00000000000000000000111001100001",
			917 => "0000000001000000000100110100000100",
			918 => "00000000010000100000111001100001",
			919 => "11111111110001000000111001100001",
			920 => "0000000000000000001010101100101000",
			921 => "0000001100000000001101010100000100",
			922 => "11111110001011100000111010110101",
			923 => "0000001101000000001001100000100000",
			924 => "0000001110000000001101101100011000",
			925 => "0000001001000000001111000000001000",
			926 => "0000001010000000001001111100000100",
			927 => "00000001111100000000111010110101",
			928 => "11111110010111000000111010110101",
			929 => "0000001100000000001001110100001000",
			930 => "0000001101000000001110010000000100",
			931 => "00000000110000000000111010110101",
			932 => "11111110111111100000111010110101",
			933 => "0000000001000000000100110100000100",
			934 => "00000001110000010000111010110101",
			935 => "11111111100011110000111010110101",
			936 => "0000000000000000001010101100000100",
			937 => "00000010011011010000111010110101",
			938 => "00000100111001100000111010110101",
			939 => "11111110011110010000111010110101",
			940 => "11111110011001100000111010110101",
			941 => "0000000100000000001011110000111100",
			942 => "0000001001000000001111000000010000",
			943 => "0000001011000000000010001000001100",
			944 => "0000000110000000000000111100001000",
			945 => "0000001000000000001001111100000100",
			946 => "11111110011111100000111101010001",
			947 => "00000001111011110000111101010001",
			948 => "11111110011000010000111101010001",
			949 => "00000000000000000000111101010001",
			950 => "0000001101000000000001000000001000",
			951 => "0000000110000000001010011000000100",
			952 => "00000000111100010000111101010001",
			953 => "11111110011100100000111101010001",
			954 => "0000001101000000000110010000011100",
			955 => "0000001110000000001011101100010000",
			956 => "0000000100000000000001011100001000",
			957 => "0000001010000000000000001000000100",
			958 => "00000000101111010000111101010001",
			959 => "00000010000100100000111101010001",
			960 => "0000001110000000001000001100000100",
			961 => "11111101100101000000111101010001",
			962 => "00000001110110010000111101010001",
			963 => "0000000111000000001000011000001000",
			964 => "0000001000000000000101000100000100",
			965 => "00000010111100000000111101010001",
			966 => "00000000000000000000111101010001",
			967 => "00000011111100110000111101010001",
			968 => "0000001100000000000100000100000100",
			969 => "11111110010000010000111101010001",
			970 => "00000000110000100000111101010001",
			971 => "0000000100000000000101000000010000",
			972 => "0000000110000000001000010000000100",
			973 => "11111110011010000000111101010001",
			974 => "0000000101000000001111010000000100",
			975 => "11111110100011000000111101010001",
			976 => "0000000001000000001010011000000100",
			977 => "00000011001111110000111101010001",
			978 => "11111110110000010000111101010001",
			979 => "11111110011000010000111101010001",
			980 => "0000000000000000000111000101000000",
			981 => "0000000110000000001101011000110000",
			982 => "0000000001000000001011111100100100",
			983 => "0000000011000000000110111100010000",
			984 => "0000000110000000001101111100000100",
			985 => "00000000000000000000111111011101",
			986 => "0000000100000000000111010100001000",
			987 => "0000001010000000000000001000000100",
			988 => "00000000000000000000111111011101",
			989 => "00000000100101000000111111011101",
			990 => "00000000000000000000111111011101",
			991 => "0000001100000000001001110100001100",
			992 => "0000000110000000001101111100000100",
			993 => "00000000000000000000111111011101",
			994 => "0000000001000000000001000100000100",
			995 => "11111111100101000000111111011101",
			996 => "00000000000000000000111111011101",
			997 => "0000001111000000000111011000000100",
			998 => "00000000000000000000111111011101",
			999 => "00000000010111100000111111011101",
			1000 => "0000001010000000000010101100001000",
			1001 => "0000000111000000001001001000000100",
			1002 => "00000000000000000000111111011101",
			1003 => "11111111010011110000111111011101",
			1004 => "00000000000000000000111111011101",
			1005 => "0000001001000000001001111100000100",
			1006 => "00000000000000000000111111011101",
			1007 => "0000001100000000000100011000000100",
			1008 => "00000000000000000000111111011101",
			1009 => "0000000011000000000110111100000100",
			1010 => "00000000000000000000111111011101",
			1011 => "00000001000100000000111111011101",
			1012 => "0000000110000000000100111100000100",
			1013 => "11111111001011010000111111011101",
			1014 => "00000000000000000000111111011101",
			1015 => "0000001111000000001100000000001100",
			1016 => "0000000100000000001100010000000100",
			1017 => "00000000000000000001000010001001",
			1018 => "0000001000000000001000100100000100",
			1019 => "11111111001111110001000010001001",
			1020 => "00000000000000000001000010001001",
			1021 => "0000000100000000000001011100100000",
			1022 => "0000001010000000000010101100010100",
			1023 => "0000000101000000001111010000001100",
			1024 => "0000000010000000001100010000000100",
			1025 => "00000000000000000001000010001001",
			1026 => "0000000101000000001100100100000100",
			1027 => "00000000000000000001000010001001",
			1028 => "11111111010111110001000010001001",
			1029 => "0000000001000000001001011000000100",
			1030 => "00000000000000000001000010001001",
			1031 => "00000000100010110001000010001001",
			1032 => "0000000000000000001111001000001000",
			1033 => "0000001101000000001110000100000100",
			1034 => "00000000000000000001000010001001",
			1035 => "00000001000011100001000010001001",
			1036 => "00000000000000000001000010001001",
			1037 => "0000000010000000001000100000001100",
			1038 => "0000000110000000001111000000001000",
			1039 => "0000000111000000001001001000000100",
			1040 => "00000000000000000001000010001001",
			1041 => "11111111001010100001000010001001",
			1042 => "00000000000000000001000010001001",
			1043 => "0000000000000000000001110100010000",
			1044 => "0000000111000000000110100100000100",
			1045 => "00000000000000000001000010001001",
			1046 => "0000000100000000001110000000001000",
			1047 => "0000000001000000001100011000000100",
			1048 => "00000000100111010001000010001001",
			1049 => "00000000000000000001000010001001",
			1050 => "00000000000000000001000010001001",
			1051 => "0000000110000000001000010000000100",
			1052 => "11111111101101000001000010001001",
			1053 => "0000000100000000000101000000001000",
			1054 => "0000001001000000001010100100000100",
			1055 => "00000000000000000001000010001001",
			1056 => "00000000001101110001000010001001",
			1057 => "00000000000000000001000010001001",
			1058 => "0000000100000000001000001100110000",
			1059 => "0000000001000000001011111100100100",
			1060 => "0000000011000000000111010100100000",
			1061 => "0000001010000000000000001000010000",
			1062 => "0000000011000000001100010000001100",
			1063 => "0000000011000000000111100000000100",
			1064 => "00000000000000000001000101001101",
			1065 => "0000000101000000001100100100000100",
			1066 => "00000000001010110001000101001101",
			1067 => "00000000000000000001000101001101",
			1068 => "00000000000000000001000101001101",
			1069 => "0000000111000000001001001000000100",
			1070 => "00000000000000000001000101001101",
			1071 => "0000000001000000001001011000000100",
			1072 => "00000000000000000001000101001101",
			1073 => "0000000000000000000101000100000100",
			1074 => "00000000000000000001000101001101",
			1075 => "00000000110101000001000101001101",
			1076 => "00000000000000000001000101001101",
			1077 => "0000001011000000000101100100001000",
			1078 => "0000001010000000000010101100000100",
			1079 => "11111111110010000001000101001101",
			1080 => "00000000000000000001000101001101",
			1081 => "00000000000000000001000101001101",
			1082 => "0000000110000000000100111100100000",
			1083 => "0000000100000000001011101100010100",
			1084 => "0000001010000000000010101100001100",
			1085 => "0000001011000000000100010000001000",
			1086 => "0000000101000000001110101000000100",
			1087 => "00000000000000000001000101001101",
			1088 => "11111111010011010001000101001101",
			1089 => "00000000000000000001000101001101",
			1090 => "0000000011000000000110111100000100",
			1091 => "00000000000000000001000101001101",
			1092 => "00000000011010000001000101001101",
			1093 => "0000001011000000001010010100001000",
			1094 => "0000000110000000001001100100000100",
			1095 => "11111110111110100001000101001101",
			1096 => "00000000000000000001000101001101",
			1097 => "00000000000000000001000101001101",
			1098 => "0000001001000000001010100000000100",
			1099 => "00000000000000000001000101001101",
			1100 => "0000000000000000001010101100001100",
			1101 => "0000001011000000001010010100001000",
			1102 => "0000001011000000001011011100000100",
			1103 => "00000000000000000001000101001101",
			1104 => "00000000011011100001000101001101",
			1105 => "00000000000000000001000101001101",
			1106 => "00000000000000000001000101001101",
			1107 => "0000001100000000000100011000011100",
			1108 => "0000001110000000000111010100010000",
			1109 => "0000000000000000001001101000001100",
			1110 => "0000001010000000000010101100001000",
			1111 => "0000001000000000001000010100000100",
			1112 => "00000000000000000001000111111001",
			1113 => "11111111101010000001000111111001",
			1114 => "00000000000000000001000111111001",
			1115 => "11111110110110110001000111111001",
			1116 => "0000000000000000000001110100001000",
			1117 => "0000001001000000000111101100000100",
			1118 => "00000000000000000001000111111001",
			1119 => "00000000010001100001000111111001",
			1120 => "00000000000000000001000111111001",
			1121 => "0000000000000000000010101000111000",
			1122 => "0000001110000000001100000000011100",
			1123 => "0000000101000000000111100000010000",
			1124 => "0000000100000000001100010000000100",
			1125 => "00000000000000000001000111111001",
			1126 => "0000001011000000000000011100000100",
			1127 => "00000000000000000001000111111001",
			1128 => "0000000101000000000111100000000100",
			1129 => "11111111011011010001000111111001",
			1130 => "00000000000000000001000111111001",
			1131 => "0000001010000000000000001000000100",
			1132 => "00000000000000000001000111111001",
			1133 => "0000000010000000001100000000000100",
			1134 => "00000000100101000001000111111001",
			1135 => "00000000000000000001000111111001",
			1136 => "0000000001000000000000111100001000",
			1137 => "0000000011000000001011111000000100",
			1138 => "00000000000000000001000111111001",
			1139 => "11111111111111110001000111111001",
			1140 => "0000000001000000001101111100001000",
			1141 => "0000000000000000000111000100000100",
			1142 => "00000001000000100001000111111001",
			1143 => "00000000000000000001000111111001",
			1144 => "0000000101000000001100100100000100",
			1145 => "11111111111101000001000111111001",
			1146 => "0000000101000000000101110000000100",
			1147 => "00000000010001110001000111111001",
			1148 => "00000000000000000001000111111001",
			1149 => "11111111110011000001000111111001",
			1150 => "0000001111000000001100000000001100",
			1151 => "0000000100000000001100010000000100",
			1152 => "00000000000000000001001010101101",
			1153 => "0000001000000000001000100100000100",
			1154 => "11111111010100000001001010101101",
			1155 => "00000000000000000001001010101101",
			1156 => "0000000100000000000001011100100000",
			1157 => "0000000110000000001101011000010100",
			1158 => "0000001011000000000110110100001000",
			1159 => "0000000101000000001100100100000100",
			1160 => "00000000000000000001001010101101",
			1161 => "11111111010000110001001010101101",
			1162 => "0000000000000000000001010100000100",
			1163 => "00000000000000000001001010101101",
			1164 => "0000001101000000000100101000000100",
			1165 => "00000000000000000001001010101101",
			1166 => "00000000100101110001001010101101",
			1167 => "0000000000000000001111001000001000",
			1168 => "0000001101000000001110000100000100",
			1169 => "00000000000000000001001010101101",
			1170 => "00000000111100110001001010101101",
			1171 => "00000000000000000001001010101101",
			1172 => "0000000010000000001000100000010000",
			1173 => "0000000110000000001111000000001100",
			1174 => "0000000111000000001001001000000100",
			1175 => "00000000000000000001001010101101",
			1176 => "0000001011000000000101100100000100",
			1177 => "00000000000000000001001010101101",
			1178 => "11111111001100110001001010101101",
			1179 => "00000000000000000001001010101101",
			1180 => "0000000000000000000001110100010000",
			1181 => "0000000111000000000110100100000100",
			1182 => "00000000000000000001001010101101",
			1183 => "0000000100000000001110000000001000",
			1184 => "0000000001000000001100011000000100",
			1185 => "00000000100101100001001010101101",
			1186 => "00000000000000000001001010101101",
			1187 => "00000000000000000001001010101101",
			1188 => "0000000110000000001000010000000100",
			1189 => "11111111101111110001001010101101",
			1190 => "0000000010000000001011110000001000",
			1191 => "0000000001000000001100011000000100",
			1192 => "00000000000000000001001010101101",
			1193 => "00000000001010110001001010101101",
			1194 => "00000000000000000001001010101101",
			1195 => "0000000000000000000010101001000100",
			1196 => "0000000001000000001001011000010000",
			1197 => "0000000110000000000000111100001000",
			1198 => "0000001001000000000001000100000100",
			1199 => "11111110101110100001001101001001",
			1200 => "00000010000110000001001101001001",
			1201 => "0000001001000000001111000000000100",
			1202 => "11111110010110110001001101001001",
			1203 => "00000000000000000001001101001001",
			1204 => "0000001101000000000110010000101100",
			1205 => "0000000111000000000110100100010100",
			1206 => "0000000000000000001111001000010000",
			1207 => "0000001100000000000100011000001000",
			1208 => "0000000010000000001100010000000100",
			1209 => "00000000110101100001001101001001",
			1210 => "11111110111101010001001101001001",
			1211 => "0000001011000000000100000100000100",
			1212 => "00000000000000000001001101001001",
			1213 => "00000001100111100001001101001001",
			1214 => "11111110011001000001001101001001",
			1215 => "0000000011000000001100111000010000",
			1216 => "0000000000000000000111000100001000",
			1217 => "0000000001000000001101111100000100",
			1218 => "00000001010010110001001101001001",
			1219 => "11111111011010110001001101001001",
			1220 => "0000001011000000001011011100000100",
			1221 => "11111110001101100001001101001001",
			1222 => "00000000000000000001001101001001",
			1223 => "0000000110000000001000010000000100",
			1224 => "00000001101111100001001101001001",
			1225 => "00000010100110010001001101001001",
			1226 => "0000000111000000000101110100000100",
			1227 => "11111110011100010001001101001001",
			1228 => "00000000110011000001001101001001",
			1229 => "0000000000000000001010101100001000",
			1230 => "0000000110000000001000010000000100",
			1231 => "11111110011101010001001101001001",
			1232 => "00000010011001110001001101001001",
			1233 => "11111110011001010001001101001001",
			1234 => "0000000000000000000010101001000000",
			1235 => "0000000011000000001100111000110000",
			1236 => "0000000000000000001111001000101000",
			1237 => "0000000110000000001011001100100000",
			1238 => "0000000010000000000111011000010000",
			1239 => "0000000001000000001001011000001000",
			1240 => "0000000000000000000110011100000100",
			1241 => "00000000000000000001001111010101",
			1242 => "11111111001010000001001111010101",
			1243 => "0000001011000000000100010000000100",
			1244 => "00000000101010110001001111010101",
			1245 => "11111111111010100001001111010101",
			1246 => "0000001100000000001011000000001000",
			1247 => "0000001100000000001010111000000100",
			1248 => "00000000000000000001001111010101",
			1249 => "11111111001011100001001111010101",
			1250 => "0000000001000000000001000100000100",
			1251 => "11111111101111010001001111010101",
			1252 => "00000000111000110001001111010101",
			1253 => "0000000011000000001010000100000100",
			1254 => "00000000000000000001001111010101",
			1255 => "00000001011001010001001111010101",
			1256 => "0000000011000000001000100000000100",
			1257 => "11111110101000010001001111010101",
			1258 => "00000000000000000001001111010101",
			1259 => "0000000010000000001101101100000100",
			1260 => "00000001001101000001001111010101",
			1261 => "0000001101000000001110010000000100",
			1262 => "00000000010010110001001111010101",
			1263 => "0000000010000000000011000000000100",
			1264 => "11111111101100110001001111010101",
			1265 => "00000000000000000001001111010101",
			1266 => "0000001001000000000010101100000100",
			1267 => "11111110100011010001001111010101",
			1268 => "00000000000000000001001111010101",
			1269 => "0000000100000000001011110000111100",
			1270 => "0000001001000000001111000000010000",
			1271 => "0000001110000000000010000100001100",
			1272 => "0000000110000000000000111100001000",
			1273 => "0000000110000000000000111100000100",
			1274 => "11111110011011110001010010111001",
			1275 => "00000001101101010001010010111001",
			1276 => "11111110010111010001010010111001",
			1277 => "00000001011011010001010010111001",
			1278 => "0000001101000000001110000100001100",
			1279 => "0000000001000000001011111100001000",
			1280 => "0000000100000000000111010100000100",
			1281 => "00000011010100010001010010111001",
			1282 => "11111110111010100001010010111001",
			1283 => "11111110010110100001010010111001",
			1284 => "0000000001000000000100110100011000",
			1285 => "0000001010000000000000001000001000",
			1286 => "0000000101000000001100100100000100",
			1287 => "00000010000100000001010010111001",
			1288 => "11111110011001100001010010111001",
			1289 => "0000000100000000000110111000001000",
			1290 => "0000000001000000001001011000000100",
			1291 => "00000000000000000001010010111001",
			1292 => "00000011011010110001010010111001",
			1293 => "0000000011000000001100111000000100",
			1294 => "11111110101111000001010010111001",
			1295 => "00000111100001100001010010111001",
			1296 => "0000001100000000001011000000000100",
			1297 => "00000000111000010001010010111001",
			1298 => "11111110011011100001010010111001",
			1299 => "0000000100000000001000110100011000",
			1300 => "0000000110000000001000010000010000",
			1301 => "0000000110000000001000010000001000",
			1302 => "0000000100000000001110000000000100",
			1303 => "11111110111100110001010010111001",
			1304 => "11111110010111000001010010111001",
			1305 => "0000000100000000001000000100000100",
			1306 => "00000000111111110001010010111001",
			1307 => "11111110101101000001010010111001",
			1308 => "0000000011000000001000101000000100",
			1309 => "11111110100001010001010010111001",
			1310 => "00000110011001010001010010111001",
			1311 => "0000000100000000000101000000011100",
			1312 => "0000000100000000000101000000010000",
			1313 => "0000001000000000000001110000000100",
			1314 => "11111110010111100001010010111001",
			1315 => "0000001000000000001100000100001000",
			1316 => "0000001000000000000001110000000100",
			1317 => "00000000110100100001010010111001",
			1318 => "11111111111110100001010010111001",
			1319 => "11111110011001010001010010111001",
			1320 => "0000001000000000000001110000000100",
			1321 => "11111110100000000001010010111001",
			1322 => "0000000001000000001101111100000100",
			1323 => "11111110100110100001010010111001",
			1324 => "00000100011011100001010010111001",
			1325 => "11111110010111000001010010111001",
			1326 => "0000000000000000000111000101000100",
			1327 => "0000000011000000000110111100011100",
			1328 => "0000001001000000001111000000001100",
			1329 => "0000001001000000001111000000000100",
			1330 => "11001001011010100001010110101101",
			1331 => "0000001010000000000000001000000100",
			1332 => "11001001110000000001010110101101",
			1333 => "11010011001000100001010110101101",
			1334 => "0000000000000000001100000100001000",
			1335 => "0000001100000000001000000000000100",
			1336 => "11110110000010010001010110101101",
			1337 => "11100101000100000001010110101101",
			1338 => "0000001101000000000101001000000100",
			1339 => "11001001011001010001010110101101",
			1340 => "11011101000110010001010110101101",
			1341 => "0000001101000000000101001000001000",
			1342 => "0000001101000000001110000100000100",
			1343 => "11001001100001000001010110101101",
			1344 => "11010101001000100001010110101101",
			1345 => "0000001001000000001111000000010000",
			1346 => "0000000110000000000100110100001000",
			1347 => "0000001000000000001000100100000100",
			1348 => "11001001100010100001010110101101",
			1349 => "11010100001011110001010110101101",
			1350 => "0000000111000000001000011000000100",
			1351 => "11001111111111100001010110101101",
			1352 => "11101000100101010001010110101101",
			1353 => "0000000001000000000100110100001100",
			1354 => "0000000100000000000110111000001000",
			1355 => "0000001000000000001000100100000100",
			1356 => "11100111000000010001010110101101",
			1357 => "11110100110111100001010110101101",
			1358 => "11100000110101010001010110101101",
			1359 => "11001001101010000001010110101101",
			1360 => "0000000000000000000001110100011000",
			1361 => "0000001000000000000101000100010100",
			1362 => "0000000110000000000100111100001100",
			1363 => "0000000110000000000100111100000100",
			1364 => "11001001011011000001010110101101",
			1365 => "0000000100000000001011110000000100",
			1366 => "11001101001010110001010110101101",
			1367 => "11001001110100110001010110101101",
			1368 => "0000000001000000001010011000000100",
			1369 => "11010101001000100001010110101101",
			1370 => "11001001110110110001010110101101",
			1371 => "11101001000011000001010110101101",
			1372 => "0000000000000000001010101100011000",
			1373 => "0000000110000000001000010000010100",
			1374 => "0000001000000000000001010100001100",
			1375 => "0000001000000000000001010100000100",
			1376 => "11001001011000100001010110101101",
			1377 => "0000000100000000001000000100000100",
			1378 => "11001101001010110001010110101101",
			1379 => "11001001011111000001010110101101",
			1380 => "0000000001000000001010011000000100",
			1381 => "11011001000111010001010110101101",
			1382 => "11001001111110110001010110101101",
			1383 => "11101101000001110001010110101101",
			1384 => "0000000000000000001010101100000100",
			1385 => "11001001101010010001010110101101",
			1386 => "11001001011000000001010110101101",
			1387 => "0000001001000000000111101101010000",
			1388 => "0000000000000000001001101000111100",
			1389 => "0000000101000000001100100100011000",
			1390 => "0000001000000000001000100100010000",
			1391 => "0000001001000000001000010000001100",
			1392 => "0000001100000000000100011000000100",
			1393 => "00000000000000000001011010101001",
			1394 => "0000000011000000001100000000000100",
			1395 => "00000000010001000001011010101001",
			1396 => "00000000000000000001011010101001",
			1397 => "11111111101010000001011010101001",
			1398 => "0000000101000000000110100000000100",
			1399 => "00000000000000000001011010101001",
			1400 => "00000000111111000001011010101001",
			1401 => "0000000101000000000111100000001100",
			1402 => "0000001111000000001111010100001000",
			1403 => "0000000110000000000100110100000100",
			1404 => "00000000000000000001011010101001",
			1405 => "00000000000001100001011010101001",
			1406 => "11111111000101000001011010101001",
			1407 => "0000000001000000000000111100010000",
			1408 => "0000000011000000001111010100001000",
			1409 => "0000001001000000001111000000000100",
			1410 => "00000000100010110001011010101001",
			1411 => "00000000000000000001011010101001",
			1412 => "0000000111000000001111011100000100",
			1413 => "11111111011001110001011010101001",
			1414 => "00000000000000000001011010101001",
			1415 => "0000001000000000000110011000000100",
			1416 => "00000000011101110001011010101001",
			1417 => "00000000000000000001011010101001",
			1418 => "0000001100000000000100011000001000",
			1419 => "0000000001000000000001111000000100",
			1420 => "11111110111110100001011010101001",
			1421 => "00000000000000000001011010101001",
			1422 => "0000000001000000000001000100000100",
			1423 => "11111111111101010001011010101001",
			1424 => "0000001001000000000100101100000100",
			1425 => "00000000010011110001011010101001",
			1426 => "00000000000000000001011010101001",
			1427 => "0000000000000000000111000100010000",
			1428 => "0000000110000000001011001100000100",
			1429 => "00000000000000000001011010101001",
			1430 => "0000000011000000000111010100000100",
			1431 => "00000000000000000001011010101001",
			1432 => "0000000101000000001001010000000100",
			1433 => "00000001000010100001011010101001",
			1434 => "00000000000000000001011010101001",
			1435 => "0000001110000000001100111000001100",
			1436 => "0000001100000000000100011000000100",
			1437 => "00000000000000000001011010101001",
			1438 => "0000000011000000000011000000000100",
			1439 => "11111111011101110001011010101001",
			1440 => "00000000000000000001011010101001",
			1441 => "0000001111000000001110000000010000",
			1442 => "0000000110000000001000010000000100",
			1443 => "00000000000000000001011010101001",
			1444 => "0000000101000000000001000000000100",
			1445 => "00000000000000000001011010101001",
			1446 => "0000001010000000001001000100000100",
			1447 => "00000000110110100001011010101001",
			1448 => "00000000000000000001011010101001",
			1449 => "00000000000000000001011010101001",
			1450 => "0000001100000000001010111000001100",
			1451 => "0000001110000000000111010100001000",
			1452 => "0000000101000000001101000100000100",
			1453 => "11111111000011000001011101110101",
			1454 => "00000000000000000001011101110101",
			1455 => "00000000000000000001011101110101",
			1456 => "0000001100000000001000000000110000",
			1457 => "0000000101000000000101001000100000",
			1458 => "0000001001000000000111101100001100",
			1459 => "0000000000000000000110001000001000",
			1460 => "0000000111000000001111011100000100",
			1461 => "00000000111000000001011101110101",
			1462 => "00000000000000000001011101110101",
			1463 => "00000000000000000001011101110101",
			1464 => "0000000110000000001011001100001000",
			1465 => "0000001001000000000000001000000100",
			1466 => "11111111011000100001011101110101",
			1467 => "00000000000000000001011101110101",
			1468 => "0000000000000000000001110100001000",
			1469 => "0000000110000000000100111100000100",
			1470 => "00000000110100110001011101110101",
			1471 => "00000000000000000001011101110101",
			1472 => "00000000000000000001011101110101",
			1473 => "0000001001000000000101010000001000",
			1474 => "0000000011000000001010000100000100",
			1475 => "00000000000000000001011101110101",
			1476 => "11111111100100000001011101110101",
			1477 => "0000000000000000001010101100000100",
			1478 => "00000000011011110001011101110101",
			1479 => "00000000000000000001011101110101",
			1480 => "0000000101000000001110000100001000",
			1481 => "0000000111000000001000011000000100",
			1482 => "11111111011001100001011101110101",
			1483 => "00000000000000000001011101110101",
			1484 => "0000001100000000001001110100010100",
			1485 => "0000001100000000001001001000001100",
			1486 => "0000000101000000000010011100001000",
			1487 => "0000001101000000001010001000000100",
			1488 => "00000000001100100001011101110101",
			1489 => "00000000000000000001011101110101",
			1490 => "00000000000000000001011101110101",
			1491 => "0000000010000000001000101000000100",
			1492 => "11111111101110110001011101110101",
			1493 => "00000000000000000001011101110101",
			1494 => "0000000010000000000010010100001100",
			1495 => "0000001111000000000111011000000100",
			1496 => "00000000000000000001011101110101",
			1497 => "0000000100000000001000110100000100",
			1498 => "00000000101011110001011101110101",
			1499 => "00000000000000000001011101110101",
			1500 => "00000000000000000001011101110101",
			1501 => "0000001100000000000100011000100100",
			1502 => "0000000100000000001010000100001100",
			1503 => "0000001110000000001110101100000100",
			1504 => "00000000000000000001100001110001",
			1505 => "0000000010000000001110110100000100",
			1506 => "00000000000100000001100001110001",
			1507 => "00000000000000000001100001110001",
			1508 => "0000001001000000000000001000001100",
			1509 => "0000000000000000001001101000001000",
			1510 => "0000000000000000001100000100000100",
			1511 => "11111111011001110001100001110001",
			1512 => "00000000000000000001100001110001",
			1513 => "11111110101101110001100001110001",
			1514 => "0000000000000000000001110100001000",
			1515 => "0000001110000000000111010100000100",
			1516 => "00000000000000000001100001110001",
			1517 => "00000000011010000001100001110001",
			1518 => "00000000000000000001100001110001",
			1519 => "0000000110000000001101111100011000",
			1520 => "0000000010000000001110110100010000",
			1521 => "0000000011000000001100000000001100",
			1522 => "0000000011000000000010000000000100",
			1523 => "00000000000000000001100001110001",
			1524 => "0000001101000000000010011100000100",
			1525 => "00000000001000010001100001110001",
			1526 => "00000000000000000001100001110001",
			1527 => "11111111111100110001100001110001",
			1528 => "0000001101000000000111111100000100",
			1529 => "00000000000000000001100001110001",
			1530 => "00000000111001010001100001110001",
			1531 => "0000001100000000000100011000010000",
			1532 => "0000000110000000000100111100001100",
			1533 => "0000000000000000000001110100001000",
			1534 => "0000001101000000000001000000000100",
			1535 => "00000000000000000001100001110001",
			1536 => "00000000110111100001100001110001",
			1537 => "00000000000000000001100001110001",
			1538 => "00000000000000000001100001110001",
			1539 => "0000000101000000000111100000010100",
			1540 => "0000001001000000000101010000001000",
			1541 => "0000001001000000001111000000000100",
			1542 => "00000000000000000001100001110001",
			1543 => "00000000000001000001100001110001",
			1544 => "0000001010000000000010101100000100",
			1545 => "11111110110111010001100001110001",
			1546 => "0000001001000000000000001000000100",
			1547 => "00000000000001110001100001110001",
			1548 => "11111111100110100001100001110001",
			1549 => "0000000001000000000101011100010000",
			1550 => "0000000110000000001010011000001000",
			1551 => "0000001100000000001001110100000100",
			1552 => "11111111111010010001100001110001",
			1553 => "00000000101000000001100001110001",
			1554 => "0000000011000000001000100000000100",
			1555 => "00000000000000000001100001110001",
			1556 => "11111111010111000001100001110001",
			1557 => "0000000000000000000001110100001000",
			1558 => "0000000011000000000010010100000100",
			1559 => "00000000111110010001100001110001",
			1560 => "00000000000000000001100001110001",
			1561 => "0000001110000000001101101100000100",
			1562 => "11111111011100110001100001110001",
			1563 => "00000000001000010001100001110001",
			1564 => "0000001100000000001010111000011000",
			1565 => "0000000000000000000110001000010100",
			1566 => "0000000010000000000111011000001100",
			1567 => "0000001100000000001010111000001000",
			1568 => "0000000111000000000110100100000100",
			1569 => "11111111011100010001100101011101",
			1570 => "00000000000000000001100101011101",
			1571 => "00000000000000000001100101011101",
			1572 => "0000001101000000000101001000000100",
			1573 => "00000000000000000001100101011101",
			1574 => "00000000110101100001100101011101",
			1575 => "11111110100010000001100101011101",
			1576 => "0000001100000000001011000000111000",
			1577 => "0000000101000000000101001000101100",
			1578 => "0000000001000000001101111100100000",
			1579 => "0000001101000000001111010000010000",
			1580 => "0000000101000000000010110100001000",
			1581 => "0000000000000000001011010100000100",
			1582 => "00000001000000000001100101011101",
			1583 => "00000000000000000001100101011101",
			1584 => "0000000101000000000110100000000100",
			1585 => "11111110110110100001100101011101",
			1586 => "00000000000000000001100101011101",
			1587 => "0000001101000000000100101000001000",
			1588 => "0000000110000000001101111100000100",
			1589 => "00000000000000000001100101011101",
			1590 => "00000001001100110001100101011101",
			1591 => "0000000101000000000111100000000100",
			1592 => "11111111011110110001100101011101",
			1593 => "00000000001101000001100101011101",
			1594 => "0000001101000000000100101000001000",
			1595 => "0000001100000000000100011000000100",
			1596 => "00000000000000000001100101011101",
			1597 => "11111111001101000001100101011101",
			1598 => "00000000000000000001100101011101",
			1599 => "0000000011000000001010000100000100",
			1600 => "00000000000000000001100101011101",
			1601 => "0000001001000000000101010000000100",
			1602 => "11111110110010000001100101011101",
			1603 => "00000000000000000001100101011101",
			1604 => "0000000010000000001110110100001100",
			1605 => "0000000001000000000000111100001000",
			1606 => "0000000100000000000010000100000100",
			1607 => "00000000000000000001100101011101",
			1608 => "11111111110000000001100101011101",
			1609 => "00000000000000000001100101011101",
			1610 => "0000001100000000000110100100010000",
			1611 => "0000001001000000000011101000001100",
			1612 => "0000000001000000001001011000000100",
			1613 => "00000000000000000001100101011101",
			1614 => "0000000000000000001010101100000100",
			1615 => "00000001001101010001100101011101",
			1616 => "00000000000000000001100101011101",
			1617 => "00000000000000000001100101011101",
			1618 => "0000001000000000001100011100001000",
			1619 => "0000000111000000001111011100000100",
			1620 => "00000000000000000001100101011101",
			1621 => "00000000101000100001100101011101",
			1622 => "11111111110010010001100101011101",
			1623 => "0000001001000000000111101101010000",
			1624 => "0000000100000000001111100101000000",
			1625 => "0000000101000000001100100100100000",
			1626 => "0000001101000000001111010000010100",
			1627 => "0000000001000000001011111100001000",
			1628 => "0000001100000000001010111000000100",
			1629 => "00000000000000000001101001101001",
			1630 => "00000000000010000001101001101001",
			1631 => "0000001010000000000010101100001000",
			1632 => "0000001100000000001010111000000100",
			1633 => "00000000000000000001101001101001",
			1634 => "11111111011010010001101001101001",
			1635 => "00000000000000000001101001101001",
			1636 => "0000000110000000001101111100000100",
			1637 => "00000000000000000001101001101001",
			1638 => "0000000010000000000010000000000100",
			1639 => "00000000000000000001101001101001",
			1640 => "00000000110001110001101001101001",
			1641 => "0000000111000000000001101000001100",
			1642 => "0000000110000000001010011000001000",
			1643 => "0000000011000000001100000000000100",
			1644 => "00000000000000000001101001101001",
			1645 => "11111111001010000001101001101001",
			1646 => "00000000000000000001101001101001",
			1647 => "0000000111000000001000011000001000",
			1648 => "0000000010000000000010000100000100",
			1649 => "00000000000000000001101001101001",
			1650 => "00000000011010100001101001101001",
			1651 => "0000000011000000000110111100000100",
			1652 => "00000000000000000001101001101001",
			1653 => "0000000111000000001111011100000100",
			1654 => "11111111101100000001101001101001",
			1655 => "00000000000000000001101001101001",
			1656 => "0000001100000000000110100100001100",
			1657 => "0000001001000000000111101100001000",
			1658 => "0000001000000000000110011000000100",
			1659 => "00000000000000000001101001101001",
			1660 => "11111110111011010001101001101001",
			1661 => "00000000000000000001101001101001",
			1662 => "00000000000000000001101001101001",
			1663 => "0000000111000000000001101000011000",
			1664 => "0000000110000000001011001100000100",
			1665 => "00000000000000000001101001101001",
			1666 => "0000000010000000001101101100010000",
			1667 => "0000000011000000001000001100000100",
			1668 => "00000000000000000001101001101001",
			1669 => "0000001010000000001000100100001000",
			1670 => "0000001101000000000101001000000100",
			1671 => "00000000000000000001101001101001",
			1672 => "00000000111011100001101001101001",
			1673 => "00000000000000000001101001101001",
			1674 => "00000000000000000001101001101001",
			1675 => "0000001110000000001100111000001100",
			1676 => "0000000100000000001011101100000100",
			1677 => "00000000000000000001101001101001",
			1678 => "0000000011000000000011000000000100",
			1679 => "11111111110010010001101001101001",
			1680 => "00000000000000000001101001101001",
			1681 => "0000001111000000001110000000010000",
			1682 => "0000000101000000001110000100000100",
			1683 => "00000000000000000001101001101001",
			1684 => "0000000111000000000000011100001000",
			1685 => "0000001100000000000110100100000100",
			1686 => "00000000010011100001101001101001",
			1687 => "00000000000000000001101001101001",
			1688 => "00000000000000000001101001101001",
			1689 => "00000000000000000001101001101001",
			1690 => "0000000000000000001010101101000000",
			1691 => "0000001100000000000111001000001100",
			1692 => "0000000111000000000110100100000100",
			1693 => "11111110011000000001101011101101",
			1694 => "0000000110000000001101111100000100",
			1695 => "00000000000000000001101011101101",
			1696 => "00000000001000010001101011101101",
			1697 => "0000001010000000001000010100110000",
			1698 => "0000000000000000001111001000011100",
			1699 => "0000000110000000001101011000010000",
			1700 => "0000000000000000001001101000001000",
			1701 => "0000001011000000000100010000000100",
			1702 => "00000000011101010001101011101101",
			1703 => "00000001101000010001101011101101",
			1704 => "0000001100000000001011000000000100",
			1705 => "11111101100101000001101011101101",
			1706 => "11111111101000010001101011101101",
			1707 => "0000001110000000001111010100001000",
			1708 => "0000000001000000000111101000000100",
			1709 => "00000001010000100001101011101101",
			1710 => "11111110100111100001101011101101",
			1711 => "00000001110101100001101011101101",
			1712 => "0000000011000000001111100100000100",
			1713 => "11111101111010110001101011101101",
			1714 => "0000000001000000000100110100001000",
			1715 => "0000000000000000000010101000000100",
			1716 => "00000001011111100001101011101101",
			1717 => "11111111000101010001101011101101",
			1718 => "0000001010000000001000010100000100",
			1719 => "11111110101100010001101011101101",
			1720 => "00000000000101110001101011101101",
			1721 => "00000011010010110001101011101101",
			1722 => "11111110011010010001101011101101",
			1723 => "0000001100000000001010111000001000",
			1724 => "0000000000000000000110001000000100",
			1725 => "00000000000000000001101110111001",
			1726 => "11111111000000100001101110111001",
			1727 => "0000001100000000001000000000110000",
			1728 => "0000001011000000000101110100101000",
			1729 => "0000000111000000000110100100011000",
			1730 => "0000000111000000001001001000001100",
			1731 => "0000000000000000001111001000001000",
			1732 => "0000000111000000001011000000000100",
			1733 => "00000000000000000001101110111001",
			1734 => "00000000101011100001101110111001",
			1735 => "00000000000000000001101110111001",
			1736 => "0000001010000000000010101100001000",
			1737 => "0000001111000000001100010000000100",
			1738 => "00000000000000000001101110111001",
			1739 => "11111111001001100001101110111001",
			1740 => "00000000000000000001101110111001",
			1741 => "0000000000000000000010101000001100",
			1742 => "0000000110000000001101111100000100",
			1743 => "00000000000000000001101110111001",
			1744 => "0000000001000000001001011000000100",
			1745 => "00000000000000000001101110111001",
			1746 => "00000001000000100001101110111001",
			1747 => "00000000000000000001101110111001",
			1748 => "0000001001000000000101010000000100",
			1749 => "11111111100110000001101110111001",
			1750 => "00000000000000000001101110111001",
			1751 => "0000001011000000000100010000001100",
			1752 => "0000000110000000001000010000001000",
			1753 => "0000001100000000001001110100000100",
			1754 => "11111111001011110001101110111001",
			1755 => "00000000000000000001101110111001",
			1756 => "00000000000000000001101110111001",
			1757 => "0000001101000000001100010100010000",
			1758 => "0000000111000000001000011000000100",
			1759 => "00000000000000000001101110111001",
			1760 => "0000001100000000000001101000001000",
			1761 => "0000000000000000001000101100000100",
			1762 => "00000000111000010001101110111001",
			1763 => "00000000000000000001101110111001",
			1764 => "00000000000000000001101110111001",
			1765 => "0000000111000000000000011100001000",
			1766 => "0000001001000000000010101100000100",
			1767 => "11111111100000000001101110111001",
			1768 => "00000000000000000001101110111001",
			1769 => "0000000001000000000111101000001000",
			1770 => "0000001011000000001110101100000100",
			1771 => "00000000010000010001101110111001",
			1772 => "00000000000000000001101110111001",
			1773 => "00000000000000000001101110111001",
			1774 => "0000000000000000001010101101000100",
			1775 => "0000001100000000000111001000001100",
			1776 => "0000000111000000000110100100000100",
			1777 => "11111110010110000001110001000101",
			1778 => "0000000110000000001101111100000100",
			1779 => "00000000000000000001110001000101",
			1780 => "00000000001010000001110001000101",
			1781 => "0000001010000000001000010100110100",
			1782 => "0000001101000000000011001000100000",
			1783 => "0000001011000000000110110100010000",
			1784 => "0000000000000000001111001000001000",
			1785 => "0000001101000000000101110000000100",
			1786 => "00000001001101000001110001000101",
			1787 => "11111111010010110001110001000101",
			1788 => "0000001101000000000101110000000100",
			1789 => "11111110001101010001110001000101",
			1790 => "00000001000111010001110001000101",
			1791 => "0000000000000000000101000100001000",
			1792 => "0000000110000000000100110100000100",
			1793 => "11111110001001100001110001000101",
			1794 => "00000000010101010001110001000101",
			1795 => "0000000011000000001010000100000100",
			1796 => "00000010001101100001110001000101",
			1797 => "00000000111010000001110001000101",
			1798 => "0000000100000000001101101100001000",
			1799 => "0000000111000000001111011100000100",
			1800 => "00000000000000000001110001000101",
			1801 => "00000001011101010001110001000101",
			1802 => "0000000111000000000101110100001000",
			1803 => "0000001010000000001000010100000100",
			1804 => "11111110001101110001110001000101",
			1805 => "11111111111100010001110001000101",
			1806 => "00000000100001000001110001000101",
			1807 => "00000011110010010001110001000101",
			1808 => "11111110011010000001110001000101",
			1809 => "0000000111000000000110100100010000",
			1810 => "0000000000000000000001010100000100",
			1811 => "00000000000000000001110100111001",
			1812 => "0000000011000000000111010100001000",
			1813 => "0000001100000000001011000000000100",
			1814 => "11111110101110110001110100111001",
			1815 => "00000000000000000001110100111001",
			1816 => "00000000000000000001110100111001",
			1817 => "0000000111000000001000011001001000",
			1818 => "0000000101000000001100100100100100",
			1819 => "0000001110000000000110010000001000",
			1820 => "0000000001000000001011111100000100",
			1821 => "00000000000000000001110100111001",
			1822 => "11111111001101010001110100111001",
			1823 => "0000000001000000000111101000001100",
			1824 => "0000000000000000000110001000001000",
			1825 => "0000001010000000000000001000000100",
			1826 => "00000000000000000001110100111001",
			1827 => "00000000111101000001110100111001",
			1828 => "00000000000000000001110100111001",
			1829 => "0000000011000000000000010000001000",
			1830 => "0000000100000000001011101100000100",
			1831 => "00000000000000000001110100111001",
			1832 => "11111111010001100001110100111001",
			1833 => "0000001010000000001000100100000100",
			1834 => "00000000110010100001110100111001",
			1835 => "00000000000000000001110100111001",
			1836 => "0000001111000000000111011000010100",
			1837 => "0000001110000000000010000100001100",
			1838 => "0000001010000000000000001000001000",
			1839 => "0000000011000000001100010000000100",
			1840 => "00000000000000000001110100111001",
			1841 => "11111111101011110001110100111001",
			1842 => "00000000000000000001110100111001",
			1843 => "0000000011000000001010000100000100",
			1844 => "00000000101110100001110100111001",
			1845 => "00000000000000000001110100111001",
			1846 => "0000001100000000001001110100001100",
			1847 => "0000001100000000001010111000000100",
			1848 => "00000000000000000001110100111001",
			1849 => "0000000111000000000110100100000100",
			1850 => "00000000000000000001110100111001",
			1851 => "11111111001100000001110100111001",
			1852 => "00000000000000000001110100111001",
			1853 => "0000000011000000001000100000010000",
			1854 => "0000000000000000000101000100000100",
			1855 => "00000000000000000001110100111001",
			1856 => "0000000100000000000011000000001000",
			1857 => "0000000111000000001000011000000100",
			1858 => "00000000000000000001110100111001",
			1859 => "00000001001010100001110100111001",
			1860 => "00000000000000000001110100111001",
			1861 => "0000000001000000000001000100000100",
			1862 => "11111111100111000001110100111001",
			1863 => "0000000010000000000010010100001100",
			1864 => "0000000001000000001010011000001000",
			1865 => "0000000011000000000001011100000100",
			1866 => "00000000000000000001110100111001",
			1867 => "00000000101110010001110100111001",
			1868 => "00000000000000000001110100111001",
			1869 => "00000000000000000001110100111001",
			1870 => "0000000111000000000110100100010000",
			1871 => "0000000100000000001010000100000100",
			1872 => "00000000000000000001111000110101",
			1873 => "0000000010000000000110111100001000",
			1874 => "0000001100000000000100011000000100",
			1875 => "11111110111000110001111000110101",
			1876 => "00000000000000000001111000110101",
			1877 => "00000000000000000001111000110101",
			1878 => "0000000110000000001101011001000000",
			1879 => "0000000100000000000110101100110000",
			1880 => "0000001010000000001010100000011100",
			1881 => "0000000001000000001001011000001100",
			1882 => "0000000110000000001101111100001000",
			1883 => "0000001100000000001011000000000100",
			1884 => "00000000000000000001111000110101",
			1885 => "00000000100000010001111000110101",
			1886 => "00000000000000000001111000110101",
			1887 => "0000000110000000000100110100001000",
			1888 => "0000001110000000000010000000000100",
			1889 => "00000000000000000001111000110101",
			1890 => "11111111001011100001111000110101",
			1891 => "0000000011000000001100010000000100",
			1892 => "11111111101110110001111000110101",
			1893 => "00000000010001100001111000110101",
			1894 => "0000001011000000000101100100001100",
			1895 => "0000001111000000000110111100001000",
			1896 => "0000000001000000000101011100000100",
			1897 => "00000000000000000001111000110101",
			1898 => "00000000000101110001111000110101",
			1899 => "11111111110000100001111000110101",
			1900 => "0000000001000000000000111100000100",
			1901 => "00000000000000000001111000110101",
			1902 => "00000000111111000001111000110101",
			1903 => "0000000111000000000111010000001100",
			1904 => "0000000101000000001100100100000100",
			1905 => "00000000000000000001111000110101",
			1906 => "0000001100000000001001110100000100",
			1907 => "11111110111010010001111000110101",
			1908 => "00000000000000000001111000110101",
			1909 => "00000000000000010001111000110101",
			1910 => "0000000000000000001111001000010000",
			1911 => "0000000001000000001101111100001100",
			1912 => "0000001100000000000100011000000100",
			1913 => "00000000000000000001111000110101",
			1914 => "0000000011000000000110111100000100",
			1915 => "00000000000000000001111000110101",
			1916 => "00000001000101010001111000110101",
			1917 => "00000000000000000001111000110101",
			1918 => "0000000001000000001101111100001000",
			1919 => "0000001100000000001011011100000100",
			1920 => "11111111011111100001111000110101",
			1921 => "00000000000000000001111000110101",
			1922 => "0000000001000000000100110100001100",
			1923 => "0000001010000000001000010100001000",
			1924 => "0000000101000000001110101000000100",
			1925 => "00000000000000000001111000110101",
			1926 => "00000000110000100001111000110101",
			1927 => "00000000000000000001111000110101",
			1928 => "0000001010000000001000010100000100",
			1929 => "11111111011101000001111000110101",
			1930 => "0000000100000000000101000000000100",
			1931 => "00000000011100100001111000110101",
			1932 => "00000000000000000001111000110101",
			1933 => "0000001001000000001111000000010000",
			1934 => "0000001000000000000100101100001100",
			1935 => "0000000100000000000111010000000100",
			1936 => "00000000000000000001111100010001",
			1937 => "0000001010000000001001100100000100",
			1938 => "00000000000100000001111100010001",
			1939 => "00000000000000000001111100010001",
			1940 => "11111110011011110001111100010001",
			1941 => "0000001100000000000001101001010100",
			1942 => "0000001100000000000100011000110000",
			1943 => "0000000101000000000111100000011100",
			1944 => "0000001001000000001010100000010000",
			1945 => "0000000111000000000110100100001000",
			1946 => "0000001010000000001010100100000100",
			1947 => "00000000011110100001111100010001",
			1948 => "11111110110010100001111100010001",
			1949 => "0000001011000000000110110100000100",
			1950 => "00000001011010010001111100010001",
			1951 => "11111111101001110001111100010001",
			1952 => "0000001011000000001011011100000100",
			1953 => "11111101111011100001111100010001",
			1954 => "0000000001000000000100110100000100",
			1955 => "00000000010101010001111100010001",
			1956 => "00000000000000000001111100010001",
			1957 => "0000001011000000000010001000010000",
			1958 => "0000000110000000001001100100001000",
			1959 => "0000001110000000000010000100000100",
			1960 => "00000000000000000001111100010001",
			1961 => "11111110001101110001111100010001",
			1962 => "0000000001000000000100110100000100",
			1963 => "00000000000000000001111100010001",
			1964 => "11111111101010000001111100010001",
			1965 => "00000000000000000001111100010001",
			1966 => "0000000001000000001001011000001000",
			1967 => "0000000011000000000110111100000100",
			1968 => "00000010001001110001111100010001",
			1969 => "00000000001110110001111100010001",
			1970 => "0000000110000000000100110100001100",
			1971 => "0000001001000000001111000000000100",
			1972 => "00000000101010110001111100010001",
			1973 => "0000001001000000000100111100000100",
			1974 => "11111110101111110001111100010001",
			1975 => "00000000100100110001111100010001",
			1976 => "0000000010000000001100010000001000",
			1977 => "0000000001000000001110010100000100",
			1978 => "00000001010111010001111100010001",
			1979 => "00000000000000000001111100010001",
			1980 => "0000001110000000001100000000000100",
			1981 => "11111110111111110001111100010001",
			1982 => "00000000101000010001111100010001",
			1983 => "0000001001000000001000010000000100",
			1984 => "11111001011101100001111100010001",
			1985 => "0000000010000000001101101100000100",
			1986 => "00000000101010100001111100010001",
			1987 => "11111110111011000001111100010001",
			1988 => "0000001100000000001010111000010000",
			1989 => "0000000000000000000110001000001100",
			1990 => "0000001011000000000000011100000100",
			1991 => "00000000000000000010000000010101",
			1992 => "0000001000000000000111110100000100",
			1993 => "00000000000000000010000000010101",
			1994 => "00000000101000000010000000010101",
			1995 => "11111110011001110010000000010101",
			1996 => "0000000010000000000111011000110000",
			1997 => "0000000001000000001011111100100100",
			1998 => "0000000011000000001111010100011000",
			1999 => "0000000000000000000101000100001100",
			2000 => "0000001011000000000110110100001000",
			2001 => "0000000100000000001100010000000100",
			2002 => "00000000111011110010000000010101",
			2003 => "00000000000000000010000000010101",
			2004 => "11111111010100010010000000010101",
			2005 => "0000001010000000000000001000000100",
			2006 => "00000000000000000010000000010101",
			2007 => "0000001001000000001001100100000100",
			2008 => "00000000000000000010000000010101",
			2009 => "00000001100001010010000000010101",
			2010 => "0000001000000000001000100100001000",
			2011 => "0000000000000000000001010100000100",
			2012 => "11111111010101010010000000010101",
			2013 => "00000000000000000010000000010101",
			2014 => "00000000110101010010000000010101",
			2015 => "0000001110000000000110010000000100",
			2016 => "11111110101111000010000000010101",
			2017 => "0000000011000000000111011000000100",
			2018 => "00000000000000000010000000010101",
			2019 => "00000000011010100010000000010101",
			2020 => "0000001110000000000111010100101100",
			2021 => "0000000100000000001111100100011000",
			2022 => "0000001010000000000010101100010000",
			2023 => "0000000111000000001111011100001000",
			2024 => "0000001111000000001111010100000100",
			2025 => "00000000000000000010000000010101",
			2026 => "11111110110101010010000000010101",
			2027 => "0000001011000000000100010000000100",
			2028 => "00000000000000000010000000010101",
			2029 => "00000000010011110010000000010101",
			2030 => "0000001001000000000111101100000100",
			2031 => "00000001000110000010000000010101",
			2032 => "00000000000000000010000000010101",
			2033 => "0000000011000000000000010000001100",
			2034 => "0000001100000000001010111000000100",
			2035 => "00000000000000000010000000010101",
			2036 => "0000000110000000001001100100000100",
			2037 => "11111110011011100010000000010101",
			2038 => "00000000000000000010000000010101",
			2039 => "0000000110000000001001100100000100",
			2040 => "00000000000000110010000000010101",
			2041 => "00000000000000000010000000010101",
			2042 => "0000000100000000000001011100000100",
			2043 => "00000001001110000010000000010101",
			2044 => "0000000011000000001000100000000100",
			2045 => "11111110111011110010000000010101",
			2046 => "0000001011000000000101110100001000",
			2047 => "0000000001000000000100110100000100",
			2048 => "00000001001100100010000000010101",
			2049 => "00000000000000000010000000010101",
			2050 => "0000000111000000000101110100000100",
			2051 => "11111111000110100010000000010101",
			2052 => "00000000000000000010000000010101",
			2053 => "0000001001000000001111000000001000",
			2054 => "0000000110000000000000111100000100",
			2055 => "00000000000000000010000100001001",
			2056 => "11111110100000100010000100001001",
			2057 => "0000001001000000000111101101001000",
			2058 => "0000000000000000001100000100101000",
			2059 => "0000000000000000000001010100011000",
			2060 => "0000001101000000000101110000001000",
			2061 => "0000001101000000000010011100000100",
			2062 => "00000001000001000010000100001001",
			2063 => "00000000000000000010000100001001",
			2064 => "0000001111000000001100000000001000",
			2065 => "0000001000000000001000100100000100",
			2066 => "11111110100101000010000100001001",
			2067 => "00000000000000000010000100001001",
			2068 => "0000000010000000001100010000000100",
			2069 => "00000000001100010010000100001001",
			2070 => "11111111001110000010000100001001",
			2071 => "0000000010000000000010000000000100",
			2072 => "11111111100111010010000100001001",
			2073 => "0000001111000000001000001100001000",
			2074 => "0000000111000000000110100100000100",
			2075 => "00000000000000000010000100001001",
			2076 => "00000001001000000010000100001001",
			2077 => "00000000000000000010000100001001",
			2078 => "0000001100000000001000011000011000",
			2079 => "0000000100000000001101101100010000",
			2080 => "0000001011000000001011011100001000",
			2081 => "0000001010000000000010101100000100",
			2082 => "11111110100000010010000100001001",
			2083 => "11111111111010010010000100001001",
			2084 => "0000000001000000000101011100000100",
			2085 => "11111111011111000010000100001001",
			2086 => "00000000110111100010000100001001",
			2087 => "0000001100000000000110100100000100",
			2088 => "11111110100101110010000100001001",
			2089 => "00000000000000000010000100001001",
			2090 => "0000000100000000000110001100000100",
			2091 => "00000000110010110010000100001001",
			2092 => "00000000000000000010000100001001",
			2093 => "0000000000000000000001110100010100",
			2094 => "0000000110000000001011001100001000",
			2095 => "0000001001000000000111101100000100",
			2096 => "00000000000000000010000100001001",
			2097 => "11111111010011000010000100001001",
			2098 => "0000001110000000001111010100000100",
			2099 => "00000000000000000010000100001001",
			2100 => "0000000111000000000000011100000100",
			2101 => "00000001010001100010000100001001",
			2102 => "00000000000000000010000100001001",
			2103 => "0000001110000000001100111000000100",
			2104 => "11111110110010100010000100001001",
			2105 => "0000000110000000001000010000001000",
			2106 => "0000001010000000001000100100000100",
			2107 => "00000000000000000010000100001001",
			2108 => "11111111100110000010000100001001",
			2109 => "0000001111000000001110000000001000",
			2110 => "0000001011000000001011110100000100",
			2111 => "00000000111111100010000100001001",
			2112 => "00000000000000000010000100001001",
			2113 => "11111111111011110010000100001001",
			2114 => "0000000000000000001010101101110000",
			2115 => "0000000111000000001000011001001100",
			2116 => "0000000111000000001000011000111000",
			2117 => "0000000101000000001100100100011000",
			2118 => "0000000001000000000111101000001100",
			2119 => "0000000011000000001010000100001000",
			2120 => "0000000001000000001011111100000100",
			2121 => "00000000011110100010000111101101",
			2122 => "11111110101111110010000111101101",
			2123 => "00000001100011100010000111101101",
			2124 => "0000000101000000001101000100000100",
			2125 => "11111110000100100010000111101101",
			2126 => "0000001100000000000100011000000100",
			2127 => "00000000010111010010000111101101",
			2128 => "11111111000101000010000111101101",
			2129 => "0000001100000000000100011000010000",
			2130 => "0000000101000000001100100100001000",
			2131 => "0000000001000000000000111100000100",
			2132 => "00000000000000000010000111101101",
			2133 => "00000000111000010010000111101101",
			2134 => "0000001101000000000010011100000100",
			2135 => "00000000000000000010000111101101",
			2136 => "11111110110101100010000111101101",
			2137 => "0000000001000000000000111100001000",
			2138 => "0000000101000000001111010000000100",
			2139 => "00000000010100100010000111101101",
			2140 => "11111110111101100010000111101101",
			2141 => "0000000000000000000001110100000100",
			2142 => "00000001100110000010000111101101",
			2143 => "11111111001000010010000111101101",
			2144 => "0000000110000000000100110100000100",
			2145 => "00000000000000000010000111101101",
			2146 => "0000000110000000001011001100001000",
			2147 => "0000000011000000001111010100000100",
			2148 => "00000000000000000010000111101101",
			2149 => "11111110010001100010000111101101",
			2150 => "0000001001000000000000001000000100",
			2151 => "00000000000000000010000111101101",
			2152 => "11111111101100100010000111101101",
			2153 => "0000001100000000000001101000011000",
			2154 => "0000001101000000001100010100010000",
			2155 => "0000000000000000000101000100000100",
			2156 => "00000000000000000010000111101101",
			2157 => "0000001011000000000100010000001000",
			2158 => "0000001011000000000010001000000100",
			2159 => "00000001001100010010000111101101",
			2160 => "00000000000000000010000111101101",
			2161 => "00000001101010010010000111101101",
			2162 => "0000000101000000000011001000000100",
			2163 => "11111111011000010010000111101101",
			2164 => "00000000000000000010000111101101",
			2165 => "0000001001000000000101010000000100",
			2166 => "11111101111011110010000111101101",
			2167 => "0000000001000000000100110100000100",
			2168 => "00000000100000110010000111101101",
			2169 => "11111111110001000010000111101101",
			2170 => "11111110011101000010000111101101",
			2171 => "0000001100000000000111001000001000",
			2172 => "0000000111000000000110100100000100",
			2173 => "11111110011101100010001011101001",
			2174 => "00000000000000000010001011101001",
			2175 => "0000000110000000001101111100100000",
			2176 => "0000001101000000000111111100011100",
			2177 => "0000001011000000001011011100001100",
			2178 => "0000001100000000000100011000000100",
			2179 => "00000000000000000010001011101001",
			2180 => "0000001101000000000010011100000100",
			2181 => "00000000111111010010001011101001",
			2182 => "00000000000000000010001011101001",
			2183 => "0000000111000000000001101000001000",
			2184 => "0000001101000000000010011100000100",
			2185 => "00000000000000000010001011101001",
			2186 => "11111111001000000010001011101001",
			2187 => "0000000001000000001001011000000100",
			2188 => "00000000000000000010001011101001",
			2189 => "00000000011110110010001011101001",
			2190 => "00000001100010000010001011101001",
			2191 => "0000000101000000001100100100101000",
			2192 => "0000000001000000000111101000010100",
			2193 => "0000001110000000000111011000010000",
			2194 => "0000000001000000001011111100001000",
			2195 => "0000001000000000001100011100000100",
			2196 => "00000001000000100010001011101001",
			2197 => "11111111101001000010001011101001",
			2198 => "0000001100000000000100011000000100",
			2199 => "00000000000000000010001011101001",
			2200 => "11111110011101110010001011101001",
			2201 => "00000001100000010010001011101001",
			2202 => "0000001101000000000010011100001100",
			2203 => "0000000111000000001001001000000100",
			2204 => "00000000000000000010001011101001",
			2205 => "0000001010000000000011101000000100",
			2206 => "00000000000000000010001011101001",
			2207 => "11111110001100000010001011101001",
			2208 => "0000001010000000001000010100000100",
			2209 => "00000000001110000010001011101001",
			2210 => "00000000000000000010001011101001",
			2211 => "0000000101000000001100100100010100",
			2212 => "0000000001000000000100110100001100",
			2213 => "0000001101000000000100101000001000",
			2214 => "0000000010000000001101101100000100",
			2215 => "00000001100000110010001011101001",
			2216 => "00000000000000000010001011101001",
			2217 => "00000000000000000010001011101001",
			2218 => "0000000111000000000001101000000100",
			2219 => "00000000000000000010001011101001",
			2220 => "11111111100101000010001011101001",
			2221 => "0000001100000000000110100100010000",
			2222 => "0000000111000000001000011000001000",
			2223 => "0000000111000000001000011000000100",
			2224 => "00000000010010010010001011101001",
			2225 => "11111111001011110010001011101001",
			2226 => "0000001101000000001100010100000100",
			2227 => "00000001001011000010001011101001",
			2228 => "11111111110000000010001011101001",
			2229 => "0000001011000000000101110100000100",
			2230 => "11111110010110000010001011101001",
			2231 => "0000000110000000001001100100000100",
			2232 => "00000000110100100010001011101001",
			2233 => "11111111000000110010001011101001",
			2234 => "0000001100000000000111001000001000",
			2235 => "0000000111000000000110100100000100",
			2236 => "11111110011100010010001111010101",
			2237 => "00000000000000000010001111010101",
			2238 => "0000001100000000000001101001100000",
			2239 => "0000001100000000001011000000110100",
			2240 => "0000000111000000000001101000011100",
			2241 => "0000000111000000000110100100010000",
			2242 => "0000000111000000001001001000001000",
			2243 => "0000000000000000001111001000000100",
			2244 => "00000000110000110010001111010101",
			2245 => "00000000000000000010001111010101",
			2246 => "0000001010000000000010101100000100",
			2247 => "11111110100011100010001111010101",
			2248 => "00000000000000000010001111010101",
			2249 => "0000001000000000000111110100000100",
			2250 => "11111111100110100010001111010101",
			2251 => "0000000000000000000001110100000100",
			2252 => "00000001010010100010001111010101",
			2253 => "11111111111110110010001111010101",
			2254 => "0000001111000000001100010000001000",
			2255 => "0000001010000000000000001000000100",
			2256 => "00000000000000000010001111010101",
			2257 => "00000001100011100010001111010101",
			2258 => "0000001100000000001010111000001000",
			2259 => "0000001101000000000101110000000100",
			2260 => "11111101101111110010001111010101",
			2261 => "00000000000000000010001111010101",
			2262 => "0000000110000000000100110100000100",
			2263 => "11111110100111110010001111010101",
			2264 => "11111111110001000010001111010101",
			2265 => "0000001101000000000010011100010000",
			2266 => "0000001100000000001000000000001100",
			2267 => "0000000000000000000110001000001000",
			2268 => "0000000001000000001001011000000100",
			2269 => "00000000000000000010001111010101",
			2270 => "00000000111110100010001111010101",
			2271 => "00000000000000000010001111010101",
			2272 => "11111110101110110010001111010101",
			2273 => "0000001101000000001110010000010000",
			2274 => "0000000110000000000100110100001000",
			2275 => "0000000110000000001101111100000100",
			2276 => "00000001001101100010001111010101",
			2277 => "11111111110110010010001111010101",
			2278 => "0000000000000000001010101100000100",
			2279 => "00000001011110010010001111010101",
			2280 => "00000000000000000010001111010101",
			2281 => "0000000111000000001000011000000100",
			2282 => "11111111000010000010001111010101",
			2283 => "0000001101000000001100010100000100",
			2284 => "00000000111110010010001111010101",
			2285 => "11111111111011000010001111010101",
			2286 => "0000001011000000000101110100000100",
			2287 => "11111100001111100010001111010101",
			2288 => "0000000110000000001001100100000100",
			2289 => "00000000101001000010001111010101",
			2290 => "0000000111000000000111010000000100",
			2291 => "00000000000000000010001111010101",
			2292 => "11111110110100110010001111010101",
			2293 => "0000000000000000001010101110000000",
			2294 => "0000000001000000000000111101000000",
			2295 => "0000000111000000001000011000100100",
			2296 => "0000000111000000000001101000011000",
			2297 => "0000000011000000001100000000010000",
			2298 => "0000001100000000000100011000001000",
			2299 => "0000000111000000000110100100000100",
			2300 => "11111110101000000010010011011011",
			2301 => "00000000000000000010010011011011",
			2302 => "0000001001000000001111000000000100",
			2303 => "00000000010000000010010011011011",
			2304 => "00000010100110010010010011011011",
			2305 => "0000000101000000001100100100000100",
			2306 => "00000000000000000010010011011011",
			2307 => "11111110100100100010010011011011",
			2308 => "0000000000000000000101000100001000",
			2309 => "0000000011000000001100000000000100",
			2310 => "00000000000000000010010011011011",
			2311 => "11111111101111100010010011011011",
			2312 => "00000010011100010010010011011011",
			2313 => "0000000011000000000110111100001100",
			2314 => "0000000111000000001000011000001000",
			2315 => "0000000010000000000110010000000100",
			2316 => "00000000001001000010010011011011",
			2317 => "00000000000000000010010011011011",
			2318 => "00000011100001100010010011011011",
			2319 => "0000000000000000000001010100000100",
			2320 => "11111101101011110010010011011011",
			2321 => "0000000111000000001000011000000100",
			2322 => "11111101110100110010010011011011",
			2323 => "0000000010000000000110111100000100",
			2324 => "00000001010011110010010011011011",
			2325 => "11111110111011010010010011011011",
			2326 => "0000000111000000000001101000100000",
			2327 => "0000001100000000001001001000011100",
			2328 => "0000000000000000001111001000001100",
			2329 => "0000000001000000001101111100001000",
			2330 => "0000000101000000000110100000000100",
			2331 => "11111111101110000010010011011011",
			2332 => "00000001001100010010010011011011",
			2333 => "11111110010000110010010011011011",
			2334 => "0000000110000000001111000000001000",
			2335 => "0000001100000000001011000000000100",
			2336 => "11111110000101110010010011011011",
			2337 => "00000000000000000010010011011011",
			2338 => "0000000101000000001100100100000100",
			2339 => "11111110101100110010010011011011",
			2340 => "00000001001110110010010011011011",
			2341 => "11111110001101010010010011011011",
			2342 => "0000001101000000000110010000011000",
			2343 => "0000001001000000000100111100001000",
			2344 => "0000000010000000000111011000000100",
			2345 => "00000000101010000010010011011011",
			2346 => "11111111110011010010010011011011",
			2347 => "0000001011000000001011011100001000",
			2348 => "0000000000000000001111001000000100",
			2349 => "00000001000110000010010011011011",
			2350 => "11111111110000010010010011011011",
			2351 => "0000000000000000001010101100000100",
			2352 => "00000001100001100010010011011011",
			2353 => "00000011000011100010010011011011",
			2354 => "0000000111000000000101110100000100",
			2355 => "11111110101000100010010011011011",
			2356 => "00000000010100000010010011011011",
			2357 => "11111110011010010010010011011011",
			2358 => "00000000000000000010010011011101",
			2359 => "00000000000000000010010011100001",
			2360 => "00000000000000000010010011100101",
			2361 => "0000001100000000001011000000000100",
			2362 => "00000000000000000010010011111001",
			2363 => "0000001100000000000110100100000100",
			2364 => "00000000000010000010010011111001",
			2365 => "00000000000000000010010011111001",
			2366 => "0000001100000000001010111000000100",
			2367 => "00000000000000000010010100001101",
			2368 => "0000000000000000000001110100000100",
			2369 => "00000000000100010010010100001101",
			2370 => "00000000000000000010010100001101",
			2371 => "0000000000000000001100000100001000",
			2372 => "0000000000000000000011101000000100",
			2373 => "00000000000000000010010100100001",
			2374 => "00000000000001110010010100100001",
			2375 => "00000000000000000010010100100001",
			2376 => "0000000101000000001100100100001000",
			2377 => "0000000101000000000110110100000100",
			2378 => "00000000000000000010010100111101",
			2379 => "00000000000101010010010100111101",
			2380 => "0000000101000000001111010000000100",
			2381 => "11111111111100100010010100111101",
			2382 => "00000000000000000010010100111101",
			2383 => "0000000100000000001101101100001000",
			2384 => "0000000010000000001101000100000100",
			2385 => "00000000000000000010010101011001",
			2386 => "00000000000010110010010101011001",
			2387 => "0000000010000000001000101000000100",
			2388 => "11111111111101000010010101011001",
			2389 => "00000000000000000010010101011001",
			2390 => "0000001110000000000111010100001100",
			2391 => "0000000111000000000001101000001000",
			2392 => "0000001001000000001001111100000100",
			2393 => "11111111110010110010010101111101",
			2394 => "00000000000000000010010101111101",
			2395 => "00000000000000000010010101111101",
			2396 => "0000000010000000001101101100000100",
			2397 => "00000000001101100010010101111101",
			2398 => "00000000000000000010010101111101",
			2399 => "0000001100000000001001110100001100",
			2400 => "0000001100000000000100011000000100",
			2401 => "00000000000000000010010110100001",
			2402 => "0000001100000000001011000000000100",
			2403 => "11111111111011110010010110100001",
			2404 => "00000000000000000010010110100001",
			2405 => "0000001100000000000110100100000100",
			2406 => "00000000000000010010010110100001",
			2407 => "00000000000000000010010110100001",
			2408 => "0000000000000000001001101000001100",
			2409 => "0000000010000000000010000100000100",
			2410 => "00000000000000000010010111001101",
			2411 => "0000001100000000000100011000000100",
			2412 => "00000000000000000010010111001101",
			2413 => "00000000010001100010010111001101",
			2414 => "0000001100000000001001110100001000",
			2415 => "0000000010000000000010010100000100",
			2416 => "11111111110001110010010111001101",
			2417 => "00000000000000000010010111001101",
			2418 => "00000000000000000010010111001101",
			2419 => "0000000100000000001100010000000100",
			2420 => "00000000000000000010010111110001",
			2421 => "0000001011000000001011110100001100",
			2422 => "0000001110000000001100111000001000",
			2423 => "0000000011000000000001011100000100",
			2424 => "11111111101010110010010111110001",
			2425 => "00000000000000000010010111110001",
			2426 => "00000000000000000010010111110001",
			2427 => "00000000000000000010010111110001",
			2428 => "0000000100000000001101101100010000",
			2429 => "0000000101000000000110100000000100",
			2430 => "00000000000000000010011000010101",
			2431 => "0000000101000000000101001000001000",
			2432 => "0000000100000000000010000000000100",
			2433 => "00000000000000000010011000010101",
			2434 => "00000000000111110010011000010101",
			2435 => "00000000000000000010011000010101",
			2436 => "00000000000000000010011000010101",
			2437 => "0000001100000000001001110100010000",
			2438 => "0000000110000000001101111100000100",
			2439 => "00000000000000000010011001000001",
			2440 => "0000000110000000001001100100001000",
			2441 => "0000001011000000000000011100000100",
			2442 => "00000000000000000010011001000001",
			2443 => "11111111101110000010011001000001",
			2444 => "00000000000000000010011001000001",
			2445 => "0000001100000000000110100100000100",
			2446 => "00000000000000100010011001000001",
			2447 => "00000000000000000010011001000001",
			2448 => "0000000110000000001101111100001000",
			2449 => "0000001100000000000100011000000100",
			2450 => "00000000000000000010011001101101",
			2451 => "00000000010000110010011001101101",
			2452 => "0000001100000000001001110100001100",
			2453 => "0000000100000000001010000100000100",
			2454 => "00000000000000000010011001101101",
			2455 => "0000000110000000001011001100000100",
			2456 => "11111111110101010010011001101101",
			2457 => "00000000000000000010011001101101",
			2458 => "00000000000000000010011001101101",
			2459 => "0000000010000000001100010000001100",
			2460 => "0000000000000000001100000100001000",
			2461 => "0000000010000000001101000100000100",
			2462 => "00000000000000000010011010100001",
			2463 => "00000000001010100010011010100001",
			2464 => "00000000000000000010011010100001",
			2465 => "0000000010000000001010000100000100",
			2466 => "11111111111000110010011010100001",
			2467 => "0000000000000000000111000100001000",
			2468 => "0000000000000000001001101000000100",
			2469 => "00000000000000000010011010100001",
			2470 => "00000000000111100010011010100001",
			2471 => "00000000000000000010011010100001",
			2472 => "0000000100000000000001011100010100",
			2473 => "0000001010000000000000001000000100",
			2474 => "00000000000000000010011011010101",
			2475 => "0000000001000000000111101000001100",
			2476 => "0000001001000000001111000000000100",
			2477 => "00000000000000000010011011010101",
			2478 => "0000001110000000000010000000000100",
			2479 => "00000000000000000010011011010101",
			2480 => "00000000010010110010011011010101",
			2481 => "00000000000000000010011011010101",
			2482 => "0000001001000000001010100100000100",
			2483 => "11111111110100110010011011010101",
			2484 => "00000000000000000010011011010101",
			2485 => "0000000000000000000111000100010100",
			2486 => "0000001100000000001010111000000100",
			2487 => "00000000000000000010011100000001",
			2488 => "0000001101000000001010001000001100",
			2489 => "0000001101000000001110000100000100",
			2490 => "00000000000000000010011100000001",
			2491 => "0000001010000000000000001000000100",
			2492 => "00000000000000000010011100000001",
			2493 => "00000000010000000010011100000001",
			2494 => "00000000000000000010011100000001",
			2495 => "00000000000000000010011100000001",
			2496 => "0000000101000000001111010000010100",
			2497 => "0000001100000000000100011000000100",
			2498 => "00000000000000000010011100101101",
			2499 => "0000000000000000000010101000001100",
			2500 => "0000001100000000001001001000001000",
			2501 => "0000001101000000001001011100000100",
			2502 => "00000000011010010010011100101101",
			2503 => "00000000000000000010011100101101",
			2504 => "00000000000000000010011100101101",
			2505 => "00000000000000000010011100101101",
			2506 => "00000000000000000010011100101101",
			2507 => "0000000001000000000000111100001100",
			2508 => "0000000010000000001100010000000100",
			2509 => "00000000000000000010011101101001",
			2510 => "0000001101000000000111111100000100",
			2511 => "00000000000000000010011101101001",
			2512 => "11111111101011110010011101101001",
			2513 => "0000001100000000000100011000000100",
			2514 => "00000000000000000010011101101001",
			2515 => "0000000010000000000110111000001100",
			2516 => "0000000001000000001010011000001000",
			2517 => "0000001101000000000010011100000100",
			2518 => "00000000000000000010011101101001",
			2519 => "00000000010110110010011101101001",
			2520 => "00000000000000000010011101101001",
			2521 => "00000000000000000010011101101001",
			2522 => "0000000101000000000110100000001000",
			2523 => "0000001110000000000111010100000100",
			2524 => "11111111110000110010011110101101",
			2525 => "00000000000000000010011110101101",
			2526 => "0000000101000000001100100100010000",
			2527 => "0000000010000000001101101100001100",
			2528 => "0000001110000000000010000000000100",
			2529 => "00000000000000000010011110101101",
			2530 => "0000000010000000000110010000000100",
			2531 => "00000000000000000010011110101101",
			2532 => "00000000010101110010011110101101",
			2533 => "00000000000000000010011110101101",
			2534 => "0000000111000000001000011000000100",
			2535 => "11111111111011010010011110101101",
			2536 => "0000000111000000000101100100000100",
			2537 => "00000000000110100010011110101101",
			2538 => "00000000000000000010011110101101",
			2539 => "0000000000000000001100000100010000",
			2540 => "0000001001000000000101010000001100",
			2541 => "0000000100000000000110111100001000",
			2542 => "0000001011000000001001110100000100",
			2543 => "00000000000000000010100000000001",
			2544 => "00000000001011010010100000000001",
			2545 => "00000000000000000010100000000001",
			2546 => "00000000000000000010100000000001",
			2547 => "0000001001000000000111101100001100",
			2548 => "0000001011000000001011110100001000",
			2549 => "0000001011000000000000011100000100",
			2550 => "00000000000000000010100000000001",
			2551 => "11111111101010100010100000000001",
			2552 => "00000000000000000010100000000001",
			2553 => "0000000000000000000001110100001100",
			2554 => "0000001011000000000101100100000100",
			2555 => "00000000000000000010100000000001",
			2556 => "0000001011000000001011110100000100",
			2557 => "00000000010000000010100000000001",
			2558 => "00000000000000000010100000000001",
			2559 => "00000000000000000010100000000001",
			2560 => "0000000100000000000001011100011000",
			2561 => "0000001001000000000100111100000100",
			2562 => "00000000000000000010100000111101",
			2563 => "0000000001000000001101111100010000",
			2564 => "0000000111000000000110100100000100",
			2565 => "00000000000000000010100000111101",
			2566 => "0000001011000000000100000100000100",
			2567 => "00000000000000000010100000111101",
			2568 => "0000001010000000000111110100000100",
			2569 => "00000000011111100010100000111101",
			2570 => "00000000000000000010100000111101",
			2571 => "00000000000000000010100000111101",
			2572 => "0000001001000000001010100000000100",
			2573 => "11111111111101010010100000111101",
			2574 => "00000000000000000010100000111101",
			2575 => "0000001110000000001100000000001000",
			2576 => "0000001101000000001001010100000100",
			2577 => "00000000000000000010100001111001",
			2578 => "11111111111110110010100001111001",
			2579 => "0000001101000000000011001000010100",
			2580 => "0000001001000000000100111100000100",
			2581 => "00000000000000000010100001111001",
			2582 => "0000001110000000000010010100001100",
			2583 => "0000001101000000001110000100000100",
			2584 => "00000000000000000010100001111001",
			2585 => "0000001001000000000010101100000100",
			2586 => "00000000001011100010100001111001",
			2587 => "00000000000000000010100001111001",
			2588 => "00000000000000000010100001111001",
			2589 => "00000000000000000010100001111001",
			2590 => "0000000001000000000000111100001000",
			2591 => "0000001010000000001001100100000100",
			2592 => "00000000000000000010100010110101",
			2593 => "11111111111010100010100010110101",
			2594 => "0000001111000000001011110000010100",
			2595 => "0000000001000000001100011000010000",
			2596 => "0000001001000000000100111100000100",
			2597 => "00000000000000000010100010110101",
			2598 => "0000001010000000001010100000000100",
			2599 => "00000000000000000010100010110101",
			2600 => "0000001010000000001001000100000100",
			2601 => "00000000001010010010100010110101",
			2602 => "00000000000000000010100010110101",
			2603 => "00000000000000000010100010110101",
			2604 => "00000000000000000010100010110101",
			2605 => "0000000110000000001001100100011100",
			2606 => "0000000100000000000110101100010000",
			2607 => "0000001100000000001011000000001000",
			2608 => "0000001100000000001010111000000100",
			2609 => "00000000000000000010100100010001",
			2610 => "00000000010010110010100100010001",
			2611 => "0000001100000000001001110100000100",
			2612 => "11111111110001100010100100010001",
			2613 => "00000000000000000010100100010001",
			2614 => "0000001011000000001011110100001000",
			2615 => "0000001010000000001010100000000100",
			2616 => "00000000000000000010100100010001",
			2617 => "11111111011011110010100100010001",
			2618 => "00000000000000000010100100010001",
			2619 => "0000000000000000000001110100010000",
			2620 => "0000000101000000000101110000001100",
			2621 => "0000001100000000001010111000000100",
			2622 => "00000000000000000010100100010001",
			2623 => "0000001110000000001010000100000100",
			2624 => "00000000000000000010100100010001",
			2625 => "00000000100100110010100100010001",
			2626 => "00000000000000000010100100010001",
			2627 => "00000000000000000010100100010001",
			2628 => "0000000100000000000001011100011000",
			2629 => "0000000011000000001000100000010100",
			2630 => "0000001100000000001010111000000100",
			2631 => "00000000000000000010100101000101",
			2632 => "0000001100000000001001001000001100",
			2633 => "0000000111000000001000011000001000",
			2634 => "0000000000000000001001101000000100",
			2635 => "00000000011011010010100101000101",
			2636 => "00000000000000000010100101000101",
			2637 => "00000000000000000010100101000101",
			2638 => "00000000000000000010100101000101",
			2639 => "00000000000000000010100101000101",
			2640 => "00000000000000000010100101000101",
			2641 => "0000000000000000000010101000011100",
			2642 => "0000001110000000001100000000001000",
			2643 => "0000000100000000001100010000000100",
			2644 => "00000000000000000010100110000001",
			2645 => "11111111111101000010100110000001",
			2646 => "0000001101000000001001010000000100",
			2647 => "00000000000000000010100110000001",
			2648 => "0000000101000000001001010000001100",
			2649 => "0000001100000000001010111000000100",
			2650 => "00000000000000000010100110000001",
			2651 => "0000001001000000000100111100000100",
			2652 => "00000000000000000010100110000001",
			2653 => "00000000100101000010100110000001",
			2654 => "00000000000000000010100110000001",
			2655 => "00000000000000000010100110000001",
			2656 => "0000001111000000001100000000001100",
			2657 => "0000001000000000001000100100001000",
			2658 => "0000000111000000000110100100000100",
			2659 => "00000000000000000010100111011101",
			2660 => "11111111100101100010100111011101",
			2661 => "00000000000000000010100111011101",
			2662 => "0000001100000000001000000000010000",
			2663 => "0000001010000000000010101100001000",
			2664 => "0000000110000000001101111100000100",
			2665 => "00000000000000000010100111011101",
			2666 => "11111111111000110010100111011101",
			2667 => "0000001010000000001000100100000100",
			2668 => "00000000000100100010100111011101",
			2669 => "00000000000000000010100111011101",
			2670 => "0000001100000000000110100100010000",
			2671 => "0000001101000000001100010100001100",
			2672 => "0000001110000000001110110100000100",
			2673 => "00000000000000000010100111011101",
			2674 => "0000001010000000001001000100000100",
			2675 => "00000000100011110010100111011101",
			2676 => "00000000000000000010100111011101",
			2677 => "00000000000000000010100111011101",
			2678 => "00000000000000000010100111011101",
			2679 => "0000000100000000001011101100100100",
			2680 => "0000001100000000001011000000010000",
			2681 => "0000001100000000000100011000000100",
			2682 => "00000000000000000010101001001001",
			2683 => "0000001010000000000111101100000100",
			2684 => "00000000000000000010101001001001",
			2685 => "0000001011000000000100000100000100",
			2686 => "00000000000000000010101001001001",
			2687 => "00000000011010000010101001001001",
			2688 => "0000001011000000000100010000010000",
			2689 => "0000000000000000001001101000001100",
			2690 => "0000001100000000001001110100001000",
			2691 => "0000000010000000000010000000000100",
			2692 => "00000000000000000010101001001001",
			2693 => "11111111100111100010101001001001",
			2694 => "00000000000000000010101001001001",
			2695 => "00000000000000000010101001001001",
			2696 => "00000000001010100010101001001001",
			2697 => "0000000010000000001000100000001100",
			2698 => "0000000000000000001011010100000100",
			2699 => "00000000000000000010101001001001",
			2700 => "0000001011000000000101100100000100",
			2701 => "00000000000000000010101001001001",
			2702 => "11111111101000100010101001001001",
			2703 => "0000000010000000001101101100000100",
			2704 => "00000000000001000010101001001001",
			2705 => "00000000000000000010101001001001",
			2706 => "0000000100000000000001011100100000",
			2707 => "0000001000000000001000100100001000",
			2708 => "0000000001000000001001011000000100",
			2709 => "00000000000000000010101010011101",
			2710 => "11111111111111110010101010011101",
			2711 => "0000000111000000000110100100000100",
			2712 => "00000000000000000010101010011101",
			2713 => "0000000110000000000100110100000100",
			2714 => "00000000000000000010101010011101",
			2715 => "0000001100000000000001101000001100",
			2716 => "0000000110000000001101011000001000",
			2717 => "0000000000000000001001101000000100",
			2718 => "00000000100010010010101010011101",
			2719 => "00000000000000000010101010011101",
			2720 => "00000000000000000010101010011101",
			2721 => "00000000000000000010101010011101",
			2722 => "0000000110000000001000010000001000",
			2723 => "0000001100000000001000011000000100",
			2724 => "11111111101001100010101010011101",
			2725 => "00000000000000000010101010011101",
			2726 => "00000000000000000010101010011101",
			2727 => "0000000100000000000001011100011100",
			2728 => "0000001010000000000000001000000100",
			2729 => "00000000000000000010101011101001",
			2730 => "0000001100000000000100011000000100",
			2731 => "00000000000000000010101011101001",
			2732 => "0000001100000000000001101000010000",
			2733 => "0000001110000000000010000000000100",
			2734 => "00000000000000000010101011101001",
			2735 => "0000001001000000001111000000000100",
			2736 => "00000000000000000010101011101001",
			2737 => "0000001101000000000001000000000100",
			2738 => "00000000000000000010101011101001",
			2739 => "00000000011110100010101011101001",
			2740 => "00000000000000000010101011101001",
			2741 => "0000000110000000000100111100001000",
			2742 => "0000001100000000000001011000000100",
			2743 => "11111111101111000010101011101001",
			2744 => "00000000000000000010101011101001",
			2745 => "00000000000000000010101011101001",
			2746 => "0000001100000000001001110100011100",
			2747 => "0000001001000000001010100000011000",
			2748 => "0000001011000000000000011100000100",
			2749 => "00000000000000000010101100101101",
			2750 => "0000000001000000001001011000000100",
			2751 => "00000000000000000010101100101101",
			2752 => "0000001111000000001001100000000100",
			2753 => "00000000000000000010101100101101",
			2754 => "0000001000000000001100011100001000",
			2755 => "0000000111000000001001001000000100",
			2756 => "00000000000000000010101100101101",
			2757 => "11111111101001000010101100101101",
			2758 => "00000000000000000010101100101101",
			2759 => "00000000000000000010101100101101",
			2760 => "0000001100000000000110100100000100",
			2761 => "00000000000000010010101100101101",
			2762 => "00000000000000000010101100101101",
			2763 => "0000001001000000001010100000100100",
			2764 => "0000001011000000000101100100010100",
			2765 => "0000001011000000001001110100000100",
			2766 => "00000000000000000010101110011001",
			2767 => "0000000001000000001101111100001100",
			2768 => "0000001111000000001011101100001000",
			2769 => "0000001110000000001110101100000100",
			2770 => "00000000000000000010101110011001",
			2771 => "00000000000111010010101110011001",
			2772 => "00000000000000000010101110011001",
			2773 => "00000000000000000010101110011001",
			2774 => "0000001011000000000110110100001100",
			2775 => "0000001111000000001001100000000100",
			2776 => "00000000000000000010101110011001",
			2777 => "0000001110000000001000001100000100",
			2778 => "11111111101001110010101110011001",
			2779 => "00000000000000000010101110011001",
			2780 => "00000000000000000010101110011001",
			2781 => "0000001011000000001010010100010000",
			2782 => "0000000101000000001110101000000100",
			2783 => "00000000000000000010101110011001",
			2784 => "0000001111000000001110000000001000",
			2785 => "0000000010000000001011110000000100",
			2786 => "00000000010100010010101110011001",
			2787 => "00000000000000000010101110011001",
			2788 => "00000000000000000010101110011001",
			2789 => "00000000000000000010101110011001",
			2790 => "0000000101000000001111010000100100",
			2791 => "0000000101000000001101000100001100",
			2792 => "0000000000000000000001010100000100",
			2793 => "00000000000000000010101111111101",
			2794 => "0000000110000000001011001100000100",
			2795 => "11111111101101000010101111111101",
			2796 => "00000000000000000010101111111101",
			2797 => "0000001100000000001001001000010100",
			2798 => "0000000110000000000100110100000100",
			2799 => "00000000000000000010101111111101",
			2800 => "0000000010000000001101101100001100",
			2801 => "0000001000000000001000100100000100",
			2802 => "00000000000000000010101111111101",
			2803 => "0000001010000000001000100100000100",
			2804 => "00000000101001100010101111111101",
			2805 => "00000000000000000010101111111101",
			2806 => "00000000000000000010101111111101",
			2807 => "00000000000000000010101111111101",
			2808 => "0000001011000000001011110100001100",
			2809 => "0000001110000000000001011100001000",
			2810 => "0000000011000000001000100000000100",
			2811 => "00000000000000000010101111111101",
			2812 => "11111111101001100010101111111101",
			2813 => "00000000000000000010101111111101",
			2814 => "00000000000000000010101111111101",
			2815 => "0000001101000000000101110000011100",
			2816 => "0000000000000000001111001000010100",
			2817 => "0000001001000000001111000000000100",
			2818 => "00000000000000000010110001111001",
			2819 => "0000000111000000000110100100000100",
			2820 => "00000000000000000010110001111001",
			2821 => "0000001011000000000110110100001000",
			2822 => "0000001101000000000001000000000100",
			2823 => "00000000000000000010110001111001",
			2824 => "00000000110101100010110001111001",
			2825 => "00000000000000000010110001111001",
			2826 => "0000001101000000000101110000000100",
			2827 => "11111111111010110010110001111001",
			2828 => "00000000000000000010110001111001",
			2829 => "0000000110000000001100011000010000",
			2830 => "0000001010000000000000001000000100",
			2831 => "00000000000000000010110001111001",
			2832 => "0000001011000000000110110100000100",
			2833 => "00000000000000000010110001111001",
			2834 => "0000000010000000000110111100000100",
			2835 => "00000000010011000010110001111001",
			2836 => "00000000000000000010110001111001",
			2837 => "0000001010000000000011101000001000",
			2838 => "0000000111000000001111011100000100",
			2839 => "11111111011110010010110001111001",
			2840 => "00000000000000000010110001111001",
			2841 => "0000000000000000000001110100001000",
			2842 => "0000000010000000001000101000000100",
			2843 => "00000000001001100010110001111001",
			2844 => "00000000000000000010110001111001",
			2845 => "00000000000000000010110001111001",
			2846 => "0000000100000000001100010000000100",
			2847 => "00000000000000000010110010110101",
			2848 => "0000001011000000000110110100011000",
			2849 => "0000001110000000001100111000010100",
			2850 => "0000001011000000000101100100000100",
			2851 => "00000000000000000010110010110101",
			2852 => "0000000111000000001001001000000100",
			2853 => "00000000000000000010110010110101",
			2854 => "0000000101000000000101001000001000",
			2855 => "0000000111000000001000011000000100",
			2856 => "11111111100110100010110010110101",
			2857 => "00000000000000000010110010110101",
			2858 => "00000000000000000010110010110101",
			2859 => "00000000000000000010110010110101",
			2860 => "00000000000000000010110010110101",
			2861 => "0000001001000000001111000000000100",
			2862 => "00000000000000000010110011110001",
			2863 => "0000000000000000001010101100011000",
			2864 => "0000001100000000000100011000000100",
			2865 => "00000000000000000010110011110001",
			2866 => "0000000101000000001110010000010000",
			2867 => "0000001010000000000000001000000100",
			2868 => "00000000000000000010110011110001",
			2869 => "0000000001000000001010011000001000",
			2870 => "0000001011000000000100000100000100",
			2871 => "00000000000000000010110011110001",
			2872 => "00000000010010100010110011110001",
			2873 => "00000000000000000010110011110001",
			2874 => "00000000000000000010110011110001",
			2875 => "00000000000000000010110011110001",
			2876 => "0000000000000000000010101000011100",
			2877 => "0000001100000000001101010100000100",
			2878 => "00000000000000000010110100101101",
			2879 => "0000001001000000001111000000000100",
			2880 => "00000000000000000010110100101101",
			2881 => "0000000111000000000110100100000100",
			2882 => "00000000000000000010110100101101",
			2883 => "0000000010000000001110110100000100",
			2884 => "00000000000000000010110100101101",
			2885 => "0000000001000000001010011000001000",
			2886 => "0000000011000000000010010100000100",
			2887 => "00000000010110000010110100101101",
			2888 => "00000000000000000010110100101101",
			2889 => "00000000000000000010110100101101",
			2890 => "00000000000000000010110100101101",
			2891 => "0000000100000000001100010000000100",
			2892 => "00000000000000000010110101111001",
			2893 => "0000000101000000001111010000011100",
			2894 => "0000001110000000000111010100010100",
			2895 => "0000001011000000000100010000010000",
			2896 => "0000001011000000000000011100000100",
			2897 => "00000000000000000010110101111001",
			2898 => "0000001100000000001010111000000100",
			2899 => "00000000000000000010110101111001",
			2900 => "0000000011000000000000010000000100",
			2901 => "11111111100011000010110101111001",
			2902 => "00000000000000000010110101111001",
			2903 => "00000000000000000010110101111001",
			2904 => "0000001010000000001000100100000100",
			2905 => "00000000000111000010110101111001",
			2906 => "00000000000000000010110101111001",
			2907 => "0000000011000000001000001100000100",
			2908 => "00000000000000100010110101111001",
			2909 => "00000000000000000010110101111001",
			2910 => "0000000000000000001001101000011100",
			2911 => "0000000001000000001011111100010000",
			2912 => "0000000111000000001011000000000100",
			2913 => "00000000000000000010111000000101",
			2914 => "0000001111000000001111010100001000",
			2915 => "0000000011000000000111010100000100",
			2916 => "00000000011110100010111000000101",
			2917 => "00000000000000000010111000000101",
			2918 => "00000000000000000010111000000101",
			2919 => "0000001010000000000010101100001000",
			2920 => "0000000111000000001001001000000100",
			2921 => "00000000000000000010111000000101",
			2922 => "11111111100111110010111000000101",
			2923 => "00000000000000000010111000000101",
			2924 => "0000001001000000000111101100010000",
			2925 => "0000000111000000000110110100001100",
			2926 => "0000000100000000001000100000001000",
			2927 => "0000000100000000000110101100000100",
			2928 => "11111111111111100010111000000101",
			2929 => "00000000000000000010111000000101",
			2930 => "11111111010000110010111000000101",
			2931 => "00000000000000000010111000000101",
			2932 => "0000001101000000000010011100010000",
			2933 => "0000000101000000000110100000000100",
			2934 => "00000000000000000010111000000101",
			2935 => "0000001110000000001010000100000100",
			2936 => "00000000000000000010111000000101",
			2937 => "0000000101000000001100100100000100",
			2938 => "11111111110110010010111000000101",
			2939 => "00000000000000000010111000000101",
			2940 => "0000001101000000001100010100001000",
			2941 => "0000001110000000000110111000000100",
			2942 => "00000000001111010010111000000101",
			2943 => "00000000000000000010111000000101",
			2944 => "00000000000000000010111000000101",
			2945 => "0000001100000000001011000000101000",
			2946 => "0000000100000000001100010000001000",
			2947 => "0000000001000000001101101000000100",
			2948 => "00000000000000000010111010000001",
			2949 => "00000000000001110010111010000001",
			2950 => "0000001001000000000100101100010000",
			2951 => "0000000111000000001000011000001100",
			2952 => "0000000110000000001101111100000100",
			2953 => "00000000000000000010111010000001",
			2954 => "0000001011000000000101100100000100",
			2955 => "00000000000000000010111010000001",
			2956 => "11111111100101010010111010000001",
			2957 => "00000000000000000010111010000001",
			2958 => "0000000001000000001101111100001100",
			2959 => "0000000111000000000001101000001000",
			2960 => "0000000111000000001000000000000100",
			2961 => "00000000000000000010111010000001",
			2962 => "00000000001001100010111010000001",
			2963 => "00000000000000000010111010000001",
			2964 => "00000000000000000010111010000001",
			2965 => "0000000000000000000101000100000100",
			2966 => "00000000000000000010111010000001",
			2967 => "0000000110000000001100011000001000",
			2968 => "0000001100000000001000000000000100",
			2969 => "00000000000000000010111010000001",
			2970 => "00000000100101000010111010000001",
			2971 => "0000000001000000000001000100000100",
			2972 => "11111111110011110010111010000001",
			2973 => "0000000001000000001010011000000100",
			2974 => "00000000010010010010111010000001",
			2975 => "00000000000000000010111010000001",
			2976 => "0000001110000000000111010100101100",
			2977 => "0000000000000000001100000100011100",
			2978 => "0000000011000000001010000100010100",
			2979 => "0000001001000000001111000000000100",
			2980 => "00000000000000000010111011111101",
			2981 => "0000000110000000001100011000001100",
			2982 => "0000000001000000001001011000000100",
			2983 => "00000000000000000010111011111101",
			2984 => "0000000000000000000101000100000100",
			2985 => "00000000000000000010111011111101",
			2986 => "00000000100100010010111011111101",
			2987 => "00000000000000000010111011111101",
			2988 => "0000001000000000001000010100000100",
			2989 => "11111111111111100010111011111101",
			2990 => "00000000000000000010111011111101",
			2991 => "0000000101000000000010110100000100",
			2992 => "00000000000000000010111011111101",
			2993 => "0000001101000000001110010000001000",
			2994 => "0000001011000000000000011100000100",
			2995 => "00000000000000000010111011111101",
			2996 => "11111111101011010010111011111101",
			2997 => "00000000000000000010111011111101",
			2998 => "0000000000000000000001110100010000",
			2999 => "0000000100000000001110000000001100",
			3000 => "0000001000000000000001010000000100",
			3001 => "00000000000000000010111011111101",
			3002 => "0000000001000000001100011000000100",
			3003 => "00000000011101100010111011111101",
			3004 => "00000000000000000010111011111101",
			3005 => "00000000000000000010111011111101",
			3006 => "00000000000000000010111011111101",
			3007 => "0000001100000000001011000000101100",
			3008 => "0000000100000000000110111100010000",
			3009 => "0000001100000000001010111000000100",
			3010 => "00000000000000000010111110000001",
			3011 => "0000000111000000001000011000001000",
			3012 => "0000000111000000001011000000000100",
			3013 => "00000000000000000010111110000001",
			3014 => "00000000001010100010111110000001",
			3015 => "00000000000000000010111110000001",
			3016 => "0000001001000000000111101100001100",
			3017 => "0000001011000000000000011100000100",
			3018 => "00000000000000000010111110000001",
			3019 => "0000001110000000001100010000000100",
			3020 => "00000000000000000010111110000001",
			3021 => "11111111011111010010111110000001",
			3022 => "0000000001000000001101111100001100",
			3023 => "0000001110000000001111010100000100",
			3024 => "00000000000000000010111110000001",
			3025 => "0000001010000000001000100100000100",
			3026 => "00000000001110010010111110000001",
			3027 => "00000000000000000010111110000001",
			3028 => "00000000000000000010111110000001",
			3029 => "0000001110000000001100000000000100",
			3030 => "00000000000000000010111110000001",
			3031 => "0000000001000000001100011000010000",
			3032 => "0000000001000000000000111100000100",
			3033 => "00000000000000000010111110000001",
			3034 => "0000000000000000000111000000001000",
			3035 => "0000001101000000000010000100000100",
			3036 => "00000000101100100010111110000001",
			3037 => "00000000000000000010111110000001",
			3038 => "00000000000000000010111110000001",
			3039 => "00000000000000000010111110000001",
			3040 => "0000000100000000001011101100110100",
			3041 => "0000001101000000000101110000011000",
			3042 => "0000000111000000000110100100000100",
			3043 => "00000000000000000011000000010101",
			3044 => "0000001001000000001111000000000100",
			3045 => "00000000000000000011000000010101",
			3046 => "0000001011000000000110110100001100",
			3047 => "0000001010000000000000001000000100",
			3048 => "00000000000000000011000000010101",
			3049 => "0000001101000000001110000100000100",
			3050 => "00000000000000000011000000010101",
			3051 => "00000000101011100011000000010101",
			3052 => "00000000000000000011000000010101",
			3053 => "0000001011000000000110110100001100",
			3054 => "0000000011000000000000010000001000",
			3055 => "0000001111000000001001100000000100",
			3056 => "00000000000000000011000000010101",
			3057 => "11111111110011000011000000010101",
			3058 => "00000000000000000011000000010101",
			3059 => "0000000011000000000111010100001000",
			3060 => "0000001111000000001100000000000100",
			3061 => "00000000000000000011000000010101",
			3062 => "00000000011101110011000000010101",
			3063 => "0000000010000000001010000100000100",
			3064 => "11111111111111110011000000010101",
			3065 => "00000000000000000011000000010101",
			3066 => "0000000011000000001111100100001100",
			3067 => "0000001110000000001000001100001000",
			3068 => "0000000000000000001011010100000100",
			3069 => "00000000000000000011000000010101",
			3070 => "11111111010111010011000000010101",
			3071 => "00000000000000000011000000010101",
			3072 => "0000000000000000000111000100001000",
			3073 => "0000000000000000001011010100000100",
			3074 => "00000000000000000011000000010101",
			3075 => "00000000010110110011000000010101",
			3076 => "00000000000000000011000000010101",
			3077 => "0000000000000000001001101000100000",
			3078 => "0000001101000000000101001000001100",
			3079 => "0000000001000000001011111100001000",
			3080 => "0000000001000000001101101000000100",
			3081 => "00000000000000000011000010101001",
			3082 => "00000000000010000011000010101001",
			3083 => "11111111110110010011000010101001",
			3084 => "0000000101000000000101001000010000",
			3085 => "0000001111000000001110110100000100",
			3086 => "00000000000000000011000010101001",
			3087 => "0000001001000000001111000000000100",
			3088 => "00000000000000000011000010101001",
			3089 => "0000001110000000000110111100000100",
			3090 => "00000000110001000011000010101001",
			3091 => "00000000000000000011000010101001",
			3092 => "00000000000000000011000010101001",
			3093 => "0000000001000000000111101000001100",
			3094 => "0000001011000000001010010100001000",
			3095 => "0000000100000000000000010000000100",
			3096 => "00000000000000000011000010101001",
			3097 => "11111111001101000011000010101001",
			3098 => "00000000000000000011000010101001",
			3099 => "0000000101000000001100100100001100",
			3100 => "0000000001000000001101111100000100",
			3101 => "00000000000000000011000010101001",
			3102 => "0000000111000000000001101000000100",
			3103 => "11111111011111100011000010101001",
			3104 => "00000000000000000011000010101001",
			3105 => "0000001101000000001100010100010000",
			3106 => "0000000001000000001010011000001100",
			3107 => "0000001011000000001011011100000100",
			3108 => "00000000000000000011000010101001",
			3109 => "0000000000000000001010101100000100",
			3110 => "00000000101001010011000010101001",
			3111 => "00000000000000000011000010101001",
			3112 => "00000000000000000011000010101001",
			3113 => "00000000000000000011000010101001",
			3114 => "0000000000000000000111000100110100",
			3115 => "0000001001000000000111101100101000",
			3116 => "0000000010000000001010000100011100",
			3117 => "0000001000000000001001000100010100",
			3118 => "0000000001000000000101011100001100",
			3119 => "0000001001000000000100111100001000",
			3120 => "0000000111000000000001101000000100",
			3121 => "11111111111110010011000100011101",
			3122 => "00000000000000000011000100011101",
			3123 => "00000000100010100011000100011101",
			3124 => "0000000111000000000001101000000100",
			3125 => "11111111010100100011000100011101",
			3126 => "00000000000000000011000100011101",
			3127 => "0000001101000000001111010000000100",
			3128 => "00000000000000000011000100011101",
			3129 => "00000000111010010011000100011101",
			3130 => "0000001011000000001011110100001000",
			3131 => "0000001001000000000100101100000100",
			3132 => "11111111001100110011000100011101",
			3133 => "00000000000000000011000100011101",
			3134 => "00000000000100100011000100011101",
			3135 => "0000000010000000001000001100000100",
			3136 => "00000000000000000011000100011101",
			3137 => "0000000011000000001000001100000100",
			3138 => "00000000000000000011000100011101",
			3139 => "00000000110011000011000100011101",
			3140 => "0000001110000000000001011100000100",
			3141 => "11111111001000110011000100011101",
			3142 => "00000000000000000011000100011101",
			3143 => "0000001110000000000111010100110100",
			3144 => "0000000000000000001100000100011100",
			3145 => "0000000011000000001010000100010100",
			3146 => "0000001001000000001111000000000100",
			3147 => "00000000000000000011000110100001",
			3148 => "0000000110000000001100011000001100",
			3149 => "0000000001000000001001011000000100",
			3150 => "00000000000000000011000110100001",
			3151 => "0000000000000000000101000100000100",
			3152 => "00000000000000000011000110100001",
			3153 => "00000000100111100011000110100001",
			3154 => "00000000000000000011000110100001",
			3155 => "0000001000000000001000010100000100",
			3156 => "11111111111110000011000110100001",
			3157 => "00000000000000000011000110100001",
			3158 => "0000000101000000000010110100000100",
			3159 => "00000000000000000011000110100001",
			3160 => "0000000111000000001001001000000100",
			3161 => "00000000000000000011000110100001",
			3162 => "0000001011000000000101110100001100",
			3163 => "0000001011000000000000011100000100",
			3164 => "00000000000000000011000110100001",
			3165 => "0000000111000000001111011100000100",
			3166 => "11111111100110000011000110100001",
			3167 => "00000000000000000011000110100001",
			3168 => "00000000000000000011000110100001",
			3169 => "0000000000000000000001110100001100",
			3170 => "0000000001000000001110010100000100",
			3171 => "00000000000000000011000110100001",
			3172 => "0000000001000000001100011000000100",
			3173 => "00000000011100100011000110100001",
			3174 => "00000000000000000011000110100001",
			3175 => "00000000000000000011000110100001",
			3176 => "0000000100000000000110111000110000",
			3177 => "0000001001000000001111000000010000",
			3178 => "0000000111000000001000011000001100",
			3179 => "0000001010000000001001100100001000",
			3180 => "0000001100000000000000001100000100",
			3181 => "11111110011101000011001001000101",
			3182 => "00000101110101100011001001000101",
			3183 => "11111110011000100011001001000101",
			3184 => "00000000011101000011001001000101",
			3185 => "0000001101000000001110000100001000",
			3186 => "0000001000000000000110011000000100",
			3187 => "00000001001001010011001001000101",
			3188 => "11111110011011010011001001000101",
			3189 => "0000000011000000001000101000010000",
			3190 => "0000000001000000001001011000000100",
			3191 => "11111111100111110011001001000101",
			3192 => "0000001010000000001000100100001000",
			3193 => "0000001010000000000000001000000100",
			3194 => "00000001101100100011001001000101",
			3195 => "00000010010101010011001001000101",
			3196 => "11111110111010000011001001000101",
			3197 => "0000000100000000000010010100000100",
			3198 => "11111110111101100011001001000101",
			3199 => "00000001010000110011001001000101",
			3200 => "0000000100000000001000110100011000",
			3201 => "0000000111000000000001101000000100",
			3202 => "11111110010111010011001001000101",
			3203 => "0000001101000000001100010100010000",
			3204 => "0000000101000000000101001000001000",
			3205 => "0000001101000000000100101000000100",
			3206 => "11111110101010010011001001000101",
			3207 => "00000001110100110011001001000101",
			3208 => "0000001111000000000010010100000100",
			3209 => "00000011010100110011001001000101",
			3210 => "00000101101000010011001001000101",
			3211 => "11111110011000110011001001000101",
			3212 => "0000000100000000000101000000001000",
			3213 => "0000000100000000000101000000000100",
			3214 => "11111110011101010011001001000101",
			3215 => "11111111011100010011001001000101",
			3216 => "11111110011000000011001001000101",
			3217 => "0000000000000000000010101000111000",
			3218 => "0000001001000000001001100100001100",
			3219 => "0000000110000000000000111100001000",
			3220 => "0000000010000000000111010000000100",
			3221 => "11111110100111000011001011001001",
			3222 => "00000001101111110011001011001001",
			3223 => "11111110011010000011001011001001",
			3224 => "0000001101000000001100010100100100",
			3225 => "0000000101000000000110100000001100",
			3226 => "0000000001000000001011111100001000",
			3227 => "0000001100000000001010111000000100",
			3228 => "11111111111110000011001011001001",
			3229 => "00000001101011110011001011001001",
			3230 => "11111110010000010011001011001001",
			3231 => "0000000110000000000100111100010000",
			3232 => "0000000000000000001111001000001000",
			3233 => "0000000001000000000000111100000100",
			3234 => "00000000011111000011001011001001",
			3235 => "00000001100101110011001011001001",
			3236 => "0000000011000000001111100100000100",
			3237 => "11111101100101000011001011001001",
			3238 => "00000001100111110011001011001001",
			3239 => "0000000010000000001000101000000100",
			3240 => "00000010010100000011001011001001",
			3241 => "00000011100111000011001011001001",
			3242 => "0000000010000000001100111000000100",
			3243 => "00000000011001110011001011001001",
			3244 => "11111110011011010011001011001001",
			3245 => "0000000000000000001010101100001000",
			3246 => "0000000110000000001000010000000100",
			3247 => "11111110011011110011001011001001",
			3248 => "00000001011010010011001011001001",
			3249 => "11111110011001000011001011001001",
			3250 => "0000000000000000000010101000111100",
			3251 => "0000000001000000001001011000010000",
			3252 => "0000001011000000000010001000001100",
			3253 => "0000000110000000000000111100001000",
			3254 => "0000000000000000000011101000000100",
			3255 => "11111110100011100011001101010101",
			3256 => "00000001110100010011001101010101",
			3257 => "11111110011001100011001101010101",
			3258 => "00000000000000000011001101010101",
			3259 => "0000001101000000001100010100100100",
			3260 => "0000000101000000000110100000001100",
			3261 => "0000000001000000001011111100001000",
			3262 => "0000001100000000001010111000000100",
			3263 => "00000000000000000011001101010101",
			3264 => "00000001110000110011001101010101",
			3265 => "11111110001111100011001101010101",
			3266 => "0000000110000000000100111100010000",
			3267 => "0000001010000000000000001000001000",
			3268 => "0000000011000000001110110100000100",
			3269 => "00000001010011100011001101010101",
			3270 => "11111110010111000011001101010101",
			3271 => "0000000000000000001111001000000100",
			3272 => "00000001101101110011001101010101",
			3273 => "00000000110010100011001101010101",
			3274 => "0000000101000000001001010000000100",
			3275 => "00000100001110100011001101010101",
			3276 => "00000010100111010011001101010101",
			3277 => "0000000010000000001100111000000100",
			3278 => "00000000011001100011001101010101",
			3279 => "11111110011000110011001101010101",
			3280 => "0000000000000000001010101100001000",
			3281 => "0000000110000000001000010000000100",
			3282 => "11111110011010100011001101010101",
			3283 => "00000001101001110011001101010101",
			3284 => "11111110011000110011001101010101",
			3285 => "0000001111000000001100000000010000",
			3286 => "0000001010000000001001100100000100",
			3287 => "00000000000000000011001111111001",
			3288 => "0000001001000000000100111100001000",
			3289 => "0000000001000000000000111100000100",
			3290 => "11111111100011010011001111111001",
			3291 => "00000000000000000011001111111001",
			3292 => "00000000000000000011001111111001",
			3293 => "0000000010000000000000010000100100",
			3294 => "0000001010000000000010101100010100",
			3295 => "0000001011000000000110110100001000",
			3296 => "0000000101000000001100100100000100",
			3297 => "00000000000000000011001111111001",
			3298 => "11111111010011000011001111111001",
			3299 => "0000001001000000001111000000000100",
			3300 => "00000000000000000011001111111001",
			3301 => "0000000001000000001001011000000100",
			3302 => "00000000000000000011001111111001",
			3303 => "00000000011101110011001111111001",
			3304 => "0000000011000000000110111100000100",
			3305 => "00000000000000000011001111111001",
			3306 => "0000001101000000001110000100000100",
			3307 => "00000000000000000011001111111001",
			3308 => "0000001010000000000111110100000100",
			3309 => "00000000111001000011001111111001",
			3310 => "00000000000000000011001111111001",
			3311 => "0000001110000000001000001100000100",
			3312 => "11111111100110100011001111111001",
			3313 => "0000001101000000001100010100010100",
			3314 => "0000000000000000000001110100001000",
			3315 => "0000000110000000001001100100000100",
			3316 => "00000000000000000011001111111001",
			3317 => "00000000011100000011001111111001",
			3318 => "0000001001000000001010100100000100",
			3319 => "11111111110110110011001111111001",
			3320 => "0000000011000000000001011100000100",
			3321 => "00000000000000000011001111111001",
			3322 => "00000000001111110011001111111001",
			3323 => "0000001011000000000001001000000100",
			3324 => "11111111111101010011001111111001",
			3325 => "00000000000000000011001111111001",
			3326 => "0000000000000000000001110100111100",
			3327 => "0000001001000000001111000000010000",
			3328 => "0000000101000000000101001000001100",
			3329 => "0000000110000000000000111100001000",
			3330 => "0000001001000000000001000100000100",
			3331 => "11111110100000010011010010011101",
			3332 => "00000010011010010011010010011101",
			3333 => "11111110011001000011010010011101",
			3334 => "11111111111101000011010010011101",
			3335 => "0000001101000000000001000000001000",
			3336 => "0000001001000000001001111100000100",
			3337 => "00000000111011010011010010011101",
			3338 => "11111110011100110011010010011101",
			3339 => "0000001101000000001100010100011100",
			3340 => "0000001010000000000000001000001100",
			3341 => "0000000011000000001100010000000100",
			3342 => "00000010001101110011010010011101",
			3343 => "0000000101000000001100100100000100",
			3344 => "00000000000000000011010010011101",
			3345 => "11111110001101100011010010011101",
			3346 => "0000001100000000001010111000001000",
			3347 => "0000000000000000000110001000000100",
			3348 => "00000001101100000011010010011101",
			3349 => "11111110001000010011010010011101",
			3350 => "0000000011000000001100111000000100",
			3351 => "00000001110110000011010010011101",
			3352 => "00000010110011010011010010011101",
			3353 => "0000000000000000001111001000000100",
			3354 => "00000000001011100011010010011101",
			3355 => "11111110011011100011010010011101",
			3356 => "0000000000000000001010101100010100",
			3357 => "0000001000000000000001010100001100",
			3358 => "0000000000000000000001110100001000",
			3359 => "0000001000000000000101000100000100",
			3360 => "11111110100111010011010010011101",
			3361 => "00000010111110100011010010011101",
			3362 => "11111110011001010011010010011101",
			3363 => "0000000110000000001000010000000100",
			3364 => "00000000000011110011010010011101",
			3365 => "00000011001110100011010010011101",
			3366 => "11111110011000010011010010011101",
			3367 => "0000000100000000001011110000110100",
			3368 => "0000000001000000001001011000001100",
			3369 => "0000000110000000000000111100001000",
			3370 => "0000001110000000001011000000000100",
			3371 => "11111110101011100011010100111001",
			3372 => "00000010011100110011010100111001",
			3373 => "11111110011011100011010100111001",
			3374 => "0000001101000000001110000100001100",
			3375 => "0000000100000000001100010000000100",
			3376 => "00000001101110110011010100111001",
			3377 => "0000000101000000001101000100000100",
			3378 => "11111110010011010011010100111001",
			3379 => "00000000001101000011010100111001",
			3380 => "0000000001000000001100011000011000",
			3381 => "0000001010000000000000001000001000",
			3382 => "0000000010000000001100010100000100",
			3383 => "00000000100111110011010100111001",
			3384 => "11111110011110010011010100111001",
			3385 => "0000000010000000001100000000001000",
			3386 => "0000000101000000001111010000000100",
			3387 => "00000001110010000011010100111001",
			3388 => "00000000011110100011010100111001",
			3389 => "0000001000000000001000010100000100",
			3390 => "11111111001111110011010100111001",
			3391 => "00000001001111000011010100111001",
			3392 => "11111110100110110011010100111001",
			3393 => "0000000001000000000100110100000100",
			3394 => "11111110011001010011010100111001",
			3395 => "0000000011000000000110111000010100",
			3396 => "0000001101000000000111111100000100",
			3397 => "11111110110110010011010100111001",
			3398 => "0000000111000000001000011000001000",
			3399 => "0000000100000000000101000000000100",
			3400 => "00000011000101110011010100111001",
			3401 => "00000000000000000011010100111001",
			3402 => "0000000110000000000101010000000100",
			3403 => "11111110111010010011010100111001",
			3404 => "00000000111100110011010100111001",
			3405 => "11111110011010110011010100111001",
			3406 => "0000000000000000001001101000101000",
			3407 => "0000001101000000000101001000001100",
			3408 => "0000000001000000001011111100001000",
			3409 => "0000000001000000001101101000000100",
			3410 => "00000000000000000011010111111101",
			3411 => "00000000000001110011010111111101",
			3412 => "11111111110110110011010111111101",
			3413 => "0000000110000000001100011000010100",
			3414 => "0000001110000000001100010000001100",
			3415 => "0000001101000000000111111100001000",
			3416 => "0000001101000000000010011100000100",
			3417 => "00000000000000000011010111111101",
			3418 => "11111111111101100011010111111101",
			3419 => "00000000100100100011010111111101",
			3420 => "0000001101000000001001011100000100",
			3421 => "11111111110000110011010111111101",
			3422 => "00000000000000000011010111111101",
			3423 => "0000000001000000000101011100000100",
			3424 => "00000000000000000011010111111101",
			3425 => "00000000110101010011010111111101",
			3426 => "0000000110000000001011001100001100",
			3427 => "0000001100000000001001110100001000",
			3428 => "0000000100000000000000010000000100",
			3429 => "00000000000000000011010111111101",
			3430 => "11111111001010010011010111111101",
			3431 => "00000000000000000011010111111101",
			3432 => "0000000111000000000001101000010000",
			3433 => "0000001011000000000000011100000100",
			3434 => "00000000000000000011010111111101",
			3435 => "0000001010000000001000010100001000",
			3436 => "0000000011000000001010000100000100",
			3437 => "00000000000000000011010111111101",
			3438 => "00000000100100000011010111111101",
			3439 => "00000000000000000011010111111101",
			3440 => "0000000011000000000001011100010000",
			3441 => "0000001010000000000011101000000100",
			3442 => "00000000000000000011010111111101",
			3443 => "0000001110000000000001011100001000",
			3444 => "0000000110000000001001100100000100",
			3445 => "00000000000000000011010111111101",
			3446 => "11111111101001100011010111111101",
			3447 => "00000000000000000011010111111101",
			3448 => "0000000100000000000101000000001100",
			3449 => "0000001101000000001100010100001000",
			3450 => "0000000101000000001110000100000100",
			3451 => "00000000000000000011010111111101",
			3452 => "00000000011011100011010111111101",
			3453 => "00000000000000000011010111111101",
			3454 => "00000000000000000011010111111101",
			3455 => "0000001100000000000100011000011100",
			3456 => "0000001110000000000111010100001000",
			3457 => "0000000000000000001001101000000100",
			3458 => "00000000000000000011011010011001",
			3459 => "11111110111101000011011010011001",
			3460 => "0000000111000000000001101000010000",
			3461 => "0000001111000000000011000000001100",
			3462 => "0000000111000000001001001000000100",
			3463 => "00000000000000000011011010011001",
			3464 => "0000000000000000000010101000000100",
			3465 => "00000000010111000011011010011001",
			3466 => "00000000000000000011011010011001",
			3467 => "00000000000000000011011010011001",
			3468 => "00000000000000000011011010011001",
			3469 => "0000000000000000000010101000110000",
			3470 => "0000001110000000001100000000011000",
			3471 => "0000001101000000000111111100010000",
			3472 => "0000000111000000000110100100000100",
			3473 => "00000000000000000011011010011001",
			3474 => "0000001011000000000000011100000100",
			3475 => "00000000000000000011011010011001",
			3476 => "0000000111000000001000011000000100",
			3477 => "11111111100000100011011010011001",
			3478 => "00000000000000000011011010011001",
			3479 => "0000000010000000001100000000000100",
			3480 => "00000000110011100011011010011001",
			3481 => "00000000000000000011011010011001",
			3482 => "0000000001000000000000111100000100",
			3483 => "00000000000000000011011010011001",
			3484 => "0000001101000000000010011100001000",
			3485 => "0000000001000000001101111100000100",
			3486 => "00000000010000100011011010011001",
			3487 => "11111111101101100011011010011001",
			3488 => "0000000101000000001110010000001000",
			3489 => "0000000001000000001100011000000100",
			3490 => "00000001000001000011011010011001",
			3491 => "00000000000000000011011010011001",
			3492 => "00000000000000000011011010011001",
			3493 => "11111111110110000011011010011001",
			3494 => "0000000000000000000010101001000000",
			3495 => "0000000011000000001100111000101100",
			3496 => "0000000000000000001111001000100100",
			3497 => "0000000110000000001011001100011100",
			3498 => "0000001111000000001111010100010000",
			3499 => "0000000000000000000001010100001000",
			3500 => "0000000101000000000111100000000100",
			3501 => "00000000011000110011011100100101",
			3502 => "11111111010000000011011100100101",
			3503 => "0000001101000000001111010000000100",
			3504 => "11111111100010010011011100100101",
			3505 => "00000000111110000011011100100101",
			3506 => "0000001011000000001011110100001000",
			3507 => "0000000001000000000001000100000100",
			3508 => "11111110111010010011011100100101",
			3509 => "11111111111001110011011100100101",
			3510 => "00000000101111100011011100100101",
			3511 => "0000000011000000001010000100000100",
			3512 => "00000000000000000011011100100101",
			3513 => "00000001011101000011011100100101",
			3514 => "0000000011000000001000100000000100",
			3515 => "11111110100010100011011100100101",
			3516 => "00000000000000000011011100100101",
			3517 => "0000000010000000001101101100000100",
			3518 => "00000001010101110011011100100101",
			3519 => "0000001000000000000101000100001000",
			3520 => "0000000100000000001110000000000100",
			3521 => "00000000000000000011011100100101",
			3522 => "11111111100001100011011100100101",
			3523 => "0000000001000000001010011000000100",
			3524 => "00000000110111100011011100100101",
			3525 => "00000000000000000011011100100101",
			3526 => "0000000001000000001100011000000100",
			3527 => "11111110100001100011011100100101",
			3528 => "00000000000000000011011100100101",
			3529 => "0000000000000000001001101000101100",
			3530 => "0000001101000000000101001000001100",
			3531 => "0000000001000000001011111100001000",
			3532 => "0000000001000000001101101000000100",
			3533 => "00000000000000000011011111110001",
			3534 => "00000000000001110011011111110001",
			3535 => "11111111110111010011011111110001",
			3536 => "0000000110000000001100011000011000",
			3537 => "0000001101000000000111111100001100",
			3538 => "0000000010000000000110010000000100",
			3539 => "00000000000000000011011111110001",
			3540 => "0000001101000000000010011100000100",
			3541 => "00000000000000000011011111110001",
			3542 => "11111111101101000011011111110001",
			3543 => "0000001010000000001010100000001000",
			3544 => "0000000001000000000000111100000100",
			3545 => "00000000101011100011011111110001",
			3546 => "00000000000000000011011111110001",
			3547 => "00000000000000000011011111110001",
			3548 => "0000000010000000001000001100000100",
			3549 => "00000000110011010011011111110001",
			3550 => "00000000000000000011011111110001",
			3551 => "0000000110000000001011001100001100",
			3552 => "0000001100000000001001110100001000",
			3553 => "0000000101000000000010110100000100",
			3554 => "00000000000000000011011111110001",
			3555 => "11111111001001010011011111110001",
			3556 => "00000000000000000011011111110001",
			3557 => "0000000111000000000001101000010000",
			3558 => "0000001011000000000000011100000100",
			3559 => "00000000000000000011011111110001",
			3560 => "0000001010000000001000010100001000",
			3561 => "0000000011000000001010000100000100",
			3562 => "00000000000000000011011111110001",
			3563 => "00000000100010010011011111110001",
			3564 => "00000000000000000011011111110001",
			3565 => "0000000111000000001000011000010000",
			3566 => "0000001001000000000000001000000100",
			3567 => "00000000000000000011011111110001",
			3568 => "0000001100000000001001110100001000",
			3569 => "0000000011000000000010010100000100",
			3570 => "11111111101000100011011111110001",
			3571 => "00000000000000000011011111110001",
			3572 => "00000000000000000011011111110001",
			3573 => "0000001101000000001100010100001100",
			3574 => "0000001001000000000111101100000100",
			3575 => "00000000000000000011011111110001",
			3576 => "0000001100000000000100011000000100",
			3577 => "00000000000000000011011111110001",
			3578 => "00000000011001100011011111110001",
			3579 => "00000000000000000011011111110001",
			3580 => "0000000101000000000001000000111000",
			3581 => "0000000010000000001000001100100100",
			3582 => "0000000000000000001001101000011000",
			3583 => "0000001010000000001010100100010000",
			3584 => "0000001011000000000101100100000100",
			3585 => "00000000000000000011100010110101",
			3586 => "0000000101000000000111100000001000",
			3587 => "0000001011000000000010001000000100",
			3588 => "11111111101000000011100010110101",
			3589 => "00000000000000000011100010110101",
			3590 => "00000000000000000011100010110101",
			3591 => "0000001101000000000101001000000100",
			3592 => "00000000000000000011100010110101",
			3593 => "00000000100111000011100010110101",
			3594 => "0000001100000000000100011000001000",
			3595 => "0000000111000000000001101000000100",
			3596 => "11111110111000010011100010110101",
			3597 => "00000000000000000011100010110101",
			3598 => "00000000000000000011100010110101",
			3599 => "0000000100000000000001011100000100",
			3600 => "00000000010111010011100010110101",
			3601 => "0000000100000000001011110000001100",
			3602 => "0000000111000000001000011000001000",
			3603 => "0000001100000000001010111000000100",
			3604 => "00000000000000000011100010110101",
			3605 => "11111111100010100011100010110101",
			3606 => "00000000000000000011100010110101",
			3607 => "00000000000000000011100010110101",
			3608 => "0000000000000000000010101000100100",
			3609 => "0000001010000000000000001000000100",
			3610 => "00000000000000000011100010110101",
			3611 => "0000001101000000001010001000001100",
			3612 => "0000001001000000001111000000000100",
			3613 => "00000000000000000011100010110101",
			3614 => "0000001100000000000100011000000100",
			3615 => "00000000000000000011100010110101",
			3616 => "00000000111101000011100010110101",
			3617 => "0000001100000000001001110100001000",
			3618 => "0000001001000000000100111100000100",
			3619 => "11111111111011010011100010110101",
			3620 => "00000000000000000011100010110101",
			3621 => "0000000010000000000001011100001000",
			3622 => "0000001001000000001010100100000100",
			3623 => "00000000010101110011100010110101",
			3624 => "00000000000000000011100010110101",
			3625 => "00000000000000000011100010110101",
			3626 => "0000001100000000001000000000000100",
			3627 => "00000000000000000011100010110101",
			3628 => "11111111111000110011100010110101",
			3629 => "0000001001000000001001100100001100",
			3630 => "0000001010000000001001100100001000",
			3631 => "0000000100000000000111010000000100",
			3632 => "00000000000000000011100101100001",
			3633 => "00000000000101110011100101100001",
			3634 => "11111110011011100011100101100001",
			3635 => "0000000100000000001100010000010000",
			3636 => "0000000011000000001100000000001100",
			3637 => "0000000001000000001001011000000100",
			3638 => "00000000000000000011100101100001",
			3639 => "0000001001000000001111000000000100",
			3640 => "00000000000000000011100101100001",
			3641 => "00000001101110010011100101100001",
			3642 => "11111111110001010011100101100001",
			3643 => "0000001110000000001100111000100100",
			3644 => "0000001100000000001001110100011000",
			3645 => "0000001101000000001010001000001100",
			3646 => "0000000011000000001100111000001000",
			3647 => "0000001001000000001010100000000100",
			3648 => "11111111111101100011100101100001",
			3649 => "11111110110111010011100101100001",
			3650 => "00000001011101100011100101100001",
			3651 => "0000000011000000001000100000001000",
			3652 => "0000000010000000001111010100000100",
			3653 => "11111111011011010011100101100001",
			3654 => "00000000011100110011100101100001",
			3655 => "11111110011111000011100101100001",
			3656 => "0000000100000000001011110000001000",
			3657 => "0000000001000000000000111100000100",
			3658 => "11111111110001000011100101100001",
			3659 => "00000001011100000011100101100001",
			3660 => "11111111011100000011100101100001",
			3661 => "0000001101000000001100010100010000",
			3662 => "0000001010000000001001000100001000",
			3663 => "0000001011000000001011011100000100",
			3664 => "00000000000000000011100101100001",
			3665 => "00000001101100110011100101100001",
			3666 => "0000001101000000000011001000000100",
			3667 => "11111111110011100011100101100001",
			3668 => "00000000000000000011100101100001",
			3669 => "0000001011000000001010010100000100",
			3670 => "00000000000000000011100101100001",
			3671 => "11111110110111000011100101100001",
			3672 => "0000000000000000000111000101001000",
			3673 => "0000000110000000001101011000110000",
			3674 => "0000000001000000001011111100100100",
			3675 => "0000001111000000001111010100010100",
			3676 => "0000001001000000000100111100010000",
			3677 => "0000001011000000000010001000001000",
			3678 => "0000000011000000001100000000000100",
			3679 => "00000000000000000011100111111101",
			3680 => "11111111110011110011100111111101",
			3681 => "0000000010000000001110110100000100",
			3682 => "00000000000000000011100111111101",
			3683 => "00000000011000000011100111111101",
			3684 => "00000000101101110011100111111101",
			3685 => "0000001011000000001011110100001100",
			3686 => "0000000001000000000001000100001000",
			3687 => "0000001100000000000100011000000100",
			3688 => "00000000000000000011100111111101",
			3689 => "11111111010111000011100111111101",
			3690 => "00000000000000000011100111111101",
			3691 => "00000000000000000011100111111101",
			3692 => "0000001010000000000010101100001000",
			3693 => "0000000111000000001001001000000100",
			3694 => "00000000000000000011100111111101",
			3695 => "11111111001101100011100111111101",
			3696 => "00000000000000000011100111111101",
			3697 => "0000001001000000001001111100000100",
			3698 => "00000000000000000011100111111101",
			3699 => "0000001100000000000100011000001100",
			3700 => "0000000111000000000110100100001000",
			3701 => "0000000111000000001001001000000100",
			3702 => "00000000000000000011100111111101",
			3703 => "00000000000010110011100111111101",
			3704 => "00000000000000000011100111111101",
			3705 => "0000000011000000000110111100000100",
			3706 => "00000000000000000011100111111101",
			3707 => "00000001000111010011100111111101",
			3708 => "0000001110000000000001011100000100",
			3709 => "11111111000101100011100111111101",
			3710 => "00000000000000000011100111111101",
			3711 => "0000000000000000000001110101001000",
			3712 => "0000000001000000001001011000100000",
			3713 => "0000000001000000001001011000010000",
			3714 => "0000001010000000001001100100001000",
			3715 => "0000000111000000000001111100000100",
			3716 => "11111110011011100011101011011001",
			3717 => "00001101011110100011101011011001",
			3718 => "0000000111000000001000011000000100",
			3719 => "11111110011000000011101011011001",
			3720 => "11111111011010110011101011011001",
			3721 => "0000001101000000000010011100001000",
			3722 => "0000001011000000000101100100000100",
			3723 => "11111111000010000011101011011001",
			3724 => "00000111100110010011101011011001",
			3725 => "0000001011000000000110110100000100",
			3726 => "11111110011100010011101011011001",
			3727 => "00000000000000000011101011011001",
			3728 => "0000001101000000001110000100001000",
			3729 => "0000000010000000000110010000000100",
			3730 => "00000001100101010011101011011001",
			3731 => "11111110011010000011101011011001",
			3732 => "0000001101000000000110010000011000",
			3733 => "0000001010000000000000001000001100",
			3734 => "0000000011000000001100010000000100",
			3735 => "00000010111111000011101011011001",
			3736 => "0000001100000000001000000000000100",
			3737 => "11111110010100000011101011011001",
			3738 => "00000000001011000011101011011001",
			3739 => "0000001100000000000111001000000100",
			3740 => "11111111111000100011101011011001",
			3741 => "0000000101000000000110100000000100",
			3742 => "00000001100101010011101011011001",
			3743 => "00000011000001000011101011011001",
			3744 => "0000000000000000000111000100000100",
			3745 => "00000000001000000011101011011001",
			3746 => "11111110100001110011101011011001",
			3747 => "0000000000000000001010101100100100",
			3748 => "0000001000000000000001010100011000",
			3749 => "0000001000000000000001010100010000",
			3750 => "0000000000000000000001110100001100",
			3751 => "0000000101000000000101110000001000",
			3752 => "0000001100000000001010111000000100",
			3753 => "11111110101000110011101011011001",
			3754 => "00000010001010000011101011011001",
			3755 => "11111110011010100011101011011001",
			3756 => "11111110010111110011101011011001",
			3757 => "0000001100000000001001110100000100",
			3758 => "00000101111011000011101011011001",
			3759 => "11111110100000110011101011011001",
			3760 => "0000000111000000000111010000001000",
			3761 => "0000001011000000000100010000000100",
			3762 => "00000001110111000011101011011001",
			3763 => "00000110001001010011101011011001",
			3764 => "11111110100110100011101011011001",
			3765 => "11111110010111010011101011011001",
			3766 => "0000000000000000001001101000111000",
			3767 => "0000001101000000000101110000010100",
			3768 => "0000001100000000001010111000000100",
			3769 => "00000000000000000011101110011101",
			3770 => "0000000001000000000111101000001100",
			3771 => "0000001011000000000110110100001000",
			3772 => "0000000111000000000011100000000100",
			3773 => "00000000000000000011101110011101",
			3774 => "00000000111010000011101110011101",
			3775 => "00000000000000000011101110011101",
			3776 => "00000000000000000011101110011101",
			3777 => "0000001100000000001000000000011000",
			3778 => "0000001011000000000110110100001100",
			3779 => "0000000101000000001100100100000100",
			3780 => "00000000000000000011101110011101",
			3781 => "0000001111000000000010000100000100",
			3782 => "00000000000000000011101110011101",
			3783 => "11111111000111100011101110011101",
			3784 => "0000000000000000000001110000001000",
			3785 => "0000000010000000001110110100000100",
			3786 => "00000000000000000011101110011101",
			3787 => "11111111110011010011101110011101",
			3788 => "00000000001001100011101110011101",
			3789 => "0000000010000000001010000100001000",
			3790 => "0000000010000000001110110100000100",
			3791 => "00000000000000000011101110011101",
			3792 => "00000000110011110011101110011101",
			3793 => "00000000000000000011101110011101",
			3794 => "0000001110000000000111011000000100",
			3795 => "11111110110001100011101110011101",
			3796 => "0000001111000000000000010000000100",
			3797 => "00000000101111100011101110011101",
			3798 => "0000000111000000000110100100001100",
			3799 => "0000000010000000001101101100001000",
			3800 => "0000001101000000001110000100000100",
			3801 => "00000000000000000011101110011101",
			3802 => "00000000010000110011101110011101",
			3803 => "00000000000000000011101110011101",
			3804 => "0000000010000000001000100000001000",
			3805 => "0000001100000000000100011000000100",
			3806 => "11111111000001000011101110011101",
			3807 => "00000000000000000011101110011101",
			3808 => "0000000010000000001101101100001000",
			3809 => "0000001000000000000101000100000100",
			3810 => "00000000100001100011101110011101",
			3811 => "00000000000000000011101110011101",
			3812 => "0000000111000000001000011000000100",
			3813 => "11111111011110000011101110011101",
			3814 => "00000000000000000011101110011101",
			3815 => "0000000111000000000110100100010000",
			3816 => "0000000100000000001100000000000100",
			3817 => "00000000000000000011110001110001",
			3818 => "0000000011000000000111010100001000",
			3819 => "0000001011000000000101100100000100",
			3820 => "11111110101011010011110001110001",
			3821 => "00000000000000000011110001110001",
			3822 => "00000000000000000011110001110001",
			3823 => "0000001011000000001011011100100100",
			3824 => "0000001011000000000101100100010000",
			3825 => "0000000001000000001101111100001100",
			3826 => "0000000011000000000110111100000100",
			3827 => "00000000000000000011110001110001",
			3828 => "0000000100000000000011000000000100",
			3829 => "00000000110100100011110001110001",
			3830 => "00000000000000000011110001110001",
			3831 => "00000000000000000011110001110001",
			3832 => "0000000111000000000110100100000100",
			3833 => "00000000000000000011110001110001",
			3834 => "0000001111000000001001100000000100",
			3835 => "00000000000000000011110001110001",
			3836 => "0000001100000000001010111000000100",
			3837 => "00000000000000000011110001110001",
			3838 => "0000000111000000001000011000000100",
			3839 => "11111111000110010011110001110001",
			3840 => "00000000000000000011110001110001",
			3841 => "0000000100000000000001011100100000",
			3842 => "0000000111000000000110100100001100",
			3843 => "0000001001000000001001111100001000",
			3844 => "0000000011000000001100000000000100",
			3845 => "00000000000000000011110001110001",
			3846 => "11111111101101000011110001110001",
			3847 => "00000000000000000011110001110001",
			3848 => "0000000001000000000000111100010000",
			3849 => "0000001010000000001010100000001000",
			3850 => "0000000011000000000111010100000100",
			3851 => "00000000011110010011110001110001",
			3852 => "00000000000000000011110001110001",
			3853 => "0000000111000000001111011100000100",
			3854 => "11111111100011100011110001110001",
			3855 => "00000000000000000011110001110001",
			3856 => "00000001001011100011110001110001",
			3857 => "0000001110000000001100111000001100",
			3858 => "0000000101000000000011001000001000",
			3859 => "0000000011000000000011000000000100",
			3860 => "11111111011100000011110001110001",
			3861 => "00000000000000000011110001110001",
			3862 => "00000000000000000011110001110001",
			3863 => "0000000100000000001000110100001000",
			3864 => "0000001101000000001100010100000100",
			3865 => "00000000100110000011110001110001",
			3866 => "00000000000000000011110001110001",
			3867 => "00000000000000000011110001110001",
			3868 => "0000000001000000001110010101000000",
			3869 => "0000000100000000001000100000111000",
			3870 => "0000001101000000000010011100010000",
			3871 => "0000000001000000001001011000000100",
			3872 => "00000000000000000011110101001101",
			3873 => "0000001101000000000101001000000100",
			3874 => "00000000000000000011110101001101",
			3875 => "0000001010000000000111101100000100",
			3876 => "00000000000000000011110101001101",
			3877 => "00000000100110100011110101001101",
			3878 => "0000000010000000000010000100010000",
			3879 => "0000001101000000000101110000000100",
			3880 => "00000000000000000011110101001101",
			3881 => "0000001010000000001010100000001000",
			3882 => "0000000010000000000110010000000100",
			3883 => "00000000000000000011110101001101",
			3884 => "11111111010110100011110101001101",
			3885 => "00000000000000000011110101001101",
			3886 => "0000000111000000000001101000001100",
			3887 => "0000001110000000001100000000001000",
			3888 => "0000001011000000000110110100000100",
			3889 => "11111111110001100011110101001101",
			3890 => "00000000000000000011110101001101",
			3891 => "00000000000000000011110101001101",
			3892 => "0000000001000000001001011000000100",
			3893 => "00000000000000000011110101001101",
			3894 => "0000000010000000001010000100000100",
			3895 => "00000000011100010011110101001101",
			3896 => "00000000000000000011110101001101",
			3897 => "0000001100000000000001101000000100",
			3898 => "11111111010001100011110101001101",
			3899 => "00000000000000000011110101001101",
			3900 => "0000001010000000001000100100010100",
			3901 => "0000000101000000001101000100000100",
			3902 => "00000000000000000011110101001101",
			3903 => "0000001100000000001010111000000100",
			3904 => "00000000000000000011110101001101",
			3905 => "0000000100000000001011110000001000",
			3906 => "0000000001000000001100011000000100",
			3907 => "00000001000000110011110101001101",
			3908 => "00000000000000000011110101001101",
			3909 => "00000000000000000011110101001101",
			3910 => "0000001110000000001100111000001000",
			3911 => "0000000111000000000110100100000100",
			3912 => "00000000000000000011110101001101",
			3913 => "11111111101111000011110101001101",
			3914 => "0000000100000000001000110100010000",
			3915 => "0000001100000000000100011000000100",
			3916 => "00000000000000000011110101001101",
			3917 => "0000000011000000001101101100000100",
			3918 => "00000000000000000011110101001101",
			3919 => "0000000111000000000111010000000100",
			3920 => "00000000011101010011110101001101",
			3921 => "00000000000000000011110101001101",
			3922 => "00000000000000000011110101001101",
			3923 => "0000001100000000001010111000010100",
			3924 => "0000000000000000000110001000010000",
			3925 => "0000000010000000000111011000001000",
			3926 => "0000001100000000001010111000000100",
			3927 => "11111111011111110011111000110001",
			3928 => "00000000000000000011111000110001",
			3929 => "0000001011000000000000011100000100",
			3930 => "00000000000000000011111000110001",
			3931 => "00000000110010010011111000110001",
			3932 => "11111110100011110011111000110001",
			3933 => "0000001100000000001011000001000000",
			3934 => "0000001101000000000100101000100100",
			3935 => "0000000001000000001101111100011100",
			3936 => "0000001101000000001111010000010000",
			3937 => "0000000101000000000010110100001000",
			3938 => "0000000000000000001011010100000100",
			3939 => "00000000111100100011111000110001",
			3940 => "00000000000000000011111000110001",
			3941 => "0000000101000000000110100000000100",
			3942 => "11111110111001110011111000110001",
			3943 => "00000000000000000011111000110001",
			3944 => "0000000110000000001101111100000100",
			3945 => "00000000000000000011111000110001",
			3946 => "0000001011000000000110110100000100",
			3947 => "00000001010001000011111000110001",
			3948 => "00000000000000000011111000110001",
			3949 => "0000001011000000001011011100000100",
			3950 => "11111111001101100011111000110001",
			3951 => "00000000000000000011111000110001",
			3952 => "0000001100000000001011000000001100",
			3953 => "0000000001000000001110010100001000",
			3954 => "0000001110000000000010000100000100",
			3955 => "00000000000000000011111000110001",
			3956 => "11111110110010110011111000110001",
			3957 => "00000000000000000011111000110001",
			3958 => "0000001100000000001011000000001100",
			3959 => "0000000101000000001111010000001000",
			3960 => "0000000101000000000001000000000100",
			3961 => "00000000000000000011111000110001",
			3962 => "00000000101101000011111000110001",
			3963 => "00000000000000000011111000110001",
			3964 => "11111111100011110011111000110001",
			3965 => "0000000010000000001110110100001100",
			3966 => "0000000001000000000000111100001000",
			3967 => "0000000100000000000010000100000100",
			3968 => "00000000000000000011111000110001",
			3969 => "11111111110000110011111000110001",
			3970 => "00000000000000000011111000110001",
			3971 => "0000000001000000001100011000010000",
			3972 => "0000000001000000001001011000000100",
			3973 => "00000000000000000011111000110001",
			3974 => "0000000100000000001000110100001000",
			3975 => "0000000101000000001101000100000100",
			3976 => "00000000000000000011111000110001",
			3977 => "00000001000010000011111000110001",
			3978 => "00000000000000000011111000110001",
			3979 => "00000000000000000011111000110001",
			3980 => "0000000101000000001101000100011100",
			3981 => "0000000000000000000001010100001100",
			3982 => "0000001100000000000100011000000100",
			3983 => "00000000000000000011111100110101",
			3984 => "0000001011000000000000011100000100",
			3985 => "00000000110001100011111100110101",
			3986 => "00000000000000000011111100110101",
			3987 => "0000001110000000000111010100001000",
			3988 => "0000000100000000000010000100000100",
			3989 => "00000000000000000011111100110101",
			3990 => "11111110011011100011111100110101",
			3991 => "0000000110000000000100111100000100",
			3992 => "00000000100000010011111100110101",
			3993 => "00000000000000000011111100110101",
			3994 => "0000000010000000000111011000110000",
			3995 => "0000000000000000000001010100100100",
			3996 => "0000000001000000001001011000010000",
			3997 => "0000000111000000000001101000000100",
			3998 => "00000000000000000011111100110101",
			3999 => "0000000011000000000110111100001000",
			4000 => "0000001110000000000110010000000100",
			4001 => "00000000000000000011111100110101",
			4002 => "00000001100001100011111100110101",
			4003 => "00000000000000000011111100110101",
			4004 => "0000000010000000000010000100010000",
			4005 => "0000000010000000000110010000001000",
			4006 => "0000001001000000001111000000000100",
			4007 => "00000000000000000011111100110101",
			4008 => "00000000001000100011111100110101",
			4009 => "0000000111000000000001101000000100",
			4010 => "00000000000000000011111100110101",
			4011 => "11111110111010100011111100110101",
			4012 => "00000000000000000011111100110101",
			4013 => "0000000001000000001001011000000100",
			4014 => "00000000000000000011111100110101",
			4015 => "0000000011000000000111010100000100",
			4016 => "00000001010011010011111100110101",
			4017 => "00000000000000000011111100110101",
			4018 => "0000001001000000000100101100011100",
			4019 => "0000001011000000000100010000001100",
			4020 => "0000000101000000001100100100000100",
			4021 => "00000000010100010011111100110101",
			4022 => "0000001100000000001001110100000100",
			4023 => "11111110101100010011111100110101",
			4024 => "00000000000000000011111100110101",
			4025 => "0000001010000000001010100100000100",
			4026 => "00000000110111000011111100110101",
			4027 => "0000001010000000001010100100000100",
			4028 => "11111111101101100011111100110101",
			4029 => "0000000010000000000110101100000100",
			4030 => "00000000010000000011111100110101",
			4031 => "00000000000000000011111100110101",
			4032 => "0000000100000000000001011100001000",
			4033 => "0000000101000000001101000100000100",
			4034 => "00000000000000000011111100110101",
			4035 => "00000001010000110011111100110101",
			4036 => "0000000011000000001000100000000100",
			4037 => "11111110110101000011111100110101",
			4038 => "0000001100000000001001001000001000",
			4039 => "0000000001000000000100110100000100",
			4040 => "00000001001000110011111100110101",
			4041 => "00000000000000000011111100110101",
			4042 => "0000000111000000000101110100000100",
			4043 => "11111111010110010011111100110101",
			4044 => "00000000000000000011111100110101",
			4045 => "0000000000000000001010101101010000",
			4046 => "0000001110000000001100111001000100",
			4047 => "0000000000000000001011010100100100",
			4048 => "0000001010000000000010101100011000",
			4049 => "0000000000000000001001101000010000",
			4050 => "0000001000000000001000100100001000",
			4051 => "0000000100000000001100010000000100",
			4052 => "00000000100111100011111111011001",
			4053 => "11111111010110110011111111011001",
			4054 => "0000001101000000001010001000000100",
			4055 => "00000000111100100011111111011001",
			4056 => "11111111110011110011111111011001",
			4057 => "0000000111000000001001001000000100",
			4058 => "00000000000000000011111111011001",
			4059 => "11111110011111010011111111011001",
			4060 => "0000000110000000001101011000000100",
			4061 => "00000000000000000011111111011001",
			4062 => "0000001011000000000000011100000100",
			4063 => "00000000000000000011111111011001",
			4064 => "00000001011111010011111111011001",
			4065 => "0000001110000000001000001100010000",
			4066 => "0000000100000000001011101100001000",
			4067 => "0000001101000000000101001000000100",
			4068 => "00000000000000000011111111011001",
			4069 => "00000001000001110011111111011001",
			4070 => "0000000111000000000001101000000100",
			4071 => "11111110001101000011111111011001",
			4072 => "00000000000000000011111111011001",
			4073 => "0000000000000000000111000100001100",
			4074 => "0000000000000000000110001000001000",
			4075 => "0000001011000000000110110100000100",
			4076 => "00000000000000000011111111011001",
			4077 => "11111110110100000011111111011001",
			4078 => "00000001010100100011111111011001",
			4079 => "11111110100110000011111111011001",
			4080 => "0000001101000000001100010100000100",
			4081 => "00000001010101110011111111011001",
			4082 => "0000001000000000000001010100000100",
			4083 => "11111111111010110011111111011001",
			4084 => "00000000000000000011111111011001",
			4085 => "11111110011111000011111111011001",
			4086 => "0000001011000000001011011101000100",
			4087 => "0000001110000000000111011000100100",
			4088 => "0000000000000000001100000100011100",
			4089 => "0000001000000000001000100100010100",
			4090 => "0000000100000000001100010000001100",
			4091 => "0000000011000000000111100000000100",
			4092 => "00000000000000000100000011111101",
			4093 => "0000000011000000001100010000000100",
			4094 => "00000000001110110100000011111101",
			4095 => "00000000000000000100000011111101",
			4096 => "0000001011000000000101100100000100",
			4097 => "11111110111100110100000011111101",
			4098 => "00000000000000000100000011111101",
			4099 => "0000000001000000000000111100000100",
			4100 => "00000000000000000100000011111101",
			4101 => "00000000110000100100000011111101",
			4102 => "0000000100000000001010000100000100",
			4103 => "00000000000000000100000011111101",
			4104 => "11111110011101010100000011111101",
			4105 => "0000001011000000000101100100001000",
			4106 => "0000000000000000001111001000000100",
			4107 => "00000001000101010100000011111101",
			4108 => "00000000000000000100000011111101",
			4109 => "0000000100000000001111100100000100",
			4110 => "00000000000000000100000011111101",
			4111 => "0000001001000000000111101100000100",
			4112 => "11111110111100000100000011111101",
			4113 => "0000001001000000001010100000001000",
			4114 => "0000001000000000000110011100000100",
			4115 => "00000000011100000100000011111101",
			4116 => "00000000000000000100000011111101",
			4117 => "0000001101000000000101110000000100",
			4118 => "11111111001111000100000011111101",
			4119 => "00000000000000000100000011111101",
			4120 => "0000000101000000000111100000011000",
			4121 => "0000000001000000001101111100010000",
			4122 => "0000001011000000000010001000001100",
			4123 => "0000000110000000001101111100000100",
			4124 => "00000000000000000100000011111101",
			4125 => "0000000000000000000010101000000100",
			4126 => "00000001010010000100000011111101",
			4127 => "00000000000000000100000011111101",
			4128 => "00000000000000000100000011111101",
			4129 => "0000000101000000001100100100000100",
			4130 => "11111111101111010100000011111101",
			4131 => "00000000000000000100000011111101",
			4132 => "0000001100000000001011000000010000",
			4133 => "0000001110000000001100010000000100",
			4134 => "00000000000000000100000011111101",
			4135 => "0000000011000000001101101100001000",
			4136 => "0000001100000000000100011000000100",
			4137 => "11111110101100110100000011111101",
			4138 => "00000000000000000100000011111101",
			4139 => "00000000000000000100000011111101",
			4140 => "0000000000000000000001010100010000",
			4141 => "0000000011000000000110111100001000",
			4142 => "0000001111000000000010000100000100",
			4143 => "00000000000000000100000011111101",
			4144 => "00000000101000000100000011111101",
			4145 => "0000000101000000001111010000000100",
			4146 => "11111111000011100100000011111101",
			4147 => "00000000000000000100000011111101",
			4148 => "0000001101000000001100010100010000",
			4149 => "0000001100000000000110100100001000",
			4150 => "0000000000000000000111000000000100",
			4151 => "00000000111011100100000011111101",
			4152 => "00000000000000000100000011111101",
			4153 => "0000000110000000001010011000000100",
			4154 => "00000000000000000100000011111101",
			4155 => "11111111110001000100000011111101",
			4156 => "0000001001000000000100101100000100",
			4157 => "00000000000000000100000011111101",
			4158 => "11111111001100000100000011111101",
			4159 => "0000001100000000001010111000011000",
			4160 => "0000000000000000000110001000010100",
			4161 => "0000000111000000001001001000001000",
			4162 => "0000000010000000001111010100000100",
			4163 => "11111111010101000100001000000001",
			4164 => "00000000000000000100001000000001",
			4165 => "0000001010000000000111101100000100",
			4166 => "00000000000000000100001000000001",
			4167 => "0000000111000000000110100100000100",
			4168 => "00000000000000000100001000000001",
			4169 => "00000000011000000100001000000001",
			4170 => "11111110100001000100001000000001",
			4171 => "0000000101000000001100100100101100",
			4172 => "0000000001000000001101111100100000",
			4173 => "0000001101000000001110000100001100",
			4174 => "0000000000000000000001010100000100",
			4175 => "00000000000000000100001000000001",
			4176 => "0000000111000000000001101000000100",
			4177 => "11111111000011010100001000000001",
			4178 => "00000000000000000100001000000001",
			4179 => "0000000000000000001111001000001000",
			4180 => "0000000110000000001101111100000100",
			4181 => "00000000000000000100001000000001",
			4182 => "00000001001101100100001000000001",
			4183 => "0000001001000000001010100000000100",
			4184 => "11111111111101100100001000000001",
			4185 => "0000000011000000001101101100000100",
			4186 => "00000000000101110100001000000001",
			4187 => "00000000000000000100001000000001",
			4188 => "0000001100000000000100011000000100",
			4189 => "00000000000000000100001000000001",
			4190 => "0000001100000000001000000000000100",
			4191 => "11111111001000000100001000000001",
			4192 => "00000000000000000100001000000001",
			4193 => "0000000101000000000111100000010000",
			4194 => "0000001101000000000111111100001100",
			4195 => "0000000011000000001111100100001000",
			4196 => "0000001111000000000110111100000100",
			4197 => "00000000000000000100001000000001",
			4198 => "11111110111011100100001000000001",
			4199 => "00000000000000000100001000000001",
			4200 => "00000000100010100100001000000001",
			4201 => "0000000001000000000000111100011000",
			4202 => "0000000011000000000110111100001000",
			4203 => "0000001000000000001000100100000100",
			4204 => "00000000000000000100001000000001",
			4205 => "00000000111101110100001000000001",
			4206 => "0000000111000000001000011000001000",
			4207 => "0000000111000000000001101000000100",
			4208 => "00000000000000000100001000000001",
			4209 => "00000000110000000100001000000001",
			4210 => "0000000000000000000001010100000100",
			4211 => "11111110111101010100001000000001",
			4212 => "00000000000000000100001000000001",
			4213 => "0000001101000000001100010100001100",
			4214 => "0000000001000000001010011000001000",
			4215 => "0000000100000000000101000000000100",
			4216 => "00000001010010000100001000000001",
			4217 => "00000000000000000100001000000001",
			4218 => "00000000000000000100001000000001",
			4219 => "0000000111000000000000011100000100",
			4220 => "11111111001001110100001000000001",
			4221 => "0000000010000000001101101100000100",
			4222 => "00000000110111010100001000000001",
			4223 => "11111111111010110100001000000001",
			4224 => "0000000000000000001010101101010100",
			4225 => "0000001110000000001100111001001000",
			4226 => "0000000000000000001011010100100100",
			4227 => "0000001000000000001000100100010000",
			4228 => "0000000110000000000100110100001100",
			4229 => "0000000111000000001111011100001000",
			4230 => "0000000110000000001101111100000100",
			4231 => "11111111110010110100001010101101",
			4232 => "00000000110000010100001010101101",
			4233 => "11111110101110010100001010101101",
			4234 => "11111110100100010100001010101101",
			4235 => "0000000010000000001100000000001000",
			4236 => "0000001101000000000001000000000100",
			4237 => "00000000000000000100001010101101",
			4238 => "00000001011000000100001010101101",
			4239 => "0000000110000000001011001100001000",
			4240 => "0000000000000000001001101000000100",
			4241 => "00000000001100000100001010101101",
			4242 => "11111111000100100100001010101101",
			4243 => "00000001011001010100001010101101",
			4244 => "0000001110000000001000001100010100",
			4245 => "0000000101000000000010110100001000",
			4246 => "0000001011000000000000011100000100",
			4247 => "11111111101011010100001010101101",
			4248 => "00000000100111110100001010101101",
			4249 => "0000000101000000000001000000001000",
			4250 => "0000000111000000001001001000000100",
			4251 => "00000000000000000100001010101101",
			4252 => "11111110010110010100001010101101",
			4253 => "00000000000000000100001010101101",
			4254 => "0000000000000000000111000100001100",
			4255 => "0000000000000000000110001000001000",
			4256 => "0000001011000000000110110100000100",
			4257 => "00000000000000000100001010101101",
			4258 => "11111110101110010100001010101101",
			4259 => "00000001010111000100001010101101",
			4260 => "11111110100011000100001010101101",
			4261 => "0000001101000000001010001000000100",
			4262 => "00000001011110010100001010101101",
			4263 => "0000001000000000000001010100000100",
			4264 => "11111111110010100100001010101101",
			4265 => "00000000000000000100001010101101",
			4266 => "11111110011110010100001010101101",
			4267 => "0000001100000000001010111000010000",
			4268 => "0000000000000000000110001000001100",
			4269 => "0000001110000000001100000000001000",
			4270 => "0000000111000000000110100100000100",
			4271 => "11111111001011110100001110110001",
			4272 => "00000000000000000100001110110001",
			4273 => "00000000011010100100001110110001",
			4274 => "11111110011110010100001110110001",
			4275 => "0000000101000000001100100100110000",
			4276 => "0000000001000000001101111100100100",
			4277 => "0000000101000000001101000100011000",
			4278 => "0000000011000000001010000100010000",
			4279 => "0000000000000000000001010100001000",
			4280 => "0000001100000000000100011000000100",
			4281 => "00000000000000000100001110110001",
			4282 => "00000000011111000100001110110001",
			4283 => "0000001100000000001010111000000100",
			4284 => "00000000000000000100001110110001",
			4285 => "11111111010011110100001110110001",
			4286 => "0000000001000000000001111000000100",
			4287 => "00000001000001000100001110110001",
			4288 => "00000000000000000100001110110001",
			4289 => "0000000110000000001101111100000100",
			4290 => "00000000000000000100001110110001",
			4291 => "0000000000000000000001110100000100",
			4292 => "00000001010100110100001110110001",
			4293 => "00000000000000000100001110110001",
			4294 => "0000001100000000000100011000000100",
			4295 => "00000000000000000100001110110001",
			4296 => "0000001100000000001000000000000100",
			4297 => "11111111000100000100001110110001",
			4298 => "00000000000000000100001110110001",
			4299 => "0000000101000000000111100000011100",
			4300 => "0000001111000000000110111100010000",
			4301 => "0000000110000000000100110100001000",
			4302 => "0000000011000000001100010000000100",
			4303 => "00000000000000000100001110110001",
			4304 => "11111111111101000100001110110001",
			4305 => "0000001110000000000110010000000100",
			4306 => "00000000000000000100001110110001",
			4307 => "00000000111111100100001110110001",
			4308 => "0000000011000000001111100100001000",
			4309 => "0000001011000000001011011100000100",
			4310 => "11111110101110110100001110110001",
			4311 => "00000000000000000100001110110001",
			4312 => "00000000000000000100001110110001",
			4313 => "0000000001000000000000111100011000",
			4314 => "0000000011000000000110111100001000",
			4315 => "0000001000000000001000100100000100",
			4316 => "00000000000000000100001110110001",
			4317 => "00000001001010100100001110110001",
			4318 => "0000000111000000001000011000001000",
			4319 => "0000000111000000000001101000000100",
			4320 => "00000000000000000100001110110001",
			4321 => "00000000110110000100001110110001",
			4322 => "0000001100000000001001110100000100",
			4323 => "11111111000100100100001110110001",
			4324 => "00000000000000000100001110110001",
			4325 => "0000000001000000001010011000001100",
			4326 => "0000000100000000000101000000001000",
			4327 => "0000000101000000001110010000000100",
			4328 => "00000000111110100100001110110001",
			4329 => "00000000000000000100001110110001",
			4330 => "00000000000000000100001110110001",
			4331 => "11111111110011010100001110110001",
			4332 => "0000001100000000000111001000001000",
			4333 => "0000000111000000000110100100000100",
			4334 => "11111110011111110100010010001101",
			4335 => "00000000000000000100010010001101",
			4336 => "0000000000000000001001101000111000",
			4337 => "0000001000000000001000100100011000",
			4338 => "0000000100000000001100010000001100",
			4339 => "0000000011000000001100010000001000",
			4340 => "0000001001000000001111000000000100",
			4341 => "00000000000000000100010010001101",
			4342 => "00000001001110000100010010001101",
			4343 => "00000000000000000100010010001101",
			4344 => "0000000010000000001110110100000100",
			4345 => "11111110100100100100010010001101",
			4346 => "0000001100000000001000000000000100",
			4347 => "11111111011001000100010010001101",
			4348 => "00000000110000110100010010001101",
			4349 => "0000001101000000001010001000010000",
			4350 => "0000001101000000000101001000001000",
			4351 => "0000000001000000001110010100000100",
			4352 => "00000000000000000100010010001101",
			4353 => "11111111001111000100010010001101",
			4354 => "0000000011000000000000010000000100",
			4355 => "00000001010111100100010010001101",
			4356 => "00000000000000000100010010001101",
			4357 => "0000000111000000001111011100001000",
			4358 => "0000000001000000000000111100000100",
			4359 => "11111110110001100100010010001101",
			4360 => "00000000010000100100010010001101",
			4361 => "0000000110000000001100011000000100",
			4362 => "00000001000111000100010010001101",
			4363 => "00000000000000000100010010001101",
			4364 => "0000001010000000000010101100000100",
			4365 => "11111110100000010100010010001101",
			4366 => "0000000000000000001011010100001100",
			4367 => "0000000110000000001101011000000100",
			4368 => "00000000000000000100010010001101",
			4369 => "0000000010000000000111011000000100",
			4370 => "00000000000000000100010010001101",
			4371 => "00000001011001010100010010001101",
			4372 => "0000001110000000001000001100010000",
			4373 => "0000000100000000001011101100001000",
			4374 => "0000001101000000000101001000000100",
			4375 => "00000000000000000100010010001101",
			4376 => "00000000111111000100010010001101",
			4377 => "0000000111000000000001101000000100",
			4378 => "11111110010000100100010010001101",
			4379 => "00000000000000000100010010001101",
			4380 => "0000000000000000000010101000001000",
			4381 => "0000000011000000001100111000000100",
			4382 => "00000000000000000100010010001101",
			4383 => "00000001010010100100010010001101",
			4384 => "0000000011000000001000101000000100",
			4385 => "11111110110010010100010010001101",
			4386 => "00000000000000000100010010001101",
			4387 => "0000001001000000001001100100010100",
			4388 => "0000000110000000000000111100010000",
			4389 => "0000000110000000000000111100000100",
			4390 => "00000000000000000100010110100001",
			4391 => "0000000000000000000011101000000100",
			4392 => "00000000000000000100010110100001",
			4393 => "0000000000000000000000110000000100",
			4394 => "00000000001011010100010110100001",
			4395 => "00000000000000000100010110100001",
			4396 => "11111110011011010100010110100001",
			4397 => "0000001100000000000100011001000000",
			4398 => "0000000000000000000110001000100000",
			4399 => "0000000111000000000110100100010000",
			4400 => "0000000111000000001001001000001000",
			4401 => "0000001101000000000001000000000100",
			4402 => "00000000000000000100010110100001",
			4403 => "00000000100101010100010110100001",
			4404 => "0000001011000000000000011100000100",
			4405 => "00000000000000000100010110100001",
			4406 => "11111110000010000100010110100001",
			4407 => "0000001101000000000100101000001100",
			4408 => "0000001001000000001111000000000100",
			4409 => "00000000000000000100010110100001",
			4410 => "0000001100000000000100011000000100",
			4411 => "00000001100010010100010110100001",
			4412 => "00000000000010000100010110100001",
			4413 => "11111111000001000100010110100001",
			4414 => "0000001011000000001011011100010000",
			4415 => "0000000111000000001000011000001100",
			4416 => "0000001001000000001010100000000100",
			4417 => "11111101110010010100010110100001",
			4418 => "0000001001000000001010100000000100",
			4419 => "00000000000000000100010110100001",
			4420 => "11111111010001010100010110100001",
			4421 => "00000000000000000100010110100001",
			4422 => "0000001100000000000100011000000100",
			4423 => "00000000000000000100010110100001",
			4424 => "0000001100000000000100011000001000",
			4425 => "0000000010000000001110000000000100",
			4426 => "00000000010100110100010110100001",
			4427 => "00000000000000000100010110100001",
			4428 => "00000000000000000100010110100001",
			4429 => "0000001101000000001100010100101000",
			4430 => "0000000011000000001011101100011100",
			4431 => "0000000000000000001111001000010000",
			4432 => "0000000110000000001011001100001000",
			4433 => "0000000010000000001000001100000100",
			4434 => "00000000001110000100010110100001",
			4435 => "11111110011110010100010110100001",
			4436 => "0000000011000000001111010100000100",
			4437 => "00000000000000000100010110100001",
			4438 => "00000001011001100100010110100001",
			4439 => "0000001100000000001000000000001000",
			4440 => "0000001100000000000100011000000100",
			4441 => "00000000000000000100010110100001",
			4442 => "11111110011011010100010110100001",
			4443 => "00000000000000000100010110100001",
			4444 => "0000000001000000001010011000001000",
			4445 => "0000000000000000000111000000000100",
			4446 => "00000001101110010100010110100001",
			4447 => "11111111111101010100010110100001",
			4448 => "11111111101111010100010110100001",
			4449 => "0000001001000000000100101100001100",
			4450 => "0000000001000000001011111100000100",
			4451 => "11111111010111100100010110100001",
			4452 => "0000001101000000001110110100000100",
			4453 => "00000000101111110100010110100001",
			4454 => "00000000000000000100010110100001",
			4455 => "11111110100101000100010110100001",
			4456 => "0000001101000000001110000100010100",
			4457 => "0000000000000000000101000100001100",
			4458 => "0000000111000000001011000000000100",
			4459 => "00000000000000000100011010110101",
			4460 => "0000000101000000001101000100000100",
			4461 => "00000000001001110100011010110101",
			4462 => "00000000000000000100011010110101",
			4463 => "0000000111000000000110100100000100",
			4464 => "11111110011101100100011010110101",
			4465 => "00000000000000000100011010110101",
			4466 => "0000001001000000000111101101010000",
			4467 => "0000000100000000000000010000110000",
			4468 => "0000001101000000000010011100010100",
			4469 => "0000001101000000000101001000001100",
			4470 => "0000001100000000000100011000001000",
			4471 => "0000000111000000000110100100000100",
			4472 => "11111111010110010100011010110101",
			4473 => "00000000000000000100011010110101",
			4474 => "00000000000000000100011010110101",
			4475 => "0000001010000000000000001000000100",
			4476 => "00000000000000000100011010110101",
			4477 => "00000001011010110100011010110101",
			4478 => "0000000000000000000001010100001100",
			4479 => "0000000101000000001111010000001000",
			4480 => "0000000010000000000110010000000100",
			4481 => "00000000000000000100011010110101",
			4482 => "11111110100110110100011010110101",
			4483 => "11111111110101100100011010110101",
			4484 => "0000000000000000001100000100001000",
			4485 => "0000001100000000000100011000000100",
			4486 => "00000000000000000100011010110101",
			4487 => "00000001000001010100011010110101",
			4488 => "0000000001000000001011111100000100",
			4489 => "11111110101111010100011010110101",
			4490 => "00000000000110100100011010110101",
			4491 => "0000001100000000001000011000010100",
			4492 => "0000000100000000001101101100010000",
			4493 => "0000001010000000000010101100001000",
			4494 => "0000000111000000001111011100000100",
			4495 => "11111110011101000100011010110101",
			4496 => "00000000000000000100011010110101",
			4497 => "0000000101000000001110101000000100",
			4498 => "11111111101100010100011010110101",
			4499 => "00000001000101010100011010110101",
			4500 => "11111110011111000100011010110101",
			4501 => "0000000001000000000001000100000100",
			4502 => "00000000000000000100011010110101",
			4503 => "0000000110000000001000010000000100",
			4504 => "00000000111000010100011010110101",
			4505 => "00000000000000000100011010110101",
			4506 => "0000000000000000000001110100001100",
			4507 => "0000001010000000000011101000000100",
			4508 => "11111111111100110100011010110101",
			4509 => "0000000101000000000111111100000100",
			4510 => "00000001010101110100011010110101",
			4511 => "00000000000000000100011010110101",
			4512 => "0000001110000000001100111000000100",
			4513 => "11111110101100010100011010110101",
			4514 => "0000000110000000001000010000001000",
			4515 => "0000001010000000001000100100000100",
			4516 => "00000000000000000100011010110101",
			4517 => "11111111011111100100011010110101",
			4518 => "0000001111000000001011110000001000",
			4519 => "0000000001000000001010011000000100",
			4520 => "00000001000101010100011010110101",
			4521 => "00000000000000000100011010110101",
			4522 => "0000001111000000001110000000000100",
			4523 => "00000000000000000100011010110101",
			4524 => "11111111110000110100011010110101",
			4525 => "0000000000000000001010101101111000",
			4526 => "0000000001000000000000111100111000",
			4527 => "0000000111000000001000011000100000",
			4528 => "0000000111000000000001101000010100",
			4529 => "0000000100000000001100010000001100",
			4530 => "0000000110000000001101111100001000",
			4531 => "0000000110000000000000111100000100",
			4532 => "00000000100100100100011110101001",
			4533 => "11111111001010000100011110101001",
			4534 => "00000010001111000100011110101001",
			4535 => "0000001001000000000100111100000100",
			4536 => "11111110011011100100011110101001",
			4537 => "00000000001101010100011110101001",
			4538 => "0000000000000000000101000100001000",
			4539 => "0000000011000000001100000000000100",
			4540 => "00000000000000000100011110101001",
			4541 => "11111111110100110100011110101001",
			4542 => "00000010001110000100011110101001",
			4543 => "0000000011000000000110111100001000",
			4544 => "0000001000000000001000100100000100",
			4545 => "00000000000000000100011110101001",
			4546 => "00000010101000100100011110101001",
			4547 => "0000000000000000000001010100000100",
			4548 => "11111101111010110100011110101001",
			4549 => "0000000111000000001000011000000100",
			4550 => "11111110000010100100011110101001",
			4551 => "0000001000000000001000010100000100",
			4552 => "00000001010001010100011110101001",
			4553 => "11111111000010000100011110101001",
			4554 => "0000000111000000000001101000100100",
			4555 => "0000000100000000000001011100010100",
			4556 => "0000000111000000000001101000010000",
			4557 => "0000000101000000000110100000001000",
			4558 => "0000000001000000000111101000000100",
			4559 => "00000000000011100100011110101001",
			4560 => "11111110010110000100011110101001",
			4561 => "0000001101000000000101110000000100",
			4562 => "00000001010010000100011110101001",
			4563 => "00000000001010010100011110101001",
			4564 => "11111110101011100100011110101001",
			4565 => "0000000011000000001111100100000100",
			4566 => "11111101111100010100011110101001",
			4567 => "0000000010000000001101101100000100",
			4568 => "00000001011000010100011110101001",
			4569 => "0000001000000000000101000100000100",
			4570 => "11111110011001100100011110101001",
			4571 => "00000000000010010100011110101001",
			4572 => "0000000101000000000111111100010000",
			4573 => "0000000001000000000000111100000100",
			4574 => "00000000000000000100011110101001",
			4575 => "0000000101000000001101000100000100",
			4576 => "00000000000000000100011110101001",
			4577 => "0000001111000000000110111000000100",
			4578 => "00000001010111000100011110101001",
			4579 => "00000010011110100100011110101001",
			4580 => "0000000111000000000101110100001000",
			4581 => "0000000101000000001110010000000100",
			4582 => "00000000000000000100011110101001",
			4583 => "11111110101011100100011110101001",
			4584 => "00000000010000010100011110101001",
			4585 => "11111110011010100100011110101001",
			4586 => "0000000111000000000110100100010100",
			4587 => "0000000100000000000111010100001100",
			4588 => "0000000001000000001011111100001000",
			4589 => "0000000001000000001101101000000100",
			4590 => "00000000000000000100100011010101",
			4591 => "00000000010000100100100011010101",
			4592 => "00000000000000000100100011010101",
			4593 => "0000000011000000001010000100000100",
			4594 => "11111110011100010100100011010101",
			4595 => "00000000000000000100100011010101",
			4596 => "0000000111000000000001101000101100",
			4597 => "0000000110000000001011001100100000",
			4598 => "0000000100000000001011101100011100",
			4599 => "0000001010000000001010100000010000",
			4600 => "0000000110000000001101111100001000",
			4601 => "0000001100000000001011000000000100",
			4602 => "00000000000000000100100011010101",
			4603 => "00000000000111010100100011010101",
			4604 => "0000001111000000001001100000000100",
			4605 => "00000000000000000100100011010101",
			4606 => "11111111100100110100100011010101",
			4607 => "0000001001000000000100111100000100",
			4608 => "00000000000000000100100011010101",
			4609 => "0000000011000000000110111100000100",
			4610 => "00000000000000000100100011010101",
			4611 => "00000000111011010100100011010101",
			4612 => "11111111010111110100100011010101",
			4613 => "0000000000000000000001110100001000",
			4614 => "0000000011000000001000001100000100",
			4615 => "00000000000000000100100011010101",
			4616 => "00000001010010110100100011010101",
			4617 => "11111111111101010100100011010101",
			4618 => "0000000110000000001100011000100100",
			4619 => "0000000011000000001010000100011000",
			4620 => "0000000010000000001110110100010000",
			4621 => "0000000100000000001100000000001000",
			4622 => "0000000010000000000010000000000100",
			4623 => "00000000000000000100100011010101",
			4624 => "00000000010110010100100011010101",
			4625 => "0000001100000000001011000000000100",
			4626 => "00000000000000000100100011010101",
			4627 => "11111111101100100100100011010101",
			4628 => "0000000101000000000001000000000100",
			4629 => "00000000000000000100100011010101",
			4630 => "00000001000001100100100011010101",
			4631 => "0000000000000000000001010100000100",
			4632 => "11111111010001100100100011010101",
			4633 => "0000001100000000001011000000000100",
			4634 => "00000000000000000100100011010101",
			4635 => "00000000011100000100100011010101",
			4636 => "0000000101000000000111100000011100",
			4637 => "0000000111000000000001101000001100",
			4638 => "0000001101000000001111010000000100",
			4639 => "00000000000000000100100011010101",
			4640 => "0000001101000000000100101000000100",
			4641 => "11111110111001100100100011010101",
			4642 => "00000000000000000100100011010101",
			4643 => "0000000111000000001000011000001000",
			4644 => "0000000110000000000100111100000100",
			4645 => "00000000010101000100100011010101",
			4646 => "00000000000000000100100011010101",
			4647 => "0000001101000000000101110000000100",
			4648 => "00000000000000000100100011010101",
			4649 => "11111111010000100100100011010101",
			4650 => "0000001101000000001010001000001000",
			4651 => "0000000000000000000010101000000100",
			4652 => "00000000110001000100100011010101",
			4653 => "00000000000000000100100011010101",
			4654 => "0000001100000000001001110100001000",
			4655 => "0000000101000000001001010000000100",
			4656 => "00000000000000000100100011010101",
			4657 => "11111111000111100100100011010101",
			4658 => "0000000001000000000000111100000100",
			4659 => "00000000000000000100100011010101",
			4660 => "00000000010101100100100011010101",
			4661 => "0000000000000000001010101101110000",
			4662 => "0000001001000000000111101101001100",
			4663 => "0000000000000000001100000100101100",
			4664 => "0000000000000000000001010100011000",
			4665 => "0000001101000000000101110000001100",
			4666 => "0000000110000000001101111100000100",
			4667 => "00000000000000000100100110111001",
			4668 => "0000000011000000001100000000000100",
			4669 => "00000001001011010100100110111001",
			4670 => "00000000000000000100100110111001",
			4671 => "0000000101000000001111010000001000",
			4672 => "0000001100000000000100011000000100",
			4673 => "00000000000000000100100110111001",
			4674 => "11111110100101110100100110111001",
			4675 => "11111111111000010100100110111001",
			4676 => "0000000101000000000110100000000100",
			4677 => "11111111010010110100100110111001",
			4678 => "0000000011000000001000001100001000",
			4679 => "0000001001000000001111000000000100",
			4680 => "00000000000000000100100110111001",
			4681 => "00000001011100010100100110111001",
			4682 => "0000001001000000000100111100000100",
			4683 => "11111111100000110100100110111001",
			4684 => "00000000010100110100100110111001",
			4685 => "0000000111000000000111010000011100",
			4686 => "0000001010000000000010101100001100",
			4687 => "0000000111000000001001001000000100",
			4688 => "00000000000000000100100110111001",
			4689 => "0000001101000000001110010000000100",
			4690 => "11111110100010010100100110111001",
			4691 => "00000000000000000100100110111001",
			4692 => "0000000100000000001011101100001000",
			4693 => "0000000111000000001001001000000100",
			4694 => "11111111100000110100100110111001",
			4695 => "00000000111000100100100110111001",
			4696 => "0000000110000000001001100100000100",
			4697 => "11111110100111110100100110111001",
			4698 => "00000000000000000100100110111001",
			4699 => "00000000100010000100100110111001",
			4700 => "0000000000000000000001110100010000",
			4701 => "0000000110000000001011001100000100",
			4702 => "11111111010000010100100110111001",
			4703 => "0000000011000000000111010100000100",
			4704 => "00000000000000000100100110111001",
			4705 => "0000000101000000000111111100000100",
			4706 => "00000001010100110100100110111001",
			4707 => "00000000000000000100100110111001",
			4708 => "0000001110000000001100111000000100",
			4709 => "11111110110000100100100110111001",
			4710 => "0000000110000000001000010000001000",
			4711 => "0000000100000000001011110000000100",
			4712 => "00000000000000000100100110111001",
			4713 => "11111111101000110100100110111001",
			4714 => "0000000111000000000000011100000100",
			4715 => "00000001000111010100100110111001",
			4716 => "00000000000000000100100110111001",
			4717 => "11111110100000110100100110111001",
			4718 => "0000000000000000001010101101100100",
			4719 => "0000000110000000000100111101011000",
			4720 => "0000000000000000001001101000111000",
			4721 => "0000000111000000001000011000011100",
			4722 => "0000000101000000000110100000001100",
			4723 => "0000000001000000001011111100001000",
			4724 => "0000000111000000001011000000000100",
			4725 => "11111111001100110100101010000101",
			4726 => "00000000101100010100101010000101",
			4727 => "11111110010010010100101010000101",
			4728 => "0000001010000000000000001000001000",
			4729 => "0000001101000000001111010000000100",
			4730 => "00000000111010010100101010000101",
			4731 => "11111110111001010100101010000101",
			4732 => "0000001111000000001010000100000100",
			4733 => "00000001011000100100101010000101",
			4734 => "00000000001011100100101010000101",
			4735 => "0000000111000000001000011000010000",
			4736 => "0000001001000000000100111100001000",
			4737 => "0000000011000000000110111100000100",
			4738 => "00000000000000000100101010000101",
			4739 => "11111101111000110100101010000101",
			4740 => "0000000011000000001000001100000100",
			4741 => "00000001010010010100101010000101",
			4742 => "11111101101000110100101010000101",
			4743 => "0000001011000000000100010000001000",
			4744 => "0000001011000000000010001000000100",
			4745 => "00000001010100110100101010000101",
			4746 => "11111111000111000100101010000101",
			4747 => "00000001110110010100101010000101",
			4748 => "0000001110000000000111011000001100",
			4749 => "0000000000000000001001101000001000",
			4750 => "0000000011000000001110110100000100",
			4751 => "00000000000000000100101010000101",
			4752 => "11111100100101000100101010000101",
			4753 => "11111110011111010100101010000101",
			4754 => "0000000100000000001000100000000100",
			4755 => "00000001100110100100101010000101",
			4756 => "0000001110000000000111010100001000",
			4757 => "0000000111000000000110100100000100",
			4758 => "00000000100100010100101010000101",
			4759 => "11111101011100010100101010000101",
			4760 => "0000000000000000000111000100000100",
			4761 => "00000000101101000100101010000101",
			4762 => "11111110100111100100101010000101",
			4763 => "0000001011000000001010010100001000",
			4764 => "0000000101000000001110000100000100",
			4765 => "00000000000000100100101010000101",
			4766 => "00000010011101010100101010000101",
			4767 => "11111111010100100100101010000101",
			4768 => "11111110011010110100101010000101",
			4769 => "0000001100000000000111001000000100",
			4770 => "11111110100110100100101110011011",
			4771 => "0000000101000000000111100000111100",
			4772 => "0000000101000000001100100100101000",
			4773 => "0000000101000000001100100100011000",
			4774 => "0000000001000000001101111100010000",
			4775 => "0000000111000000000110100100001000",
			4776 => "0000000000000000001111001000000100",
			4777 => "00000000101101100100101110011011",
			4778 => "00000000000000000100101110011011",
			4779 => "0000000101000000000110100000000100",
			4780 => "11111110110011100100101110011011",
			4781 => "00000000000000110100101110011011",
			4782 => "0000001101000000000101110000000100",
			4783 => "11111110011100010100101110011011",
			4784 => "00000000000000000100101110011011",
			4785 => "0000001011000000000110110100001100",
			4786 => "0000000000000000000001110100001000",
			4787 => "0000000110000000001101111100000100",
			4788 => "00000000000000000100101110011011",
			4789 => "00000001011001100100101110011011",
			4790 => "00000000000000000100101110011011",
			4791 => "00000000000000000100101110011011",
			4792 => "0000001101000000000010011100000100",
			4793 => "00000000000000000100101110011011",
			4794 => "0000000001000000000001111000001100",
			4795 => "0000001011000000000010001000001000",
			4796 => "0000000011000000000111011000000100",
			4797 => "00000000000000000100101110011011",
			4798 => "11111110100100100100101110011011",
			4799 => "00000000000000000100101110011011",
			4800 => "00000000000000000100101110011011",
			4801 => "0000000101000000001111010000100000",
			4802 => "0000000000000000000101000100001100",
			4803 => "0000001101000000000101110000000100",
			4804 => "00000000000000000100101110011011",
			4805 => "0000000111000000000001101000000100",
			4806 => "00000000000000000100101110011011",
			4807 => "11111111101010110100101110011011",
			4808 => "0000000001000000000100110100001100",
			4809 => "0000000100000000000111011000000100",
			4810 => "00000000000000000100101110011011",
			4811 => "0000001101000000001010001000000100",
			4812 => "00000001001111000100101110011011",
			4813 => "00000000000000000100101110011011",
			4814 => "0000001101000000001010001000000100",
			4815 => "11111111111111110100101110011011",
			4816 => "00000000000000000100101110011011",
			4817 => "0000000001000000000000111100010000",
			4818 => "0000000010000000001100000000001000",
			4819 => "0000000100000000000110111100000100",
			4820 => "11111111100111110100101110011011",
			4821 => "00000000110010110100101110011011",
			4822 => "0000000111000000001111011100000100",
			4823 => "11111110110111010100101110011011",
			4824 => "00000000000000000100101110011011",
			4825 => "0000001101000000001100010100001100",
			4826 => "0000000000000000001010101100001000",
			4827 => "0000001011000000000100010000000100",
			4828 => "00000000000000000100101110011011",
			4829 => "00000001001011000100101110011011",
			4830 => "00000000000000000100101110011011",
			4831 => "0000001100000000001000011000001000",
			4832 => "0000000101000000000011001000000100",
			4833 => "11111111000111010100101110011011",
			4834 => "00000000000000000100101110011011",
			4835 => "0000000001000000000111101000000100",
			4836 => "00000000010001100100101110011011",
			4837 => "00000000000000000100101110011011",
			4838 => "00000000000000000100101110011101",
			4839 => "00000000000000000100101110100001",
			4840 => "0000001100000000001011000000000100",
			4841 => "11111111111111110100101110110101",
			4842 => "0000001100000000000110100100000100",
			4843 => "00000000000001100100101110110101",
			4844 => "00000000000000000100101110110101",
			4845 => "0000001011000000000100010000001000",
			4846 => "0000001011000000000000011100000100",
			4847 => "00000000000000000100101111001001",
			4848 => "11111111111100000100101111001001",
			4849 => "00000000000000000100101111001001",
			4850 => "0000000000000000001100000100001000",
			4851 => "0000000100000000000110110100000100",
			4852 => "00000000000000000100101111011101",
			4853 => "00000000000001100100101111011101",
			4854 => "00000000000000000100101111011101",
			4855 => "0000000000000000001100000100001000",
			4856 => "0000000000000000000011101000000100",
			4857 => "00000000000000000100101111110001",
			4858 => "00000000000000110100101111110001",
			4859 => "00000000000000000100101111110001",
			4860 => "0000000101000000001100100100001000",
			4861 => "0000000101000000000110110100000100",
			4862 => "00000000000000000100110000001101",
			4863 => "00000000000101000100110000001101",
			4864 => "0000000101000000001111010000000100",
			4865 => "11111111111100110100110000001101",
			4866 => "00000000000000000100110000001101",
			4867 => "0000001011000000001011011100000100",
			4868 => "00000000000000000100110000101001",
			4869 => "0000000010000000001100000000001000",
			4870 => "0000000010000000000010000000000100",
			4871 => "00000000000000000100110000101001",
			4872 => "00000000001100110100110000101001",
			4873 => "00000000000000000100110000101001",
			4874 => "0000000010000000001100010000001100",
			4875 => "0000000100000000000111010100001000",
			4876 => "0000000010000000001101000100000100",
			4877 => "00000000000000000100110001001101",
			4878 => "00000000000111010100110001001101",
			4879 => "00000000000000000100110001001101",
			4880 => "0000000010000000001010000100000100",
			4881 => "11111111111010100100110001001101",
			4882 => "00000000000000000100110001001101",
			4883 => "0000000000000000001001101000001100",
			4884 => "0000000010000000001101000100000100",
			4885 => "00000000000000000100110001110001",
			4886 => "0000000010000000001010000100000100",
			4887 => "00000000000100010100110001110001",
			4888 => "00000000000000000100110001110001",
			4889 => "0000000010000000001000101000000100",
			4890 => "11111111111101000100110001110001",
			4891 => "00000000000000000100110001110001",
			4892 => "0000000000000000001100000100001100",
			4893 => "0000000010000000001100000000001000",
			4894 => "0000000010000000001110110100000100",
			4895 => "00000000000000000100110010011101",
			4896 => "00000000001100100100110010011101",
			4897 => "00000000000000000100110010011101",
			4898 => "0000000110000000001000010000001000",
			4899 => "0000000110000000000100110100000100",
			4900 => "00000000000000000100110010011101",
			4901 => "11111111111111010100110010011101",
			4902 => "00000000000000000100110010011101",
			4903 => "0000000000000000000001110100010000",
			4904 => "0000000101000000001100100100001100",
			4905 => "0000000111000000000001101000001000",
			4906 => "0000000111000000001011000000000100",
			4907 => "00000000000000000100110011000001",
			4908 => "00000000001110110100110011000001",
			4909 => "00000000000000000100110011000001",
			4910 => "00000000000000000100110011000001",
			4911 => "00000000000000000100110011000001",
			4912 => "0000001100000000001001110100010000",
			4913 => "0000000100000000001100010000000100",
			4914 => "00000000000000000100110011100101",
			4915 => "0000000110000000001011001100001000",
			4916 => "0000001100000000001010111000000100",
			4917 => "00000000000000000100110011100101",
			4918 => "11111111101101010100110011100101",
			4919 => "00000000000000000100110011100101",
			4920 => "00000000000000000100110011100101",
			4921 => "0000001001000000001111000000001000",
			4922 => "0000001010000000001001100100000100",
			4923 => "00000000000000000100110100010001",
			4924 => "11111111110110100100110100010001",
			4925 => "0000001010000000001001000100001100",
			4926 => "0000001010000000000000001000000100",
			4927 => "00000000000000000100110100010001",
			4928 => "0000001001000000000010101100000100",
			4929 => "00000000000101110100110100010001",
			4930 => "00000000000000000100110100010001",
			4931 => "00000000000000000100110100010001",
			4932 => "0000001011000000001011011100000100",
			4933 => "00000000000000000100110100111101",
			4934 => "0000000101000000001111010000001000",
			4935 => "0000000101000000001100100100000100",
			4936 => "00000000000000000100110100111101",
			4937 => "00000000010001100100110100111101",
			4938 => "0000001011000000001011110100001000",
			4939 => "0000001011000000000010001000000100",
			4940 => "00000000000000000100110100111101",
			4941 => "11111111111000100100110100111101",
			4942 => "00000000000000000100110100111101",
			4943 => "0000001001000000000111101100001100",
			4944 => "0000001001000000001111000000001000",
			4945 => "0000001001000000001111000000000100",
			4946 => "00000000000000000100110101110001",
			4947 => "00000000000100010100110101110001",
			4948 => "11111111111110100100110101110001",
			4949 => "0000000101000000000111111100001100",
			4950 => "0000001001000000000010101100001000",
			4951 => "0000000101000000000010110100000100",
			4952 => "00000000000000000100110101110001",
			4953 => "00000000000111000100110101110001",
			4954 => "00000000000000000100110101110001",
			4955 => "00000000000000000100110101110001",
			4956 => "0000001100000000000100011000001000",
			4957 => "0000001001000000000000001000000100",
			4958 => "11111111111111010100110110100101",
			4959 => "00000000000000000100110110100101",
			4960 => "0000001011000000001011011100000100",
			4961 => "00000000000000000100110110100101",
			4962 => "0000000100000000001101101100001100",
			4963 => "0000001111000000001110110100000100",
			4964 => "00000000000000000100110110100101",
			4965 => "0000000001000000001001011000000100",
			4966 => "00000000000000000100110110100101",
			4967 => "00000000010100000100110110100101",
			4968 => "00000000000000000100110110100101",
			4969 => "0000000000000000000001110100010100",
			4970 => "0000000101000000001100100100010000",
			4971 => "0000001001000000001010100000001100",
			4972 => "0000000101000000000110110100000100",
			4973 => "00000000000000000100110111010001",
			4974 => "0000000000000000001111001000000100",
			4975 => "00000000001101110100110111010001",
			4976 => "00000000000000000100110111010001",
			4977 => "00000000000000000100110111010001",
			4978 => "00000000000000000100110111010001",
			4979 => "00000000000000000100110111010001",
			4980 => "0000001100000000001001110100010100",
			4981 => "0000000100000000001100010000000100",
			4982 => "00000000000000000100110111111101",
			4983 => "0000000110000000001011001100001100",
			4984 => "0000001100000000001010111000000100",
			4985 => "00000000000000000100110111111101",
			4986 => "0000000111000000001001001000000100",
			4987 => "00000000000000000100110111111101",
			4988 => "11111111101111010100110111111101",
			4989 => "00000000000000000100110111111101",
			4990 => "00000000000000000100110111111101",
			4991 => "0000000000000000001001101000010100",
			4992 => "0000001111000000000111011000000100",
			4993 => "00000000000000000100111001000001",
			4994 => "0000000000000000000001010100000100",
			4995 => "00000000000000000100111001000001",
			4996 => "0000001100000000000110100100001000",
			4997 => "0000001011000000000101100100000100",
			4998 => "00000000000000000100111001000001",
			4999 => "00000000101101000100111001000001",
			5000 => "00000000000000000100111001000001",
			5001 => "0000001110000000000111010100000100",
			5002 => "11111111110110010100111001000001",
			5003 => "0000001000000000000101000100001000",
			5004 => "0000001000000000000001010000000100",
			5005 => "00000000000000000100111001000001",
			5006 => "00000000000111010100111001000001",
			5007 => "00000000000000000100111001000001",
			5008 => "0000001100000000001001110100010000",
			5009 => "0000000100000000001100010000000100",
			5010 => "00000000000000000100111010000101",
			5011 => "0000001110000000001100111000001000",
			5012 => "0000001011000000000101100100000100",
			5013 => "00000000000000000100111010000101",
			5014 => "11111111101000110100111010000101",
			5015 => "00000000000000000100111010000101",
			5016 => "0000000010000000000110111000010000",
			5017 => "0000000000000000000001010100000100",
			5018 => "00000000000000000100111010000101",
			5019 => "0000001011000000000010001000000100",
			5020 => "00000000000000000100111010000101",
			5021 => "0000001101000000000010000100000100",
			5022 => "00000000001100110100111010000101",
			5023 => "00000000000000000100111010000101",
			5024 => "00000000000000000100111010000101",
			5025 => "0000000000000000000111000100011000",
			5026 => "0000001001000000001111000000000100",
			5027 => "00000000000000000100111011000001",
			5028 => "0000001101000000001110000100000100",
			5029 => "00000000000000000100111011000001",
			5030 => "0000001101000000001010001000001100",
			5031 => "0000001010000000000000001000000100",
			5032 => "00000000000000000100111011000001",
			5033 => "0000000111000000000110100100000100",
			5034 => "00000000000000000100111011000001",
			5035 => "00000000100000000100111011000001",
			5036 => "00000000000000000100111011000001",
			5037 => "0000000110000000001000010000000100",
			5038 => "11111111111011100100111011000001",
			5039 => "00000000000000000100111011000001",
			5040 => "0000000100000000000001011100011000",
			5041 => "0000001010000000000000001000000100",
			5042 => "00000000000000000100111011111101",
			5043 => "0000000001000000001101111100010000",
			5044 => "0000000001000000001001011000000100",
			5045 => "00000000000000000100111011111101",
			5046 => "0000001011000000000000011100000100",
			5047 => "00000000000000000100111011111101",
			5048 => "0000001000000000001100011100000100",
			5049 => "00000000010110100100111011111101",
			5050 => "00000000000000000100111011111101",
			5051 => "00000000000000000100111011111101",
			5052 => "0000000110000000000100111100000100",
			5053 => "11111111111101110100111011111101",
			5054 => "00000000000000000100111011111101",
			5055 => "0000001110000000001100000000001000",
			5056 => "0000001101000000001001010100000100",
			5057 => "00000000000000000100111100111001",
			5058 => "11111111111111100100111100111001",
			5059 => "0000001101000000000011001000010100",
			5060 => "0000001001000000000100111100000100",
			5061 => "00000000000000000100111100111001",
			5062 => "0000001110000000000010010100001100",
			5063 => "0000001101000000001110000100000100",
			5064 => "00000000000000000100111100111001",
			5065 => "0000001001000000000010101100000100",
			5066 => "00000000001011000100111100111001",
			5067 => "00000000000000000100111100111001",
			5068 => "00000000000000000100111100111001",
			5069 => "00000000000000000100111100111001",
			5070 => "0000000110000000001101111100001000",
			5071 => "0000001100000000000100011000000100",
			5072 => "00000000000000000100111101110101",
			5073 => "00000000010110110100111101110101",
			5074 => "0000000111000000001000011000010100",
			5075 => "0000000101000000001100100100000100",
			5076 => "00000000000000000100111101110101",
			5077 => "0000001100000000001001110100001100",
			5078 => "0000001001000000001010100100001000",
			5079 => "0000001101000000000010011100000100",
			5080 => "00000000000000000100111101110101",
			5081 => "11111111101011000100111101110101",
			5082 => "00000000000000000100111101110101",
			5083 => "00000000000000000100111101110101",
			5084 => "00000000000000000100111101110101",
			5085 => "0000000000000000000001110100011000",
			5086 => "0000000101000000001100100100010100",
			5087 => "0000001001000000001010100000010000",
			5088 => "0000000101000000000110100000000100",
			5089 => "00000000000000000100111110101001",
			5090 => "0000001001000000001111000000000100",
			5091 => "00000000000000000100111110101001",
			5092 => "0000000000000000001111001000000100",
			5093 => "00000000010110100100111110101001",
			5094 => "00000000000000000100111110101001",
			5095 => "00000000000000000100111110101001",
			5096 => "00000000000000000100111110101001",
			5097 => "00000000000000000100111110101001",
			5098 => "0000000101000000001111010000011000",
			5099 => "0000001100000000000100011000000100",
			5100 => "00000000000000000100111111011101",
			5101 => "0000000000000000000010101000010000",
			5102 => "0000001100000000001001001000001100",
			5103 => "0000000111000000000110100100000100",
			5104 => "00000000000000000100111111011101",
			5105 => "0000000111000000001111011100000100",
			5106 => "00000000011010010100111111011101",
			5107 => "00000000000000000100111111011101",
			5108 => "00000000000000000100111111011101",
			5109 => "00000000000000000100111111011101",
			5110 => "00000000000000000100111111011101",
			5111 => "0000000001000000000000111100010000",
			5112 => "0000001110000000001110110100000100",
			5113 => "00000000000000000101000000101001",
			5114 => "0000000101000000000101110000001000",
			5115 => "0000001101000000000101110000000100",
			5116 => "00000000000000000101000000101001",
			5117 => "11111111110110010101000000101001",
			5118 => "00000000000000000101000000101001",
			5119 => "0000001100000000000100011000000100",
			5120 => "00000000000000000101000000101001",
			5121 => "0000000000000000000001110100010000",
			5122 => "0000001110000000001100000000000100",
			5123 => "00000000000000000101000000101001",
			5124 => "0000000001000000000100110100001000",
			5125 => "0000000101000000000110100000000100",
			5126 => "00000000000000000101000000101001",
			5127 => "00000000011011100101000000101001",
			5128 => "00000000000000000101000000101001",
			5129 => "00000000000000000101000000101001",
			5130 => "0000000100000000000111010100010100",
			5131 => "0000001000000000001000100100000100",
			5132 => "00000000000000000101000010001101",
			5133 => "0000001111000000001111010100001100",
			5134 => "0000001100000000000111001000000100",
			5135 => "00000000000000000101000010001101",
			5136 => "0000001111000000000110010000000100",
			5137 => "00000000000000000101000010001101",
			5138 => "00000000001110100101000010001101",
			5139 => "00000000000000000101000010001101",
			5140 => "0000000110000000000100111100010000",
			5141 => "0000000111000000000000011100001100",
			5142 => "0000001000000000001000010100000100",
			5143 => "00000000000000000101000010001101",
			5144 => "0000000110000000001111000000000100",
			5145 => "11111111100000110101000010001101",
			5146 => "00000000000000000101000010001101",
			5147 => "00000000000000000101000010001101",
			5148 => "0000000000000000001010101100001100",
			5149 => "0000000001000000001010011000001000",
			5150 => "0000001001000000001010100000000100",
			5151 => "00000000000000000101000010001101",
			5152 => "00000000001110000101000010001101",
			5153 => "00000000000000000101000010001101",
			5154 => "00000000000000000101000010001101",
			5155 => "0000000000000000001100000100011000",
			5156 => "0000001010000000000000001000010000",
			5157 => "0000001000000000000111110100000100",
			5158 => "00000000000000000101000011111001",
			5159 => "0000000110000000000100110100001000",
			5160 => "0000001111000000001001100000000100",
			5161 => "00000000000000000101000011111001",
			5162 => "11111111101101100101000011111001",
			5163 => "00000000000000000101000011111001",
			5164 => "0000001111000000000110010000000100",
			5165 => "00000000000000000101000011111001",
			5166 => "00000000000111010101000011111001",
			5167 => "0000001010000000000010101100001100",
			5168 => "0000001011000000000101110100001000",
			5169 => "0000000110000000001101111100000100",
			5170 => "00000000000000000101000011111001",
			5171 => "11111111101000010101000011111001",
			5172 => "00000000000000000101000011111001",
			5173 => "0000001010000000001000100100010000",
			5174 => "0000000010000000001101101100001100",
			5175 => "0000001000000000000101000100001000",
			5176 => "0000000010000000001100000000000100",
			5177 => "00000000000000000101000011111001",
			5178 => "00000000001011010101000011111001",
			5179 => "00000000000000000101000011111001",
			5180 => "00000000000000000101000011111001",
			5181 => "00000000000000000101000011111001",
			5182 => "0000000100000000000001011100100000",
			5183 => "0000001000000000001000100100001000",
			5184 => "0000000001000000001001011000000100",
			5185 => "00000000000000000101000101001101",
			5186 => "11111111111111110101000101001101",
			5187 => "0000000111000000000110100100000100",
			5188 => "00000000000000000101000101001101",
			5189 => "0000000001000000001001011000000100",
			5190 => "00000000000000000101000101001101",
			5191 => "0000000111000000001000011000001100",
			5192 => "0000000001000000000111101000001000",
			5193 => "0000001101000000000001000000000100",
			5194 => "00000000000000000101000101001101",
			5195 => "00000000010111110101000101001101",
			5196 => "00000000000000000101000101001101",
			5197 => "00000000000000000101000101001101",
			5198 => "0000000001000000001100011000001000",
			5199 => "0000000111000000000001011000000100",
			5200 => "11111111110000100101000101001101",
			5201 => "00000000000000000101000101001101",
			5202 => "00000000000000000101000101001101",
			5203 => "0000001011000000001011011100001100",
			5204 => "0000001110000000000111011000001000",
			5205 => "0000000011000000001010000100000100",
			5206 => "11111111110011010101000110011001",
			5207 => "00000000000000000101000110011001",
			5208 => "00000000000000000101000110011001",
			5209 => "0000000100000000001101101100011000",
			5210 => "0000000111000000000110100100000100",
			5211 => "00000000000000000101000110011001",
			5212 => "0000000001000000001001011000000100",
			5213 => "00000000000000000101000110011001",
			5214 => "0000000000000000000101000100000100",
			5215 => "00000000000000000101000110011001",
			5216 => "0000000100000000000111011000000100",
			5217 => "00000000000000000101000110011001",
			5218 => "0000000010000000001110110100000100",
			5219 => "00000000000000000101000110011001",
			5220 => "00000000011111110101000110011001",
			5221 => "00000000000000000101000110011001",
			5222 => "0000000100000000001101101100011100",
			5223 => "0000000001000000001001011000000100",
			5224 => "00000000000000000101000111011101",
			5225 => "0000001101000000001110000100000100",
			5226 => "00000000000000000101000111011101",
			5227 => "0000000011000000001000100000010000",
			5228 => "0000001001000000001111000000000100",
			5229 => "00000000000000000101000111011101",
			5230 => "0000001111000000001100000000000100",
			5231 => "00000000000000000101000111011101",
			5232 => "0000000001000000001101111100000100",
			5233 => "00000000011000000101000111011101",
			5234 => "00000000000000000101000111011101",
			5235 => "00000000000000000101000111011101",
			5236 => "0000001001000000001010100000000100",
			5237 => "11111111111000000101000111011101",
			5238 => "00000000000000000101000111011101",
			5239 => "0000001111000000001100000000001100",
			5240 => "0000001010000000001010100000001000",
			5241 => "0000000111000000000110100100000100",
			5242 => "00000000000000000101001001001001",
			5243 => "11111111100100100101001001001001",
			5244 => "00000000000000000101001001001001",
			5245 => "0000001100000000001000000000011000",
			5246 => "0000001010000000000010101100001100",
			5247 => "0000000111000000001000011000001000",
			5248 => "0000001100000000001010111000000100",
			5249 => "00000000000000000101001001001001",
			5250 => "11111111101000100101001001001001",
			5251 => "00000000000000000101001001001001",
			5252 => "0000001010000000001000100100001000",
			5253 => "0000000111000000001001001000000100",
			5254 => "00000000000000000101001001001001",
			5255 => "00000000001000110101001001001001",
			5256 => "00000000000000000101001001001001",
			5257 => "0000001100000000000110100100010000",
			5258 => "0000001101000000001100010100001100",
			5259 => "0000000001000000000000111100000100",
			5260 => "00000000000000000101001001001001",
			5261 => "0000000000000000000111000000000100",
			5262 => "00000000101101100101001001001001",
			5263 => "00000000000000000101001001001001",
			5264 => "00000000000000000101001001001001",
			5265 => "00000000000000000101001001001001",
			5266 => "0000000101000000000110100000001000",
			5267 => "0000001110000000000111010100000100",
			5268 => "11111111110001110101001010101101",
			5269 => "00000000000000000101001010101101",
			5270 => "0000001001000000001001111100011000",
			5271 => "0000000010000000001100010000001100",
			5272 => "0000001110000000000110010000000100",
			5273 => "00000000000000000101001010101101",
			5274 => "0000000010000000000110010000000100",
			5275 => "00000000000000000101001010101101",
			5276 => "00000000000110100101001010101101",
			5277 => "0000001110000000001010000100001000",
			5278 => "0000000010000000001100000000000100",
			5279 => "00000000000000000101001010101101",
			5280 => "11111111110010110101001010101101",
			5281 => "00000000000000000101001010101101",
			5282 => "0000000010000000000110111000010000",
			5283 => "0000001001000000000010101100001100",
			5284 => "0000001110000000001100010000000100",
			5285 => "00000000000000000101001010101101",
			5286 => "0000000111000000001001001000000100",
			5287 => "00000000000000000101001010101101",
			5288 => "00000000010011110101001010101101",
			5289 => "00000000000000000101001010101101",
			5290 => "00000000000000000101001010101101",
			5291 => "0000001001000000001111000000001100",
			5292 => "0000000110000000001101111100000100",
			5293 => "00000000000000000101001100000001",
			5294 => "0000001010000000000000001000000100",
			5295 => "00000000000000000101001100000001",
			5296 => "11111111110111110101001100000001",
			5297 => "0000000000000000000001110100011100",
			5298 => "0000000111000000000110100100000100",
			5299 => "00000000000000000101001100000001",
			5300 => "0000001100000000001001001000010000",
			5301 => "0000001101000000001010001000001100",
			5302 => "0000000101000000001001010000001000",
			5303 => "0000001000000000001000100100000100",
			5304 => "00000000000000000101001100000001",
			5305 => "00000000011101010101001100000001",
			5306 => "00000000000000000101001100000001",
			5307 => "00000000000000000101001100000001",
			5308 => "0000001100000000001001110100000100",
			5309 => "11111111111111100101001100000001",
			5310 => "00000000000000000101001100000001",
			5311 => "00000000000000000101001100000001",
			5312 => "0000001110000000000111010100011100",
			5313 => "0000001011000000000101110100011000",
			5314 => "0000000100000000000110010000000100",
			5315 => "00000000000000000101001100111101",
			5316 => "0000001010000000000010101100010000",
			5317 => "0000000111000000001001001000000100",
			5318 => "00000000000000000101001100111101",
			5319 => "0000000101000000001111010000001000",
			5320 => "0000000111000000001111011100000100",
			5321 => "11111111101011000101001100111101",
			5322 => "00000000000000000101001100111101",
			5323 => "00000000000000000101001100111101",
			5324 => "00000000000000000101001100111101",
			5325 => "00000000000000000101001100111101",
			5326 => "00000000000000000101001100111101",
			5327 => "0000001001000000001111000000000100",
			5328 => "00000000000000000101001101111001",
			5329 => "0000000100000000000101000000011000",
			5330 => "0000001100000000000100011000000100",
			5331 => "00000000000000000101001101111001",
			5332 => "0000000101000000001110010000010000",
			5333 => "0000001010000000000000001000000100",
			5334 => "00000000000000000101001101111001",
			5335 => "0000001001000000000010101100001000",
			5336 => "0000001011000000000100000100000100",
			5337 => "00000000000000000101001101111001",
			5338 => "00000000010000010101001101111001",
			5339 => "00000000000000000101001101111001",
			5340 => "00000000000000000101001101111001",
			5341 => "00000000000000000101001101111001",
			5342 => "0000000000000000000010101000011100",
			5343 => "0000001001000000001111000000000100",
			5344 => "00000000000000000101001110110101",
			5345 => "0000000111000000000110100100000100",
			5346 => "00000000000000000101001110110101",
			5347 => "0000000000000000000001010100000100",
			5348 => "00000000000000000101001110110101",
			5349 => "0000000001000000001010011000001100",
			5350 => "0000001100000000001010111000000100",
			5351 => "00000000000000000101001110110101",
			5352 => "0000000001000000000000111100000100",
			5353 => "00000000000000000101001110110101",
			5354 => "00000000100001100101001110110101",
			5355 => "00000000000000000101001110110101",
			5356 => "00000000000000000101001110110101",
			5357 => "0000001001000000001111000000000100",
			5358 => "00000000000000000101010000000001",
			5359 => "0000000100000000001111100100011000",
			5360 => "0000000101000000001111010000010100",
			5361 => "0000001101000000001010001000010000",
			5362 => "0000001100000000001001001000001100",
			5363 => "0000000111000000000110100100000100",
			5364 => "00000000000000000101010000000001",
			5365 => "0000001010000000000000001000000100",
			5366 => "00000000000000000101010000000001",
			5367 => "00000000100000110101010000000001",
			5368 => "00000000000000000101010000000001",
			5369 => "00000000000000000101010000000001",
			5370 => "00000000000000000101010000000001",
			5371 => "0000001001000000000111101100001000",
			5372 => "0000000110000000001101011000000100",
			5373 => "00000000000000000101010000000001",
			5374 => "11111111110101000101010000000001",
			5375 => "00000000000000000101010000000001",
			5376 => "0000000100000000001111100100011000",
			5377 => "0000001111000000001110110100000100",
			5378 => "00000000000000000101010001110101",
			5379 => "0000000011000000000000010000010000",
			5380 => "0000000110000000000100110100000100",
			5381 => "00000000000000000101010001110101",
			5382 => "0000000111000000000110100100000100",
			5383 => "00000000000000000101010001110101",
			5384 => "0000001010000000000011101000000100",
			5385 => "00000000101011100101010001110101",
			5386 => "00000000000000000101010001110101",
			5387 => "00000000000000000101010001110101",
			5388 => "0000000011000000001111100100010000",
			5389 => "0000001100000000001010111000000100",
			5390 => "00000000000000000101010001110101",
			5391 => "0000000101000000000010110100000100",
			5392 => "00000000000000000101010001110101",
			5393 => "0000000101000000000111100000000100",
			5394 => "11111111011111010101010001110101",
			5395 => "00000000000000000101010001110101",
			5396 => "0000000001000000000001000100000100",
			5397 => "00000000000000000101010001110101",
			5398 => "0000001111000000001110000000001100",
			5399 => "0000000001000000001010011000001000",
			5400 => "0000001010000000001001000100000100",
			5401 => "00000000001010000101010001110101",
			5402 => "00000000000000000101010001110101",
			5403 => "00000000000000000101010001110101",
			5404 => "00000000000000000101010001110101",
			5405 => "0000000100000000001011101100110000",
			5406 => "0000001101000000000101110000011000",
			5407 => "0000000111000000000110100100000100",
			5408 => "00000000000000000101010100000001",
			5409 => "0000001001000000001111000000000100",
			5410 => "00000000000000000101010100000001",
			5411 => "0000001011000000000110110100001100",
			5412 => "0000001010000000000000001000000100",
			5413 => "00000000000000000101010100000001",
			5414 => "0000001101000000001110000100000100",
			5415 => "00000000000000000101010100000001",
			5416 => "00000000101001000101010100000001",
			5417 => "00000000000000000101010100000001",
			5418 => "0000001011000000000110110100001100",
			5419 => "0000000011000000000000010000001000",
			5420 => "0000001111000000001001100000000100",
			5421 => "00000000000000000101010100000001",
			5422 => "11111111110100000101010100000001",
			5423 => "00000000000000000101010100000001",
			5424 => "0000000011000000000111010100001000",
			5425 => "0000001111000000001100000000000100",
			5426 => "00000000000000000101010100000001",
			5427 => "00000000011011110101010100000001",
			5428 => "00000000000000000101010100000001",
			5429 => "0000000011000000001111100100001100",
			5430 => "0000001110000000001000001100001000",
			5431 => "0000000000000000001011010100000100",
			5432 => "00000000000000000101010100000001",
			5433 => "11111111011010100101010100000001",
			5434 => "00000000000000000101010100000001",
			5435 => "0000000000000000000111000100001000",
			5436 => "0000000000000000001011010100000100",
			5437 => "00000000000000000101010100000001",
			5438 => "00000000010100100101010100000001",
			5439 => "00000000000000000101010100000001",
			5440 => "0000000000000000000001110100101000",
			5441 => "0000001001000000001111000000001000",
			5442 => "0000000111000000001000011000000100",
			5443 => "11111110011010100101010110000101",
			5444 => "00000001001111100101010110000101",
			5445 => "0000001101000000000001000000001000",
			5446 => "0000000010000000000110010000000100",
			5447 => "00000011000011100101010110000101",
			5448 => "11111110011000100101010110000101",
			5449 => "0000001101000000000110010000010100",
			5450 => "0000001000000000000101000100001100",
			5451 => "0000000110000000001101111100000100",
			5452 => "11111110100111100101010110000101",
			5453 => "0000000100000000000001011100000100",
			5454 => "00000100010011010101010110000101",
			5455 => "00000011000101000101010110000101",
			5456 => "0000000100000000000110111000000100",
			5457 => "00000100101101010101010110000101",
			5458 => "00001001101110100101010110000101",
			5459 => "11111110011000000101010110000101",
			5460 => "0000000000000000001010101100010100",
			5461 => "0000001000000000000001010100001100",
			5462 => "0000001000000000000001010100000100",
			5463 => "11111110010110110101010110000101",
			5464 => "0000000100000000001000000100000100",
			5465 => "00000001111011100101010110000101",
			5466 => "11111110011110100101010110000101",
			5467 => "0000000110000000001000010000000100",
			5468 => "11111110110000100101010110000101",
			5469 => "00000111100001100101010110000101",
			5470 => "0000000000000000001010101100000100",
			5471 => "11111110101100000101010110000101",
			5472 => "11111110010110100101010110000101",
			5473 => "0000001001000000000100111100010100",
			5474 => "0000001010000000001010100000001100",
			5475 => "0000000011000000000111010100001000",
			5476 => "0000000011000000000111100000000100",
			5477 => "00000000000000000101011000010001",
			5478 => "00000000000010100101011000010001",
			5479 => "00000000000000000101011000010001",
			5480 => "0000000001000000000000111100000100",
			5481 => "11111111101000000101011000010001",
			5482 => "00000000000000000101011000010001",
			5483 => "0000001111000000001111010100010000",
			5484 => "0000000000000000001001101000001100",
			5485 => "0000001101000000001010001000001000",
			5486 => "0000001101000000000111100000000100",
			5487 => "00000000000000000101011000010001",
			5488 => "00000000101001110101011000010001",
			5489 => "00000000000000000101011000010001",
			5490 => "00000000000000000101011000010001",
			5491 => "0000000011000000001010000100001100",
			5492 => "0000001111000000001010000100001000",
			5493 => "0000000101000000001110101000000100",
			5494 => "00000000000000000101011000010001",
			5495 => "11111111011110110101011000010001",
			5496 => "00000000000000000101011000010001",
			5497 => "0000000000000000000001110100010000",
			5498 => "0000000000000000001001101000000100",
			5499 => "00000000000000000101011000010001",
			5500 => "0000000101000000001101000100000100",
			5501 => "00000000000000000101011000010001",
			5502 => "0000001001000000000101010000000100",
			5503 => "00000000000000000101011000010001",
			5504 => "00000000101000000101011000010001",
			5505 => "0000000011000000001000101000000100",
			5506 => "11111111111101100101011000010001",
			5507 => "00000000000000000101011000010001",
			5508 => "0000000100000000001101101100101000",
			5509 => "0000001111000000001010000100100100",
			5510 => "0000000111000000000001101000010100",
			5511 => "0000000100000000001100010000000100",
			5512 => "00000000000000000101011001111101",
			5513 => "0000001101000000000111111100001100",
			5514 => "0000000111000000001001001000000100",
			5515 => "00000000000000000101011001111101",
			5516 => "0000001011000000000000011100000100",
			5517 => "00000000000000000101011001111101",
			5518 => "11111111101001100101011001111101",
			5519 => "00000000000000000101011001111101",
			5520 => "0000000000000000000101000100000100",
			5521 => "00000000000000000101011001111101",
			5522 => "0000001001000000001111000000000100",
			5523 => "00000000000000000101011001111101",
			5524 => "0000000111000000001111011100000100",
			5525 => "00000000011010000101011001111101",
			5526 => "00000000000000000101011001111101",
			5527 => "00000000101101100101011001111101",
			5528 => "0000001001000000001010100000001100",
			5529 => "0000001100000000001011011100001000",
			5530 => "0000001000000000000001010000000100",
			5531 => "00000000000000000101011001111101",
			5532 => "11111111101000010101011001111101",
			5533 => "00000000000000000101011001111101",
			5534 => "00000000000000000101011001111101",
			5535 => "0000000100000000001011101100101100",
			5536 => "0000001011000000000101100100010100",
			5537 => "0000000010000000001111010100010000",
			5538 => "0000001001000000000101010000000100",
			5539 => "00000000000000000101011100010001",
			5540 => "0000001100000000001101010100000100",
			5541 => "00000000000000000101011100010001",
			5542 => "0000001101000000001110000100000100",
			5543 => "00000000000000000101011100010001",
			5544 => "11111111011110100101011100010001",
			5545 => "00000000000000000101011100010001",
			5546 => "0000001101000000000101001000000100",
			5547 => "00000000000000000101011100010001",
			5548 => "0000000001000000001001011000000100",
			5549 => "00000000000000000101011100010001",
			5550 => "0000000010000000001000001100001100",
			5551 => "0000001101000000001010001000001000",
			5552 => "0000001000000000001000100100000100",
			5553 => "00000000000000000101011100010001",
			5554 => "00000000100100010101011100010001",
			5555 => "00000000000000000101011100010001",
			5556 => "00000000000000000101011100010001",
			5557 => "0000000110000000001001100100001100",
			5558 => "0000001100000000001001110100001000",
			5559 => "0000000000000000001011010100000100",
			5560 => "00000000000000000101011100010001",
			5561 => "11111111010010010101011100010001",
			5562 => "00000000000000000101011100010001",
			5563 => "0000000000000000000001110100001100",
			5564 => "0000000010000000001101101100001000",
			5565 => "0000001111000000000110101100000100",
			5566 => "00000000000000000101011100010001",
			5567 => "00000000011100110101011100010001",
			5568 => "00000000000000000101011100010001",
			5569 => "0000001000000000000001110000000100",
			5570 => "00000000000000000101011100010001",
			5571 => "00000000000000000101011100010001",
			5572 => "0000000100000000001011101100110000",
			5573 => "0000000111000000001000011000011000",
			5574 => "0000001100000000001010111000000100",
			5575 => "00000000000000000101011110000101",
			5576 => "0000001001000000000111101100010000",
			5577 => "0000000001000000001001011000000100",
			5578 => "00000000000000000101011110000101",
			5579 => "0000001100000000001001001000001000",
			5580 => "0000001011000000000111010000000100",
			5581 => "00000000000000000101011110000101",
			5582 => "00000000100000010101011110000101",
			5583 => "00000000000000000101011110000101",
			5584 => "00000000000000000101011110000101",
			5585 => "0000001011000000000100010000010100",
			5586 => "0000000101000000001001010000010000",
			5587 => "0000000101000000001100100100000100",
			5588 => "00000000000000000101011110000101",
			5589 => "0000001100000000000100011000000100",
			5590 => "00000000000000000101011110000101",
			5591 => "0000001100000000001001110100000100",
			5592 => "11111111100011110101011110000101",
			5593 => "00000000000000000101011110000101",
			5594 => "00000000000000000101011110000101",
			5595 => "00000000000000000101011110000101",
			5596 => "0000001100000000001001110100001000",
			5597 => "0000000110000000000100111100000100",
			5598 => "11111111011101010101011110000101",
			5599 => "00000000000000000101011110000101",
			5600 => "00000000000000000101011110000101",
			5601 => "0000001101000000000101110000011000",
			5602 => "0000000000000000001111001000010000",
			5603 => "0000001001000000001111000000000100",
			5604 => "00000000000000000101100000011001",
			5605 => "0000001011000000000110110100001000",
			5606 => "0000001101000000000001000000000100",
			5607 => "00000000000000000101100000011001",
			5608 => "00000000110001110101100000011001",
			5609 => "00000000000000000101100000011001",
			5610 => "0000000011000000001000100000000100",
			5611 => "11111111110110000101100000011001",
			5612 => "00000000000000000101100000011001",
			5613 => "0000000101000000000111100000001100",
			5614 => "0000001000000000000001010000001000",
			5615 => "0000001100000000000100011000000100",
			5616 => "00000000000000000101100000011001",
			5617 => "11111111010011000101100000011001",
			5618 => "00000000000000000101100000011001",
			5619 => "0000001101000000001010001000010100",
			5620 => "0000001100000000000100011000000100",
			5621 => "00000000000000000101100000011001",
			5622 => "0000000010000000001110110100000100",
			5623 => "00000000000000000101100000011001",
			5624 => "0000001011000000000101110100001000",
			5625 => "0000000000000000001010101100000100",
			5626 => "00000000110011110101100000011001",
			5627 => "00000000000000000101100000011001",
			5628 => "00000000000000000101100000011001",
			5629 => "0000000011000000001011111000000100",
			5630 => "00000000000000000101100000011001",
			5631 => "0000001100000000001000011000001100",
			5632 => "0000000101000000001111010000000100",
			5633 => "00000000000000000101100000011001",
			5634 => "0000000101000000000011001000000100",
			5635 => "11111111011101100101100000011001",
			5636 => "00000000000000000101100000011001",
			5637 => "00000000000000000101100000011001",
			5638 => "0000000110000000001101111100010000",
			5639 => "0000001100000000000100011000000100",
			5640 => "00000000000000000101100010100101",
			5641 => "0000001100000000001001110100001000",
			5642 => "0000000001000000000000111100000100",
			5643 => "00000000011000010101100010100101",
			5644 => "00000000000000000101100010100101",
			5645 => "00000000000000000101100010100101",
			5646 => "0000000111000000001000011000100000",
			5647 => "0000001001000000000100101100010100",
			5648 => "0000000101000000001100100100000100",
			5649 => "00000000000000000101100010100101",
			5650 => "0000001101000000001001011100001100",
			5651 => "0000001100000000000100011000000100",
			5652 => "00000000000000000101100010100101",
			5653 => "0000001101000000000010011100000100",
			5654 => "00000000000000000101100010100101",
			5655 => "11111111011001010101100010100101",
			5656 => "00000000000000000101100010100101",
			5657 => "0000000001000000001101111100001000",
			5658 => "0000000111000000001000000000000100",
			5659 => "00000000000000000101100010100101",
			5660 => "00000000000111100101100010100101",
			5661 => "00000000000000000101100010100101",
			5662 => "0000001100000000001011000000000100",
			5663 => "00000000000000000101100010100101",
			5664 => "0000001101000000000110010000010000",
			5665 => "0000001100000000000001101000001100",
			5666 => "0000001101000000001100010100001000",
			5667 => "0000000110000000000101010000000100",
			5668 => "00000000100110010101100010100101",
			5669 => "00000000000000000101100010100101",
			5670 => "00000000000000000101100010100101",
			5671 => "00000000000000000101100010100101",
			5672 => "00000000000000000101100010100101",
			5673 => "0000000000000000000010101000111100",
			5674 => "0000000001000000001001011000010000",
			5675 => "0000000110000000000000111100001000",
			5676 => "0000001111000000001010011100000100",
			5677 => "11111110101000110101100100111001",
			5678 => "00000010111001000101100100111001",
			5679 => "0000001001000000001111000000000100",
			5680 => "11111110010101100101100100111001",
			5681 => "00000000000000000101100100111001",
			5682 => "0000001101000000000110010000100100",
			5683 => "0000001101000000001110000100001100",
			5684 => "0000000000000000000001010100000100",
			5685 => "00000001110110010101100100111001",
			5686 => "0000000101000000001101000100000100",
			5687 => "11111110010001110101100100111001",
			5688 => "00000000010010100101100100111001",
			5689 => "0000001010000000000000001000001100",
			5690 => "0000000011000000000010000100001000",
			5691 => "0000001000000000000111110100000100",
			5692 => "00000000000000000101100100111001",
			5693 => "00000000111001110101100100111001",
			5694 => "11111110011011100101100100111001",
			5695 => "0000000110000000000100111100001000",
			5696 => "0000000000000000000110001000000100",
			5697 => "00000001011111100101100100111001",
			5698 => "00000000101000100101100100111001",
			5699 => "00000011000101000101100100111001",
			5700 => "0000000111000000000100010000000100",
			5701 => "11111110011010100101100100111001",
			5702 => "00000000111100010101100100111001",
			5703 => "0000000000000000001010101100001100",
			5704 => "0000001000000000000001010100000100",
			5705 => "11111110011010110101100100111001",
			5706 => "0000000110000000001000010000000100",
			5707 => "00000000000000000101100100111001",
			5708 => "00000010100000100101100100111001",
			5709 => "11111110011001000101100100111001",
			5710 => "0000001111000000001100000000001100",
			5711 => "0000001001000000000100111100001000",
			5712 => "0000000001000000000000111100000100",
			5713 => "11111111100101110101100111000101",
			5714 => "00000000000000000101100111000101",
			5715 => "00000000000000000101100111000101",
			5716 => "0000001100000000001000000000100100",
			5717 => "0000000110000000001011001100010100",
			5718 => "0000000111000000001000011000010000",
			5719 => "0000000101000000001110101000000100",
			5720 => "00000000000000000101100111000101",
			5721 => "0000000110000000001101111100000100",
			5722 => "00000000000000000101100111000101",
			5723 => "0000001100000000000100011000000100",
			5724 => "00000000000000000101100111000101",
			5725 => "11111111011011110101100111000101",
			5726 => "00000000000000000101100111000101",
			5727 => "0000000111000000000001101000001100",
			5728 => "0000000000000000000001110100001000",
			5729 => "0000000111000000001001001000000100",
			5730 => "00000000000000000101100111000101",
			5731 => "00000000001010110101100111000101",
			5732 => "00000000000000000101100111000101",
			5733 => "00000000000000000101100111000101",
			5734 => "0000001101000000000110010000010100",
			5735 => "0000000001000000001001011000000100",
			5736 => "00000000000000000101100111000101",
			5737 => "0000001100000000000110100100001100",
			5738 => "0000001101000000001100010100001000",
			5739 => "0000001110000000001110110100000100",
			5740 => "00000000000000000101100111000101",
			5741 => "00000000101010110101100111000101",
			5742 => "00000000000000000101100111000101",
			5743 => "00000000000000000101100111000101",
			5744 => "00000000000000000101100111000101",
			5745 => "0000001001000000001001111100101100",
			5746 => "0000000000000000001100000100100100",
			5747 => "0000001010000000001010100000011100",
			5748 => "0000001101000000000101110000010000",
			5749 => "0000000101000000000111100000001100",
			5750 => "0000000001000000001101101000000100",
			5751 => "00000000000000000101101001111001",
			5752 => "0000000011000000001100000000000100",
			5753 => "00000000010110110101101001111001",
			5754 => "00000000000000000101101001111001",
			5755 => "00000000000000000101101001111001",
			5756 => "0000001101000000000111111100001000",
			5757 => "0000000010000000000110010000000100",
			5758 => "00000000000000000101101001111001",
			5759 => "11111111010100000101101001111001",
			5760 => "00000000000000000101101001111001",
			5761 => "0000000001000000000000111100000100",
			5762 => "00000000000000000101101001111001",
			5763 => "00000000101100010101101001111001",
			5764 => "0000001100000000001000011000000100",
			5765 => "11111111010001010101101001111001",
			5766 => "00000000000000000101101001111001",
			5767 => "0000000000000000001111001000001100",
			5768 => "0000000011000000000110111100000100",
			5769 => "00000000000000000101101001111001",
			5770 => "0000000101000000000110100000000100",
			5771 => "00000000000000000101101001111001",
			5772 => "00000001000111010101101001111001",
			5773 => "0000001110000000001100111000010000",
			5774 => "0000000111000000001000011000001100",
			5775 => "0000001100000000001010111000000100",
			5776 => "00000000000000000101101001111001",
			5777 => "0000000110000000001000010000000100",
			5778 => "11111111011111110101101001111001",
			5779 => "00000000000000000101101001111001",
			5780 => "00000000000000000101101001111001",
			5781 => "0000000100000000001000110100010000",
			5782 => "0000001100000000000100011000000100",
			5783 => "00000000000000000101101001111001",
			5784 => "0000001101000000000101110000000100",
			5785 => "00000000000000000101101001111001",
			5786 => "0000001001000000000010101100000100",
			5787 => "00000000110111000101101001111001",
			5788 => "00000000000000000101101001111001",
			5789 => "00000000000000000101101001111001",
			5790 => "0000001101000000000101110000100000",
			5791 => "0000000000000000001111001000011000",
			5792 => "0000001001000000001111000000000100",
			5793 => "00000000000000000101101100011101",
			5794 => "0000000111000000000110100100000100",
			5795 => "00000000000000000101101100011101",
			5796 => "0000001011000000000110110100001100",
			5797 => "0000001101000000000001000000000100",
			5798 => "00000000000000000101101100011101",
			5799 => "0000000101000000000001000000000100",
			5800 => "00000000111000100101101100011101",
			5801 => "00000000000000000101101100011101",
			5802 => "00000000000000000101101100011101",
			5803 => "0000000011000000001000100000000100",
			5804 => "11111111110110010101101100011101",
			5805 => "00000000000000000101101100011101",
			5806 => "0000000101000000000111100000001100",
			5807 => "0000001000000000000001010000001000",
			5808 => "0000001100000000000100011000000100",
			5809 => "00000000000000000101101100011101",
			5810 => "11111111010111100101101100011101",
			5811 => "00000000000000000101101100011101",
			5812 => "0000001101000000001010001000010100",
			5813 => "0000001100000000000100011000000100",
			5814 => "00000000000000000101101100011101",
			5815 => "0000000000000000000001010100000100",
			5816 => "00000000000000000101101100011101",
			5817 => "0000000000000000001010101100001000",
			5818 => "0000001100000000000110100100000100",
			5819 => "00000000101110110101101100011101",
			5820 => "00000000000000000101101100011101",
			5821 => "00000000000000000101101100011101",
			5822 => "0000000011000000001000100000000100",
			5823 => "00000000000000000101101100011101",
			5824 => "0000001100000000001000011000001100",
			5825 => "0000000101000000001111010000000100",
			5826 => "00000000000000000101101100011101",
			5827 => "0000000101000000000011001000000100",
			5828 => "11111111011100010101101100011101",
			5829 => "00000000000000000101101100011101",
			5830 => "00000000000000000101101100011101",
			5831 => "0000000000000000000010101000111100",
			5832 => "0000001001000000001001100100001100",
			5833 => "0000000110000000000000111100001000",
			5834 => "0000000001000000000111100100000100",
			5835 => "11111110100101000101101110101001",
			5836 => "00000001111010010101101110101001",
			5837 => "11111110011001100101101110101001",
			5838 => "0000000101000000000110100000001000",
			5839 => "0000000001000000001011111100000100",
			5840 => "00000001000110010101101110101001",
			5841 => "11111110010000010101101110101001",
			5842 => "0000000101000000000101110000011000",
			5843 => "0000000110000000000100111100010000",
			5844 => "0000001100000000001010111000001000",
			5845 => "0000000000000000000110001000000100",
			5846 => "00000001000010010101101110101001",
			5847 => "11111101111111110101101110101001",
			5848 => "0000001010000000000000001000000100",
			5849 => "11111111100001110101101110101001",
			5850 => "00000001100011110101101110101001",
			5851 => "0000000101000000001001010000000100",
			5852 => "00000011110001100101101110101001",
			5853 => "00000010011010000101101110101001",
			5854 => "0000000100000000001101101100000100",
			5855 => "00000001111100010101101110101001",
			5856 => "0000000111000000000101110100001000",
			5857 => "0000000111000000000000011100000100",
			5858 => "11111101010100000101101110101001",
			5859 => "11111110101110000101101110101001",
			5860 => "00000001000100010101101110101001",
			5861 => "0000000000000000001010101100001000",
			5862 => "0000000110000000001000010000000100",
			5863 => "11111110011011000101101110101001",
			5864 => "00000001100001110101101110101001",
			5865 => "11111110011000110101101110101001",
			5866 => "0000000100000000001000001100100100",
			5867 => "0000001100000000001010111000000100",
			5868 => "00000000000000000101110001011101",
			5869 => "0000000111000000001000011000010000",
			5870 => "0000000001000000001011111100001100",
			5871 => "0000000001000000001001011000000100",
			5872 => "00000000000000000101110001011101",
			5873 => "0000001001000000001111000000000100",
			5874 => "00000000000000000101110001011101",
			5875 => "00000000111111010101110001011101",
			5876 => "00000000000000000101110001011101",
			5877 => "0000000000000000000001010100001000",
			5878 => "0000000000000000000101000100000100",
			5879 => "00000000000000000101110001011101",
			5880 => "11111111101100010101110001011101",
			5881 => "0000000000000000000001010100000100",
			5882 => "00000000000000000101110001011101",
			5883 => "00000000010011010101110001011101",
			5884 => "0000000011000000001010000100010000",
			5885 => "0000001100000000001011000000001100",
			5886 => "0000000111000000000001101000001000",
			5887 => "0000001110000000001111010100000100",
			5888 => "11111110110110100101110001011101",
			5889 => "00000000000000000101110001011101",
			5890 => "00000000000000000101110001011101",
			5891 => "00000000000000000101110001011101",
			5892 => "0000000010000000001000001100001000",
			5893 => "0000000001000000000000111100000100",
			5894 => "00000000000000000101110001011101",
			5895 => "00000000111011010101110001011101",
			5896 => "0000001110000000000111010100001100",
			5897 => "0000001100000000001011000000001000",
			5898 => "0000000111000000000110100100000100",
			5899 => "00000000000000000101110001011101",
			5900 => "11111111000001000101110001011101",
			5901 => "00000000000000000101110001011101",
			5902 => "0000000010000000001011111000000100",
			5903 => "00000000101000110101110001011101",
			5904 => "0000001011000000000101110100001000",
			5905 => "0000000111000000001000011000000100",
			5906 => "11111111110010110101110001011101",
			5907 => "00000000011110010101110001011101",
			5908 => "0000001100000000001000011000000100",
			5909 => "11111111010000100101110001011101",
			5910 => "00000000000000000101110001011101",
			5911 => "0000001001000000000100101100111000",
			5912 => "0000000000000000001100000100101000",
			5913 => "0000000011000000001010000100011100",
			5914 => "0000001010000000000000001000010100",
			5915 => "0000000100000000001100010000001100",
			5916 => "0000000101000000001100100100001000",
			5917 => "0000001100000000000100011000000100",
			5918 => "00000000000000000101110100101001",
			5919 => "00000000010011110101110100101001",
			5920 => "00000000000000000101110100101001",
			5921 => "0000000100000000000111011000000100",
			5922 => "11111111100110010101110100101001",
			5923 => "00000000000000000101110100101001",
			5924 => "0000001001000000001111000000000100",
			5925 => "00000000000000000101110100101001",
			5926 => "00000000110011110101110100101001",
			5927 => "0000001100000000001001001000001000",
			5928 => "0000001000000000001000010100000100",
			5929 => "11111111011000100101110100101001",
			5930 => "00000000000000000101110100101001",
			5931 => "00000000000000000101110100101001",
			5932 => "0000001100000000001000011000001100",
			5933 => "0000001000000000001000010100000100",
			5934 => "00000000000000000101110100101001",
			5935 => "0000001010000000001010100000000100",
			5936 => "00000000000000000101110100101001",
			5937 => "11111111001101110101110100101001",
			5938 => "00000000000000000101110100101001",
			5939 => "0000001010000000000010101100001000",
			5940 => "0000001001000000000100101100000100",
			5941 => "00000000000000000101110100101001",
			5942 => "11111111011000000101110100101001",
			5943 => "0000000000000000000001110100011100",
			5944 => "0000000101000000001101000100010000",
			5945 => "0000000111000000000110100100001000",
			5946 => "0000000111000000001001001000000100",
			5947 => "00000000000000000101110100101001",
			5948 => "00000000010001100101110100101001",
			5949 => "0000000100000000001011101100000100",
			5950 => "00000000000000000101110100101001",
			5951 => "11111111100111010101110100101001",
			5952 => "0000000011000000000010010100001000",
			5953 => "0000001001000000000010101100000100",
			5954 => "00000000110011110101110100101001",
			5955 => "00000000000000000101110100101001",
			5956 => "00000000000000000101110100101001",
			5957 => "0000000011000000001000101000001000",
			5958 => "0000001000000000000001010100000100",
			5959 => "11111111100100000101110100101001",
			5960 => "00000000000000000101110100101001",
			5961 => "00000000000000000101110100101001",
			5962 => "0000000000000000000010101001000100",
			5963 => "0000000001000000001001011000010100",
			5964 => "0000001010000000001001100100001100",
			5965 => "0000000010000000000001101000000100",
			5966 => "11111111001000110101110111011101",
			5967 => "0000001001000000001110010100000100",
			5968 => "00000001000001000101110111011101",
			5969 => "00000000000000000101110111011101",
			5970 => "0000001001000000001111000000000100",
			5971 => "11111110011100110101110111011101",
			5972 => "00000000000000000101110111011101",
			5973 => "0000000000000000001111001000011000",
			5974 => "0000001000000000001100011100010000",
			5975 => "0000000001000000001101111100001100",
			5976 => "0000000011000000001000100000001000",
			5977 => "0000001101000000000101110000000100",
			5978 => "00000001010000000101110111011101",
			5979 => "00000000100110110101110111011101",
			5980 => "11111111010001010101110111011101",
			5981 => "11111100001010100101110111011101",
			5982 => "0000000011000000001000001100000100",
			5983 => "00000000000000000101110111011101",
			5984 => "00000001111111010101110111011101",
			5985 => "0000000011000000001111100100000100",
			5986 => "11111101110110010101110111011101",
			5987 => "0000001101000000001010001000001000",
			5988 => "0000001011000000001011011100000100",
			5989 => "00000000000000000101110111011101",
			5990 => "00000001100010010101110111011101",
			5991 => "0000001010000000001000010100001000",
			5992 => "0000000100000000000010010100000100",
			5993 => "00000000001111010101110111011101",
			5994 => "11111110101011010101110111011101",
			5995 => "00000001000100000101110111011101",
			5996 => "0000000000000000001010101100010100",
			5997 => "0000000000000000001010101100000100",
			5998 => "11111110111111110101110111011101",
			5999 => "0000000001000000001010011000001100",
			6000 => "0000001001000000000010101100000100",
			6001 => "11111111101111110101110111011101",
			6002 => "0000000001000000001100011000000100",
			6003 => "00000000110111000101110111011101",
			6004 => "00000000000000000101110111011101",
			6005 => "11111111100010000101110111011101",
			6006 => "11111110011001110101110111011101",
			6007 => "0000000000000000000001110101000000",
			6008 => "0000001001000000001111000000010100",
			6009 => "0000000001000000001001011000010000",
			6010 => "0000000110000000000000111100001000",
			6011 => "0000000001000000000111100100000100",
			6012 => "11111110011101100101111010100001",
			6013 => "00001001011111100101111010100001",
			6014 => "0000001011000000000010001000000100",
			6015 => "11111110011000100101111010100001",
			6016 => "11111111101110000101111010100001",
			6017 => "00000001110011000101111010100001",
			6018 => "0000000101000000000110100000001100",
			6019 => "0000000011000000000111010100001000",
			6020 => "0000000001000000001011111100000100",
			6021 => "00000001111101100101111010100001",
			6022 => "11111110010110000101111010100001",
			6023 => "00000100110100110101111010100001",
			6024 => "0000000011000000000010010100011100",
			6025 => "0000000001000000001001011000001100",
			6026 => "0000001010000000000000001000001000",
			6027 => "0000000101000000001100100100000100",
			6028 => "00000100111100000101111010100001",
			6029 => "11111110010011000101111010100001",
			6030 => "00000010010011100101111010100001",
			6031 => "0000000000000000001111001000001000",
			6032 => "0000001001000000001111000000000100",
			6033 => "00000101000100100101111010100001",
			6034 => "00000010100111010101111010100001",
			6035 => "0000000011000000001111100100000100",
			6036 => "11111101110000110101111010100001",
			6037 => "00000010101111110101111010100001",
			6038 => "11111110100010000101111010100001",
			6039 => "0000000000000000000010101000010000",
			6040 => "0000001000000000000001010100001100",
			6041 => "0000000100000000001011110000001000",
			6042 => "0000001000000000000101000100000100",
			6043 => "11111110011110110101111010100001",
			6044 => "00000001001110010101111010100001",
			6045 => "11111110011001000101111010100001",
			6046 => "00000110110111000101111010100001",
			6047 => "0000000000000000001010101100010000",
			6048 => "0000001000000000000001110000001100",
			6049 => "0000000110000000001000010000000100",
			6050 => "11111110011000010101111010100001",
			6051 => "0000001000000000000001010100000100",
			6052 => "11111110111001100101111010100001",
			6053 => "00000000010101010101111010100001",
			6054 => "00000100011100100101111010100001",
			6055 => "11111110010111100101111010100001",
			6056 => "0000001001000000001001111100110100",
			6057 => "0000000000000000001100000100101100",
			6058 => "0000001010000000001010100000011100",
			6059 => "0000001101000000000101110000010000",
			6060 => "0000001011000000000110110100001100",
			6061 => "0000000001000000001101101000000100",
			6062 => "00000000000000000101111101100101",
			6063 => "0000000011000000001100000000000100",
			6064 => "00000000010010000101111101100101",
			6065 => "00000000000000000101111101100101",
			6066 => "00000000000000000101111101100101",
			6067 => "0000001101000000000111111100001000",
			6068 => "0000001001000000001111000000000100",
			6069 => "00000000000000000101111101100101",
			6070 => "11111111010011010101111101100101",
			6071 => "00000000000000000101111101100101",
			6072 => "0000000011000000001000001100001100",
			6073 => "0000000111000000000110100100000100",
			6074 => "00000000000000000101111101100101",
			6075 => "0000001111000000001001100000000100",
			6076 => "00000000000000000101111101100101",
			6077 => "00000000110010010101111101100101",
			6078 => "00000000000000000101111101100101",
			6079 => "0000001100000000001000011000000100",
			6080 => "11111111010110000101111101100101",
			6081 => "00000000000000000101111101100101",
			6082 => "0000000000000000000111000100011000",
			6083 => "0000000011000000000110111100000100",
			6084 => "00000000000000000101111101100101",
			6085 => "0000001100000000000100011000001100",
			6086 => "0000001100000000001010111000001000",
			6087 => "0000001100000000000111001000000100",
			6088 => "00000000000000000101111101100101",
			6089 => "00000000000110000101111101100101",
			6090 => "00000000000000000101111101100101",
			6091 => "0000001101000000001110000100000100",
			6092 => "00000000000000000101111101100101",
			6093 => "00000001000100010101111101100101",
			6094 => "0000000011000000001100111000000100",
			6095 => "11111111101010110101111101100101",
			6096 => "0000000100000000001000110100010000",
			6097 => "0000000110000000000100111100000100",
			6098 => "00000000000000000101111101100101",
			6099 => "0000000100000000001011110000000100",
			6100 => "00000000000000000101111101100101",
			6101 => "0000000011000000000110111000000100",
			6102 => "00000000101001110101111101100101",
			6103 => "00000000000000000101111101100101",
			6104 => "00000000000000000101111101100101",
			6105 => "0000000000000000000010101001000000",
			6106 => "0000000011000000001100111000110000",
			6107 => "0000000000000000000111000100101000",
			6108 => "0000001001000000000111101100100000",
			6109 => "0000001111000000001111010100010000",
			6110 => "0000000001000000001001011000001000",
			6111 => "0000000110000000000100110100000100",
			6112 => "11111111011001000101111111110001",
			6113 => "00000000000000000101111111110001",
			6114 => "0000001011000000000100010000000100",
			6115 => "00000000100110100101111111110001",
			6116 => "11111111111001110101111111110001",
			6117 => "0000001100000000001011000000001000",
			6118 => "0000001001000000000100101100000100",
			6119 => "11111110110011110101111111110001",
			6120 => "11111111111001000101111111110001",
			6121 => "0000000001000000000001000100000100",
			6122 => "11111111101010100101111111110001",
			6123 => "00000000111111010101111111110001",
			6124 => "0000000011000000001010000100000100",
			6125 => "00000000000000000101111111110001",
			6126 => "00000001010100000101111111110001",
			6127 => "0000001100000000000100011000000100",
			6128 => "00000000000000000101111111110001",
			6129 => "11111110101010110101111111110001",
			6130 => "0000000010000000001101101100000100",
			6131 => "00000001010001100101111111110001",
			6132 => "0000001101000000001110010000000100",
			6133 => "00000000010100100101111111110001",
			6134 => "0000000010000000000011000000000100",
			6135 => "11111111101100010101111111110001",
			6136 => "00000000000000000101111111110001",
			6137 => "0000001001000000000010101100000100",
			6138 => "11111110100010010101111111110001",
			6139 => "00000000000000000101111111110001",
			6140 => "0000000000000000000001110101000000",
			6141 => "0000001001000000001111000000010000",
			6142 => "0000001011000000000010001000001100",
			6143 => "0000000110000000000000111100001000",
			6144 => "0000000001000000000111100100000100",
			6145 => "11111110100001110110000010100101",
			6146 => "00000010010011010110000010100101",
			6147 => "11111110011001010110000010100101",
			6148 => "00000000000000000110000010100101",
			6149 => "0000001011000000000100000100001000",
			6150 => "0000000010000000001001100000000100",
			6151 => "00000000001010000110000010100101",
			6152 => "11111110011101000110000010100101",
			6153 => "0000001101000000001100010100100000",
			6154 => "0000000001000000000000111100010000",
			6155 => "0000000111000000001000011000001000",
			6156 => "0000000101000000000111100000000100",
			6157 => "00000001001000110110000010100101",
			6158 => "11111110101110110110000010100101",
			6159 => "0000001011000000000100010000000100",
			6160 => "00000001010000010110000010100101",
			6161 => "00000011000111100110000010100101",
			6162 => "0000000000000000001111001000001000",
			6163 => "0000001101000000000111100000000100",
			6164 => "11111111001100100110000010100101",
			6165 => "00000001110110010110000010100101",
			6166 => "0000000011000000001111100100000100",
			6167 => "11111101110000100110000010100101",
			6168 => "00000010001001000110000010100101",
			6169 => "0000000000000000001111001000000100",
			6170 => "00000000001010110110000010100101",
			6171 => "11111110011101000110000010100101",
			6172 => "0000000000000000001010101100011000",
			6173 => "0000001000000000000001010100010000",
			6174 => "0000000000000000000001110100001100",
			6175 => "0000000001000000000100110100001000",
			6176 => "0000000011000000000110010000000100",
			6177 => "00000000000000000110000010100101",
			6178 => "00000011101010010110000010100101",
			6179 => "11111110101001100110000010100101",
			6180 => "11111110011001110110000010100101",
			6181 => "0000000110000000001000010000000100",
			6182 => "00000000000101000110000010100101",
			6183 => "00000010111111010110000010100101",
			6184 => "11111110011000100110000010100101",
			6185 => "0000000100000000001111100101000000",
			6186 => "0000001010000000001010100000100000",
			6187 => "0000001101000000000101110000001000",
			6188 => "0000001001000000001111000000000100",
			6189 => "00000000000000000110000110011001",
			6190 => "00000000011111110110000110011001",
			6191 => "0000000010000000000010000100001100",
			6192 => "0000001000000000001000100100001000",
			6193 => "0000001100000000000100011000000100",
			6194 => "00000000000000000110000110011001",
			6195 => "11111110110110100110000110011001",
			6196 => "00000000000000000110000110011001",
			6197 => "0000000011000000000111010100001000",
			6198 => "0000001100000000001000000000000100",
			6199 => "00000000000000000110000110011001",
			6200 => "00000000110001100110000110011001",
			6201 => "11111111101001000110000110011001",
			6202 => "0000000011000000001011111000011000",
			6203 => "0000001101000000001110000100001000",
			6204 => "0000000000000000001100000100000100",
			6205 => "00000000000000000110000110011001",
			6206 => "11111111101110000110000110011001",
			6207 => "0000000001000000000000111100000100",
			6208 => "00000000000000000110000110011001",
			6209 => "0000000001000000000111101000001000",
			6210 => "0000000011000000001100000000000100",
			6211 => "00000000000000000110000110011001",
			6212 => "00000001010110010110000110011001",
			6213 => "00000000000000000110000110011001",
			6214 => "0000001011000000001011110100000100",
			6215 => "11111111101001010110000110011001",
			6216 => "00000000000000000110000110011001",
			6217 => "0000000001000000000111101000010100",
			6218 => "0000001100000000001001110100001100",
			6219 => "0000001000000000000110011000000100",
			6220 => "00000000000000000110000110011001",
			6221 => "0000001001000000000100101100000100",
			6222 => "11111110100001010110000110011001",
			6223 => "00000000000000000110000110011001",
			6224 => "0000001000000000001100011100000100",
			6225 => "00000000100110110110000110011001",
			6226 => "00000000000000000110000110011001",
			6227 => "0000000000000000000110001000001000",
			6228 => "0000000011000000001000001100000100",
			6229 => "11111111101010100110000110011001",
			6230 => "00000001001000100110000110011001",
			6231 => "0000000011000000001111100100001000",
			6232 => "0000001011000000000000011100000100",
			6233 => "00000000000000000110000110011001",
			6234 => "11111110110011110110000110011001",
			6235 => "0000000000000000000111000100001000",
			6236 => "0000000001000000001100011000000100",
			6237 => "00000000110111010110000110011001",
			6238 => "00000000000000000110000110011001",
			6239 => "0000001110000000001100111000001000",
			6240 => "0000000000000000000001110100000100",
			6241 => "00000000000000000110000110011001",
			6242 => "11111110111110000110000110011001",
			6243 => "0000000110000000001000010000000100",
			6244 => "00000000000000000110000110011001",
			6245 => "00000000100110110110000110011001",
			6246 => "0000000100000000001011101101000000",
			6247 => "0000001010000000000010101100111000",
			6248 => "0000000001000000001110010100110000",
			6249 => "0000000111000000000001101000011100",
			6250 => "0000000100000000001100010000001100",
			6251 => "0000000011000000001100010000001000",
			6252 => "0000001100000000001101010100000100",
			6253 => "00000000000000000110001001011101",
			6254 => "00000000001100110110001001011101",
			6255 => "00000000000000000110001001011101",
			6256 => "0000000110000000001010011000001000",
			6257 => "0000001011000000000101100100000100",
			6258 => "00000000000000000110001001011101",
			6259 => "11111111010010100110001001011101",
			6260 => "0000000010000000000010000100000100",
			6261 => "00000000000000000110001001011101",
			6262 => "00000000000010110110001001011101",
			6263 => "0000000111000000001000011000001000",
			6264 => "0000000001000000001001011000000100",
			6265 => "00000000000000000110001001011101",
			6266 => "00000000101000010110001001011101",
			6267 => "0000000001000000000000111100001000",
			6268 => "0000000001000000001001011000000100",
			6269 => "00000000000000000110001001011101",
			6270 => "11111111110110010110001001011101",
			6271 => "00000000001010000110001001011101",
			6272 => "0000001100000000000100011000000100",
			6273 => "00000000000000000110001001011101",
			6274 => "11111111010011110110001001011101",
			6275 => "0000000011000000000110111100000100",
			6276 => "00000000000000000110001001011101",
			6277 => "00000000110110100110001001011101",
			6278 => "0000000110000000001111000000001100",
			6279 => "0000000000000000001011010100000100",
			6280 => "00000000000000000110001001011101",
			6281 => "0000001100000000001000011000000100",
			6282 => "11111111000010010110001001011101",
			6283 => "00000000000000000110001001011101",
			6284 => "0000000000000000000001110100010000",
			6285 => "0000000111000000000110100100000100",
			6286 => "00000000000000000110001001011101",
			6287 => "0000001011000000001011110100001000",
			6288 => "0000000011000000001011111000000100",
			6289 => "00000000000000000110001001011101",
			6290 => "00000000110100110110001001011101",
			6291 => "00000000000000000110001001011101",
			6292 => "0000000110000000001000010000000100",
			6293 => "11111111101010110110001001011101",
			6294 => "00000000000000000110001001011101",
			6295 => "0000000100000000001111100101000100",
			6296 => "0000001010000000001010100000100100",
			6297 => "0000001101000000000101110000001000",
			6298 => "0000001001000000001111000000000100",
			6299 => "00000000000000000110001101000001",
			6300 => "00000000100000100110001101000001",
			6301 => "0000000010000000000010000100001100",
			6302 => "0000001000000000001000100100001000",
			6303 => "0000001100000000000100011000000100",
			6304 => "00000000000000000110001101000001",
			6305 => "11111110101111100110001101000001",
			6306 => "00000000000000000110001101000001",
			6307 => "0000000011000000001010000100001000",
			6308 => "0000001100000000001000000000000100",
			6309 => "00000000000000000110001101000001",
			6310 => "00000000110001110110001101000001",
			6311 => "0000001011000000000100010000000100",
			6312 => "11111111011101110110001101000001",
			6313 => "00000000000000000110001101000001",
			6314 => "0000000011000000001011111000011000",
			6315 => "0000001101000000001111010000010000",
			6316 => "0000001100000000000100011000001000",
			6317 => "0000001010000000001010100000000100",
			6318 => "00000000000000000110001101000001",
			6319 => "11111111100101100110001101000001",
			6320 => "0000001100000000000100011000000100",
			6321 => "00000000010100000110001101000001",
			6322 => "00000000000000000110001101000001",
			6323 => "0000000001000000000000111100000100",
			6324 => "00000000000000000110001101000001",
			6325 => "00000001011001010110001101000001",
			6326 => "0000001011000000001011110100000100",
			6327 => "11111111100000100110001101000001",
			6328 => "00000000000000000110001101000001",
			6329 => "0000001110000000000111010100001000",
			6330 => "0000001011000000000110110100000100",
			6331 => "11111110101110010110001101000001",
			6332 => "00000000000000000110001101000001",
			6333 => "0000000100000000001101101100000100",
			6334 => "00000001000111100110001101000001",
			6335 => "0000000001000000001110010100001000",
			6336 => "0000001100000000001000011000000100",
			6337 => "11111110100101010110001101000001",
			6338 => "00000000000000000110001101000001",
			6339 => "0000000011000000001000101000010000",
			6340 => "0000000000000000000111000100001000",
			6341 => "0000000010000000001111100100000100",
			6342 => "00000000000000000110001101000001",
			6343 => "00000000110100100110001101000001",
			6344 => "0000001110000000001100111000000100",
			6345 => "11111110110111100110001101000001",
			6346 => "00000000000000000110001101000001",
			6347 => "0000001111000000001110000000001000",
			6348 => "0000000000000000001010101100000100",
			6349 => "00000001000011000110001101000001",
			6350 => "00000000000000000110001101000001",
			6351 => "00000000000000000110001101000001",
			6352 => "0000001001000000000111101101010000",
			6353 => "0000000000000000001001101000111100",
			6354 => "0000001101000000000010011100010000",
			6355 => "0000001101000000000101001000001000",
			6356 => "0000001001000000000101010000000100",
			6357 => "00000000000000000110010000111101",
			6358 => "11111111111101010110010000111101",
			6359 => "0000001001000000001111000000000100",
			6360 => "00000000000000000110010000111101",
			6361 => "00000001000011100110010000111101",
			6362 => "0000001011000000000110110100010000",
			6363 => "0000001011000000000101100100000100",
			6364 => "00000000000000000110010000111101",
			6365 => "0000001010000000000010101100001000",
			6366 => "0000000010000000000110010000000100",
			6367 => "00000000000000000110010000111101",
			6368 => "11111110111011110110010000111101",
			6369 => "00000000000000000110010000111101",
			6370 => "0000000110000000000100110100010000",
			6371 => "0000000001000000001001011000001000",
			6372 => "0000001011000000000010001000000100",
			6373 => "00000000000000000110010000111101",
			6374 => "00000000010111110110010000111101",
			6375 => "0000001100000000001001110100000100",
			6376 => "11111111001111100110010000111101",
			6377 => "00000000000000000110010000111101",
			6378 => "0000000011000000001011111000001000",
			6379 => "0000001001000000001111000000000100",
			6380 => "00000000000000000110010000111101",
			6381 => "00000000111010000110010000111101",
			6382 => "00000000000000000110010000111101",
			6383 => "0000001100000000000001101000001000",
			6384 => "0000000001000000000001111000000100",
			6385 => "11111111000010000110010000111101",
			6386 => "00000000000000000110010000111101",
			6387 => "0000000001000000000001000100000100",
			6388 => "00000000000000000110010000111101",
			6389 => "0000000001000000000111101000000100",
			6390 => "00000000000110110110010000111101",
			6391 => "00000000000000000110010000111101",
			6392 => "0000000000000000000111000100010000",
			6393 => "0000000110000000001011001100000100",
			6394 => "00000000000000000110010000111101",
			6395 => "0000000011000000000111010100000100",
			6396 => "00000000000000000110010000111101",
			6397 => "0000001011000000000101110100000100",
			6398 => "00000001000101000110010000111101",
			6399 => "00000000000000000110010000111101",
			6400 => "0000001110000000001100111000001100",
			6401 => "0000001100000000000100011000000100",
			6402 => "00000000000000000110010000111101",
			6403 => "0000000011000000000011000000000100",
			6404 => "11111111011010100110010000111101",
			6405 => "00000000000000000110010000111101",
			6406 => "0000001111000000001110000000010000",
			6407 => "0000000110000000001000010000000100",
			6408 => "00000000000000000110010000111101",
			6409 => "0000001100000000000100011000000100",
			6410 => "00000000000000000110010000111101",
			6411 => "0000000011000000001101101100000100",
			6412 => "00000000000000000110010000111101",
			6413 => "00000000111000000110010000111101",
			6414 => "00000000000000000110010000111101",
			6415 => "0000000111000000000110100100010100",
			6416 => "0000000100000000000111010100001100",
			6417 => "0000000001000000001011111100001000",
			6418 => "0000000001000000001101101000000100",
			6419 => "00000000000000000110010100100001",
			6420 => "00000000001111010110010100100001",
			6421 => "00000000000000000110010100100001",
			6422 => "0000000110000000001011001100000100",
			6423 => "11111110100011000110010100100001",
			6424 => "00000000000000000110010100100001",
			6425 => "0000000111000000000001101000101000",
			6426 => "0000000110000000001011001100011100",
			6427 => "0000000100000000001011101100011000",
			6428 => "0000001010000000001010100000001100",
			6429 => "0000000110000000001101111100000100",
			6430 => "00000000000000000110010100100001",
			6431 => "0000001111000000001001100000000100",
			6432 => "00000000000000000110010100100001",
			6433 => "11111111101001010110010100100001",
			6434 => "0000001001000000000100111100000100",
			6435 => "00000000000000000110010100100001",
			6436 => "0000000011000000000110111100000100",
			6437 => "00000000000000000110010100100001",
			6438 => "00000000111000010110010100100001",
			6439 => "11111111011101010110010100100001",
			6440 => "0000000000000000000001110100001000",
			6441 => "0000000011000000001000001100000100",
			6442 => "00000000000000000110010100100001",
			6443 => "00000001010000000110010100100001",
			6444 => "11111111111110110110010100100001",
			6445 => "0000001011000000001011011100010000",
			6446 => "0000001011000000000101100100000100",
			6447 => "00000000000000000110010100100001",
			6448 => "0000000011000000000000010000001000",
			6449 => "0000001111000000001001100000000100",
			6450 => "00000000000000000110010100100001",
			6451 => "11111110110000010110010100100001",
			6452 => "00000000000000000110010100100001",
			6453 => "0000000100000000001101101100010100",
			6454 => "0000000001000000000000111100010000",
			6455 => "0000000011000000001010000100001000",
			6456 => "0000001100000000001001110100000100",
			6457 => "00000000100110100110010100100001",
			6458 => "00000000000000000110010100100001",
			6459 => "0000000111000000001111011100000100",
			6460 => "11111111100010000110010100100001",
			6461 => "00000000000000000110010100100001",
			6462 => "00000001000101000110010100100001",
			6463 => "0000000011000000001101101100001000",
			6464 => "0000000101000000000111100000000100",
			6465 => "00000000000000000110010100100001",
			6466 => "11111111000110000110010100100001",
			6467 => "0000000101000000000111111100001000",
			6468 => "0000000000000000000111000000000100",
			6469 => "00000000101001100110010100100001",
			6470 => "00000000000000000110010100100001",
			6471 => "00000000000000000110010100100001",
			6472 => "0000000000000000001010101101000000",
			6473 => "0000001100000000000111001000001100",
			6474 => "0000000111000000000110100100000100",
			6475 => "11111110010100000110010110100101",
			6476 => "0000000110000000001101111100000100",
			6477 => "00000000000000000110010110100101",
			6478 => "00000000001110000110010110100101",
			6479 => "0000001010000000001000010100110000",
			6480 => "0000001101000000000011001000011100",
			6481 => "0000000000000000001111001000001100",
			6482 => "0000001110000000000111010100001000",
			6483 => "0000000100000000001011101100000100",
			6484 => "00000000110011100110010110100101",
			6485 => "11111110101010000110010110100101",
			6486 => "00000001111001100110010110100101",
			6487 => "0000001101000000000101110000001000",
			6488 => "0000001111000000001011101100000100",
			6489 => "11111101110000010110010110100101",
			6490 => "11111111011100000110010110100101",
			6491 => "0000001110000000001100111000000100",
			6492 => "00000000101000010110010110100101",
			6493 => "00000001111110100110010110100101",
			6494 => "0000000100000000001101101100001000",
			6495 => "0000000111000000001111011100000100",
			6496 => "00000000000000000110010110100101",
			6497 => "00000001100000100110010110100101",
			6498 => "0000000111000000000101110100001000",
			6499 => "0000001000000000000001010100000100",
			6500 => "11111110001010000110010110100101",
			6501 => "00000000000000000110010110100101",
			6502 => "00000000100111000110010110100101",
			6503 => "00000100001110110110010110100101",
			6504 => "11111110011010000110010110100101",
			6505 => "0000001100000000000100011000101100",
			6506 => "0000000000000000001011010100011100",
			6507 => "0000001111000000000110111100011000",
			6508 => "0000001100000000001010111000001000",
			6509 => "0000000111000000000110100100000100",
			6510 => "11111111011001110110011010111001",
			6511 => "00000000000000000110011010111001",
			6512 => "0000000100000000000111010100001100",
			6513 => "0000000011000000000110111100001000",
			6514 => "0000000111000000001011000000000100",
			6515 => "00000000000000000110011010111001",
			6516 => "00000000010001000110011010111001",
			6517 => "00000000000000000110011010111001",
			6518 => "00000000000000000110011010111001",
			6519 => "00000000110111010110011010111001",
			6520 => "0000000111000000001000011000001100",
			6521 => "0000000100000000001011101100000100",
			6522 => "00000000000000000110011010111001",
			6523 => "0000001011000000000110110100000100",
			6524 => "11111110011101100110011010111001",
			6525 => "00000000000000000110011010111001",
			6526 => "00000000000000000110011010111001",
			6527 => "0000001100000000001011000000111100",
			6528 => "0000001101000000000100101000101100",
			6529 => "0000000100000000001000101000011100",
			6530 => "0000000110000000000100110100010000",
			6531 => "0000000100000000001100010000001000",
			6532 => "0000000110000000001101111100000100",
			6533 => "00000000000000000110011010111001",
			6534 => "00000000100001110110011010111001",
			6535 => "0000001111000000000010000100000100",
			6536 => "00000000000000000110011010111001",
			6537 => "11111111010011100110011010111001",
			6538 => "0000000000000000001111001000001000",
			6539 => "0000000011000000001100000000000100",
			6540 => "00000000000000000110011010111001",
			6541 => "00000001010000010110011010111001",
			6542 => "00000000000000000110011010111001",
			6543 => "0000000011000000001000100000001000",
			6544 => "0000001011000000000001011000000100",
			6545 => "00000000000000000110011010111001",
			6546 => "11111111000011110110011010111001",
			6547 => "0000000010000000001101101100000100",
			6548 => "00000000111011010110011010111001",
			6549 => "00000000000000000110011010111001",
			6550 => "0000000010000000001100010000001000",
			6551 => "0000001011000000000010001000000100",
			6552 => "11111111110011110110011010111001",
			6553 => "00000000100111010110011010111001",
			6554 => "0000000110000000001011001100000100",
			6555 => "11111110111100100110011010111001",
			6556 => "00000000000000000110011010111001",
			6557 => "0000000010000000001110110100001000",
			6558 => "0000001101000000000100101000000100",
			6559 => "00000000000000000110011010111001",
			6560 => "11111111110011000110011010111001",
			6561 => "0000001100000000000110100100010000",
			6562 => "0000000000000000001010101100001100",
			6563 => "0000000101000000001101000100000100",
			6564 => "00000000000000000110011010111001",
			6565 => "0000001101000000001100010100000100",
			6566 => "00000001001010110110011010111001",
			6567 => "00000000000000000110011010111001",
			6568 => "00000000000000000110011010111001",
			6569 => "0000001000000000001100011100001000",
			6570 => "0000001011000000000101110100000100",
			6571 => "00000000000000000110011010111001",
			6572 => "00000000101100010110011010111001",
			6573 => "11111111101111110110011010111001",
			6574 => "0000001001000000001111000000010000",
			6575 => "0000001010000000001001100100001100",
			6576 => "0000000010000000000001101000000100",
			6577 => "11111110101111000110011110001101",
			6578 => "0000000110000000000101011100000100",
			6579 => "00000001111101010110011110001101",
			6580 => "00000000000000000110011110001101",
			6581 => "11111110011000110110011110001101",
			6582 => "0000001101000000001100010101000100",
			6583 => "0000000111000000000110100100100100",
			6584 => "0000000010000000001100000000001100",
			6585 => "0000000101000000000010110100000100",
			6586 => "11111111000101010110011110001101",
			6587 => "0000000101000000001100100100000100",
			6588 => "00000001100101100110011110001101",
			6589 => "00000000010010010110011110001101",
			6590 => "0000001100000000000100011000001100",
			6591 => "0000001010000000000010101100000100",
			6592 => "11111100011000010110011110001101",
			6593 => "0000001010000000000011101000000100",
			6594 => "00000000110000110110011110001101",
			6595 => "11111110000100000110011110001101",
			6596 => "0000001101000000001111010000000100",
			6597 => "11111110011000010110011110001101",
			6598 => "0000000100000000000110111000000100",
			6599 => "00000001011101110110011110001101",
			6600 => "00000000000000000110011110001101",
			6601 => "0000001010000000001001000100011100",
			6602 => "0000001110000000001100111000010000",
			6603 => "0000001000000000001000100100001000",
			6604 => "0000000100000000001100010000000100",
			6605 => "00000001101001010110011110001101",
			6606 => "11111110101110110110011110001101",
			6607 => "0000000001000000001101111100000100",
			6608 => "00000001001110000110011110001101",
			6609 => "11111111110111010110011110001101",
			6610 => "0000001110000000000011000000001000",
			6611 => "0000000100000000001000110100000100",
			6612 => "00000010011010110110011110001101",
			6613 => "00000000000000000110011110001101",
			6614 => "00000101110101100110011110001101",
			6615 => "11111110100010110110011110001101",
			6616 => "0000001001000000000100101100010100",
			6617 => "0000001100000000001001110100000100",
			6618 => "11111111010010100110011110001101",
			6619 => "0000000111000000000101100100001000",
			6620 => "0000001011000000000001001000000100",
			6621 => "00000001110100010110011110001101",
			6622 => "00000000000000000110011110001101",
			6623 => "0000001100000000000100000100000100",
			6624 => "11111111100010110110011110001101",
			6625 => "00000000000000000110011110001101",
			6626 => "11111110011100100110011110001101",
			6627 => "0000001100000000001010111000010000",
			6628 => "0000000000000000000110001000001100",
			6629 => "0000001110000000001100000000001000",
			6630 => "0000000111000000000110100100000100",
			6631 => "11111111010000000110100010000001",
			6632 => "00000000000000000110100010000001",
			6633 => "00000000011000010110100010000001",
			6634 => "11111110011111010110100010000001",
			6635 => "0000001001000000000100101101000100",
			6636 => "0000000010000000001100010000100100",
			6637 => "0000001101000000000101001000001000",
			6638 => "0000000000000000000001010100000100",
			6639 => "00000000000000000110100010000001",
			6640 => "11111111010000000110100010000001",
			6641 => "0000000000000000000101000100010000",
			6642 => "0000000011000000001100000000001000",
			6643 => "0000001010000000000111101100000100",
			6644 => "00000000000000000110100010000001",
			6645 => "00000000110100000110100010000001",
			6646 => "0000000001000000000000111100000100",
			6647 => "11111111000111110110100010000001",
			6648 => "00000000000000000110100010000001",
			6649 => "0000001010000000000000001000000100",
			6650 => "00000000000000000110100010000001",
			6651 => "0000000011000000001010000100000100",
			6652 => "00000001010100100110100010000001",
			6653 => "00000000000000000110100010000001",
			6654 => "0000001100000000001001110100010000",
			6655 => "0000001100000000000100011000000100",
			6656 => "00000000000000000110100010000001",
			6657 => "0000001011000000000101100100000100",
			6658 => "00000000000000000110100010000001",
			6659 => "0000001101000000000010011100000100",
			6660 => "00000000000000000110100010000001",
			6661 => "11111111001000100110100010000001",
			6662 => "0000001010000000001010100100000100",
			6663 => "00000001000001010110100010000001",
			6664 => "0000000001000000000000111100000100",
			6665 => "11111111001100110110100010000001",
			6666 => "0000000010000000001101101100000100",
			6667 => "00000000110011100110100010000001",
			6668 => "00000000000000000110100010000001",
			6669 => "0000000100000000000001011100001100",
			6670 => "0000000011000000000110111100000100",
			6671 => "11111111101111100110100010000001",
			6672 => "0000000001000000001101111100000100",
			6673 => "00000001010110000110100010000001",
			6674 => "00000000000000000110100010000001",
			6675 => "0000000010000000001000100000001000",
			6676 => "0000001011000000000101100100000100",
			6677 => "00000000000000000110100010000001",
			6678 => "11111110101111000110100010000001",
			6679 => "0000000000000000000001110100001000",
			6680 => "0000000001000000001100011000000100",
			6681 => "00000001001011110110100010000001",
			6682 => "00000000000000000110100010000001",
			6683 => "0000001110000000001100111000000100",
			6684 => "11111111000011010110100010000001",
			6685 => "0000001111000000001011110000000100",
			6686 => "00000000111100100110100010000001",
			6687 => "00000000000000000110100010000001",
			6688 => "0000001001000000001001100100001100",
			6689 => "0000001010000000001001100100001000",
			6690 => "0000000100000000000111010000000100",
			6691 => "00000000000000000110100101001101",
			6692 => "00000000001000010110100101001101",
			6693 => "11111110011011000110100101001101",
			6694 => "0000000100000000001100010000001100",
			6695 => "0000000011000000001100000000001000",
			6696 => "0000001001000000001111000000000100",
			6697 => "00000000000000000110100101001101",
			6698 => "00000001110000010110100101001101",
			6699 => "11111111101000000110100101001101",
			6700 => "0000000111000000000110100100101000",
			6701 => "0000000011000000001010000100011100",
			6702 => "0000000100000000000111010100010000",
			6703 => "0000000001000000001011111100001000",
			6704 => "0000001001000000001000010000000100",
			6705 => "00000000000000000110100101001101",
			6706 => "00000000100111010110100101001101",
			6707 => "0000000111000000001001001000000100",
			6708 => "00000000000000000110100101001101",
			6709 => "11111111011001100110100101001101",
			6710 => "0000000111000000001001001000001000",
			6711 => "0000000111000000001001001000000100",
			6712 => "11111111101111100110100101001101",
			6713 => "00000000000000000110100101001101",
			6714 => "11111101101000010110100101001101",
			6715 => "0000000100000000000011000000000100",
			6716 => "00000001000110000110100101001101",
			6717 => "0000001011000000001011011100000100",
			6718 => "11111110101010110110100101001101",
			6719 => "00000000000000000110100101001101",
			6720 => "0000001000000000001000100100001100",
			6721 => "0000001111000000001100000000001000",
			6722 => "0000001010000000000000001000000100",
			6723 => "11111110001110010110100101001101",
			6724 => "00000000000000000110100101001101",
			6725 => "00000000011111100110100101001101",
			6726 => "0000000010000000001100000000001100",
			6727 => "0000001011000000000101110100001000",
			6728 => "0000000011000000000010000100000100",
			6729 => "00000000000000000110100101001101",
			6730 => "00000001011100100110100101001101",
			6731 => "00000000000000000110100101001101",
			6732 => "0000001110000000001100000000001000",
			6733 => "0000001011000000000100010000000100",
			6734 => "11111110101001110110100101001101",
			6735 => "00000000000011000110100101001101",
			6736 => "0000000010000000001000001100000100",
			6737 => "00000000111111110110100101001101",
			6738 => "11111111111101010110100101001101",
			6739 => "0000001100000000001010111000001000",
			6740 => "0000000000000000000110001000000100",
			6741 => "00000000000000000110101000100001",
			6742 => "11111111000011000110101000100001",
			6743 => "0000001100000000001000000000110100",
			6744 => "0000001011000000000101110100101100",
			6745 => "0000000111000000000110100100011000",
			6746 => "0000000111000000001001001000001100",
			6747 => "0000000000000000001111001000001000",
			6748 => "0000000111000000001011000000000100",
			6749 => "00000000000000000110101000100001",
			6750 => "00000000101000110110101000100001",
			6751 => "00000000000000000110101000100001",
			6752 => "0000000011000000001000001100001000",
			6753 => "0000000100000000001000001100000100",
			6754 => "00000000000000000110101000100001",
			6755 => "11111111010000100110101000100001",
			6756 => "00000000000000000110101000100001",
			6757 => "0000000000000000000010101000010000",
			6758 => "0000000001000000000000111100001000",
			6759 => "0000000111000000001000011000000100",
			6760 => "00000000001011000110101000100001",
			6761 => "00000000000000000110101000100001",
			6762 => "0000001011000000000000011100000100",
			6763 => "00000000000000000110101000100001",
			6764 => "00000001000111110110101000100001",
			6765 => "00000000000000000110101000100001",
			6766 => "0000001001000000000101010000000100",
			6767 => "11111111101000110110101000100001",
			6768 => "00000000000000000110101000100001",
			6769 => "0000001011000000000100010000001100",
			6770 => "0000000110000000001000010000001000",
			6771 => "0000001100000000001001110100000100",
			6772 => "11111111001111110110101000100001",
			6773 => "00000000000000000110101000100001",
			6774 => "00000000000000000110101000100001",
			6775 => "0000001101000000001100010100010000",
			6776 => "0000000111000000001000011000000100",
			6777 => "00000000000000000110101000100001",
			6778 => "0000001100000000000001101000001000",
			6779 => "0000000000000000001000101100000100",
			6780 => "00000000110100010110101000100001",
			6781 => "00000000000000000110101000100001",
			6782 => "00000000000000000110101000100001",
			6783 => "0000000111000000000000011100001000",
			6784 => "0000001001000000000010101100000100",
			6785 => "11111111100010000110101000100001",
			6786 => "00000000000000000110101000100001",
			6787 => "0000000001000000000111101000001000",
			6788 => "0000001011000000001110101100000100",
			6789 => "00000000001111000110101000100001",
			6790 => "00000000000000000110101000100001",
			6791 => "00000000000000000110101000100001",
			6792 => "0000000000000000000010101001110000",
			6793 => "0000001100000000000100011000111100",
			6794 => "0000000000000000000110001000101000",
			6795 => "0000001001000000000100111100010000",
			6796 => "0000001100000000000100011000000100",
			6797 => "11111110011011100110101100101101",
			6798 => "0000001100000000000100011000000100",
			6799 => "00000001010010010110101100101101",
			6800 => "0000001100000000000100011000000100",
			6801 => "00000000000000000110101100101101",
			6802 => "11111110000001110110101100101101",
			6803 => "0000001101000000000101110000010000",
			6804 => "0000001101000000001110000100001000",
			6805 => "0000000000000000001100000100000100",
			6806 => "00000000110100000110101100101101",
			6807 => "11111110110011100110101100101101",
			6808 => "0000000001000000000111101000000100",
			6809 => "00000001110100010110101100101101",
			6810 => "00000000101111000110101100101101",
			6811 => "0000000100000000001000001100000100",
			6812 => "00000001001001100110101100101101",
			6813 => "11111110101111010110101100101101",
			6814 => "0000000110000000001001100100001100",
			6815 => "0000001000000000001100011100001000",
			6816 => "0000001111000000001010000100000100",
			6817 => "11111111011101100110101100101101",
			6818 => "11111011110010100110101100101101",
			6819 => "11111110011000110110101100101101",
			6820 => "0000000011000000001011111000000100",
			6821 => "11111110101110110110101100101101",
			6822 => "00000001000100100110101100101101",
			6823 => "0000000101000000000101110000100100",
			6824 => "0000000001000000001001011000001000",
			6825 => "0000001001000000001111000000000100",
			6826 => "11111110100000000110101100101101",
			6827 => "11111111111101100110101100101101",
			6828 => "0000001100000000001000000000010000",
			6829 => "0000000001000000000000111100001000",
			6830 => "0000000011000000001010000100000100",
			6831 => "00000001000001010110101100101101",
			6832 => "11111110000010010110101100101101",
			6833 => "0000000100000000001000101000000100",
			6834 => "00000001011000100110101100101101",
			6835 => "00000000000111010110101100101101",
			6836 => "0000001111000000001110110100000100",
			6837 => "11111110110111100110101100101101",
			6838 => "0000000101000000001001010000000100",
			6839 => "00000010000111110110101100101101",
			6840 => "00000000110110100110101100101101",
			6841 => "0000000100000000001101101100000100",
			6842 => "00000001010110100110101100101101",
			6843 => "0000001100000000001000011000000100",
			6844 => "11111101011100010110101100101101",
			6845 => "0000000011000000000010010100000100",
			6846 => "00000001001111000110101100101101",
			6847 => "11111110110011100110101100101101",
			6848 => "0000000000000000001010101100010100",
			6849 => "0000000000000000001010101100000100",
			6850 => "11111110111011000110101100101101",
			6851 => "0000000001000000001010011000001100",
			6852 => "0000001001000000000010101100000100",
			6853 => "11111111101011000110101100101101",
			6854 => "0000000001000000001100011000000100",
			6855 => "00000000111010100110101100101101",
			6856 => "00000000000000000110101100101101",
			6857 => "11111111011011010110101100101101",
			6858 => "11111110011001110110101100101101",
			6859 => "0000000000000000000010101001111100",
			6860 => "0000001100000000000100011000110100",
			6861 => "0000000000000000000110001000100100",
			6862 => "0000001001000000000100111100001100",
			6863 => "0000000110000000000000111100001000",
			6864 => "0000001100000000000110000100000100",
			6865 => "11111111000000100110110001001001",
			6866 => "00000000111100110110110001001001",
			6867 => "11111110011111010110110001001001",
			6868 => "0000001101000000000101110000010000",
			6869 => "0000001101000000001110000100001000",
			6870 => "0000000010000000000010000000000100",
			6871 => "00000000110111100110110001001001",
			6872 => "11111110110000010110110001001001",
			6873 => "0000001000000000001010110000000100",
			6874 => "00000001010011010110110001001001",
			6875 => "00000010010110100110110001001001",
			6876 => "0000000111000000000001101000000100",
			6877 => "11111110100010010110110001001001",
			6878 => "00000001001100010110110001001001",
			6879 => "0000001000000000001100011100001000",
			6880 => "0000001111000000000111010100000100",
			6881 => "11111111010111100110110001001001",
			6882 => "11111010110101110110110001001001",
			6883 => "0000001011000000001011011100000100",
			6884 => "11111110010011110110110001001001",
			6885 => "00000000101001110110110001001001",
			6886 => "0000000101000000001111010000100100",
			6887 => "0000000101000000001111010000011100",
			6888 => "0000001001000000001111000000001100",
			6889 => "0000000000000000000001010100001000",
			6890 => "0000001011000000000010001000000100",
			6891 => "11111110101010110110110001001001",
			6892 => "11111100010110010110110001001001",
			6893 => "00000000010110000110110001001001",
			6894 => "0000001100000000001011000000001000",
			6895 => "0000000000000000001111001000000100",
			6896 => "00000001000001110110110001001001",
			6897 => "11111110111010100110110001001001",
			6898 => "0000000110000000001101111100000100",
			6899 => "11111111101001100110110001001001",
			6900 => "00000001100101100110110001001001",
			6901 => "0000000001000000000000111100000100",
			6902 => "00000011100000100110110001001001",
			6903 => "00000001100110010110110001001001",
			6904 => "0000000111000000001000011000010000",
			6905 => "0000000001000000000000111100001000",
			6906 => "0000001000000000001000100100000100",
			6907 => "00000000010101100110110001001001",
			6908 => "11111101000100110110110001001001",
			6909 => "0000000011000000001011101100000100",
			6910 => "00000001011001010110110001001001",
			6911 => "00000000000000000110110001001001",
			6912 => "0000000010000000000110101100001000",
			6913 => "0000001011000000000100010000000100",
			6914 => "00000000010010010110110001001001",
			6915 => "00000001101010010110110001001001",
			6916 => "0000000001000000001110010100000100",
			6917 => "11111110010010010110110001001001",
			6918 => "0000000001000000000100110100000100",
			6919 => "00000001100110110110110001001001",
			6920 => "11111110111010110110110001001001",
			6921 => "0000000000000000001010101100010000",
			6922 => "0000000000000000001010101100000100",
			6923 => "11111111000100000110110001001001",
			6924 => "0000000001000000001010011000001000",
			6925 => "0000000001000000001100011000000100",
			6926 => "00000000000000000110110001001001",
			6927 => "00000000011101110110110001001001",
			6928 => "00000000000000000110110001001001",
			6929 => "11111110011001110110110001001001",
			6930 => "0000001100000000000111001000001000",
			6931 => "0000000111000000000110100100000100",
			6932 => "11111110011010110110110011110101",
			6933 => "00000000000000000110110011110101",
			6934 => "0000000100000000001000110101001100",
			6935 => "0000001011000000000110110100101100",
			6936 => "0000000001000000001101111100011100",
			6937 => "0000001101000000000101110000010000",
			6938 => "0000000011000000000111010100001000",
			6939 => "0000000001000000000111101000000100",
			6940 => "00000000101000010110110011110101",
			6941 => "11111101110011110110110011110101",
			6942 => "0000000000000000001111001000000100",
			6943 => "00000001101010110110110011110101",
			6944 => "00000000000000000110110011110101",
			6945 => "0000001000000000000001010000001000",
			6946 => "0000001100000000000100011000000100",
			6947 => "00000000000000000110110011110101",
			6948 => "11111110010111100110110011110101",
			6949 => "00000001010110000110110011110101",
			6950 => "0000000011000000001111100100000100",
			6951 => "11111101010110110110110011110101",
			6952 => "0000000000000000000111000100000100",
			6953 => "00000001001110000110110011110101",
			6954 => "0000001100000000000100011000000100",
			6955 => "00000000000000000110110011110101",
			6956 => "11111110110011100110110011110101",
			6957 => "0000000010000000001110110100001000",
			6958 => "0000001100000000001011000000000100",
			6959 => "00000000000000000110110011110101",
			6960 => "11111110100101000110110011110101",
			6961 => "0000000011000000001010000100001000",
			6962 => "0000001100000000001011000000000100",
			6963 => "00000000000000000110110011110101",
			6964 => "00000001110011100110110011110101",
			6965 => "0000000001000000000101011100001000",
			6966 => "0000001100000000001011000000000100",
			6967 => "11111110100010000110110011110101",
			6968 => "00000000010111110110110011110101",
			6969 => "0000001101000000001100010100000100",
			6970 => "00000001100011100110110011110101",
			6971 => "11111111101011000110110011110101",
			6972 => "11111110101010010110110011110101",
			6973 => "0000000000000000001010101101101100",
			6974 => "0000000111000000001000011001001000",
			6975 => "0000000111000000001000011000111000",
			6976 => "0000000111000000000110100100011000",
			6977 => "0000000111000000001001001000001100",
			6978 => "0000000111000000001011000000000100",
			6979 => "11111111000001000110110111010001",
			6980 => "0000001101000000001001010000000100",
			6981 => "00000000101101110110110111010001",
			6982 => "00000000000000000110110111010001",
			6983 => "0000000010000000000110010000000100",
			6984 => "00000000000000000110110111010001",
			6985 => "0000001011000000000000011100000100",
			6986 => "00000000000000000110110111010001",
			6987 => "11111110100011110110110111010001",
			6988 => "0000000101000000001101000100010000",
			6989 => "0000001011000000000000011100001000",
			6990 => "0000001011000000000100000100000100",
			6991 => "00000000000000000110110111010001",
			6992 => "00000001100001000110110111010001",
			6993 => "0000000001000000001011111100000100",
			6994 => "00000000001000000110110111010001",
			6995 => "11111101111100110110110111010001",
			6996 => "0000000001000000001101111100001000",
			6997 => "0000001000000000001000010100000100",
			6998 => "00000000000000000110110111010001",
			6999 => "00000000111111010110110111010001",
			7000 => "0000001011000000001011011100000100",
			7001 => "11111110100010110110110111010001",
			7002 => "00000000001111010110110111010001",
			7003 => "0000000110000000000100110100000100",
			7004 => "00000000000000000110110111010001",
			7005 => "0000001101000000000101110000000100",
			7006 => "00000000000000000110110111010001",
			7007 => "0000000110000000001011001100000100",
			7008 => "11111110011110010110110111010001",
			7009 => "00000000000000000110110111010001",
			7010 => "0000001101000000001010001000001000",
			7011 => "0000001000000000001000100100000100",
			7012 => "00000000000000000110110111010001",
			7013 => "00000001011010000110110111010001",
			7014 => "0000001011000000000101110100001000",
			7015 => "0000000101000000001001010000000100",
			7016 => "00000000000010010110110111010001",
			7017 => "11111110001110000110110111010001",
			7018 => "0000001101000000001100010100001000",
			7019 => "0000001101000000001110010000000100",
			7020 => "00000000000000000110110111010001",
			7021 => "00000001010101110110110111010001",
			7022 => "0000000111000000000101110100001000",
			7023 => "0000000110000000001000010000000100",
			7024 => "11111111010001100110110111010001",
			7025 => "00000000000000000110110111010001",
			7026 => "00000000000000000110110111010001",
			7027 => "11111110011101100110110111010001",
			7028 => "0000001100000000000111001000001000",
			7029 => "0000000111000000000110100100000100",
			7030 => "11111110110001010110111011010101",
			7031 => "00000000000000000110111011010101",
			7032 => "0000000010000000001000001101001000",
			7033 => "0000001010000000001010100000100000",
			7034 => "0000000101000000001110101000001000",
			7035 => "0000001100000000001010111000000100",
			7036 => "00000000000000000110111011010101",
			7037 => "00000000011100110110111011010101",
			7038 => "0000000010000000000010000100001100",
			7039 => "0000001000000000001000100100001000",
			7040 => "0000000010000000000110010000000100",
			7041 => "00000000000000000110111011010101",
			7042 => "11111110111010010110111011010101",
			7043 => "00000000000000000110111011010101",
			7044 => "0000000010000000001100000000001000",
			7045 => "0000000001000000001001011000000100",
			7046 => "00000000000000000110111011010101",
			7047 => "00000000111010000110111011010101",
			7048 => "11111111001111110110111011010101",
			7049 => "0000000101000000001101000100011000",
			7050 => "0000000101000000000010110100001100",
			7051 => "0000000111000000000110100100000100",
			7052 => "00000000000000000110111011010101",
			7053 => "0000000000000000000110001000000100",
			7054 => "00000000101101010110111011010101",
			7055 => "00000000000000000110111011010101",
			7056 => "0000001001000000000100101100001000",
			7057 => "0000001011000000000101100100000100",
			7058 => "00000000010001010110111011010101",
			7059 => "00000000000000000110111011010101",
			7060 => "11111111000010110110111011010101",
			7061 => "0000000011000000001011111000001000",
			7062 => "0000000001000000000000111100000100",
			7063 => "00000000000000000110111011010101",
			7064 => "00000001010110110110111011010101",
			7065 => "0000000010000000001010000100000100",
			7066 => "11111111101001010110111011010101",
			7067 => "00000000000000000110111011010101",
			7068 => "0000001110000000000111010100010000",
			7069 => "0000000110000000001101011000000100",
			7070 => "00000000000000000110111011010101",
			7071 => "0000000111000000001001001000000100",
			7072 => "00000000000000000110111011010101",
			7073 => "0000001111000000001000001100000100",
			7074 => "00000000000000000110111011010101",
			7075 => "11111110101100000110111011010101",
			7076 => "0000000010000000001011111000000100",
			7077 => "00000000111100010110111011010101",
			7078 => "0000001110000000001100111000010000",
			7079 => "0000001011000000001010010100001000",
			7080 => "0000000111000000000001101000000100",
			7081 => "00000000000000000110111011010101",
			7082 => "11111111000001110110111011010101",
			7083 => "0000000010000000000001011100000100",
			7084 => "00000000011000110110111011010101",
			7085 => "00000000000000000110111011010101",
			7086 => "0000000110000000001000010000001000",
			7087 => "0000000000000000000001110100000100",
			7088 => "00000000000000000110111011010101",
			7089 => "11111111111000110110111011010101",
			7090 => "0000000000000000001010101100000100",
			7091 => "00000001000000110110111011010101",
			7092 => "00000000000000000110111011010101",
			7093 => "0000000000000000001010101101111100",
			7094 => "0000001011000000000110110101000000",
			7095 => "0000000100000000001100010000010100",
			7096 => "0000001001000000001111000000001100",
			7097 => "0000001000000000000100101100001000",
			7098 => "0000001011000000001110110000000100",
			7099 => "11111111111101010110111111010001",
			7100 => "00000001000000100110111111010001",
			7101 => "11111110111001110110111111010001",
			7102 => "0000000101000000001100100100000100",
			7103 => "00000001100100000110111111010001",
			7104 => "00000000000000000110111111010001",
			7105 => "0000001110000000000111010100011100",
			7106 => "0000000010000000001000001100010000",
			7107 => "0000001110000000000111011000001000",
			7108 => "0000000000000000001001101000000100",
			7109 => "11111111110111110110111111010001",
			7110 => "11111101101101110110111111010001",
			7111 => "0000001100000000000100011000000100",
			7112 => "11111111111001100110111111010001",
			7113 => "00000001101000100110111111010001",
			7114 => "0000000111000000000001101000001000",
			7115 => "0000001100000000001010111000000100",
			7116 => "00000000000000000110111111010001",
			7117 => "11111110001101010110111111010001",
			7118 => "11111011111001000110111111010001",
			7119 => "0000000000000000000111000100001000",
			7120 => "0000001001000000000111101100000100",
			7121 => "11111111100001010110111111010001",
			7122 => "00000001101010000110111111010001",
			7123 => "0000000010000000001000101000000100",
			7124 => "11111110100010100110111111010001",
			7125 => "00000000000000000110111111010001",
			7126 => "0000000101000000001111010000011100",
			7127 => "0000001000000000001000100100000100",
			7128 => "11111110111010100110111111010001",
			7129 => "0000001011000000000101110100010000",
			7130 => "0000001100000000001011000000001000",
			7131 => "0000001100000000000100011000000100",
			7132 => "00000000100000110110111111010001",
			7133 => "11111111101100100110111111010001",
			7134 => "0000001100000000001001110100000100",
			7135 => "00000001111001010110111111010001",
			7136 => "00000000000000000110111111010001",
			7137 => "0000001111000000000110111100000100",
			7138 => "11111111010000110110111111010001",
			7139 => "00000000100110010110111111010001",
			7140 => "0000001000000000000001010100011000",
			7141 => "0000001100000000001001110100001100",
			7142 => "0000000101000000000010011100001000",
			7143 => "0000001001000000000100111100000100",
			7144 => "11111111000110110110111111010001",
			7145 => "00000001000010010110111111010001",
			7146 => "11111110010100100110111111010001",
			7147 => "0000000000000000000111000100001000",
			7148 => "0000001111000000000110111100000100",
			7149 => "11111111010111000110111111010001",
			7150 => "00000001001111010110111111010001",
			7151 => "11111110111110000110111111010001",
			7152 => "0000001011000000001010010100000100",
			7153 => "00000010001000100110111111010001",
			7154 => "00000000000000000110111111010001",
			7155 => "11111110011011000110111111010001",
			7156 => "0000000000000000001010101101111000",
			7157 => "0000000111000000000110100100100100",
			7158 => "0000000100000000001010000100001100",
			7159 => "0000000001000000000000111100001000",
			7160 => "0000000110000000000000111100000100",
			7161 => "00000000000000000111000011000101",
			7162 => "11111111100111100111000011000101",
			7163 => "00000000110001110111000011000101",
			7164 => "0000000110000000001011001100001000",
			7165 => "0000001010000000001010100000000100",
			7166 => "00000000000000000111000011000101",
			7167 => "11111110101001100111000011000101",
			7168 => "0000001010000000001000100100001100",
			7169 => "0000001011000000000000011100000100",
			7170 => "00000000000000000111000011000101",
			7171 => "0000001110000000000111011000000100",
			7172 => "00000000000000000111000011000101",
			7173 => "00000000111111100111000011000101",
			7174 => "11111110111011100111000011000101",
			7175 => "0000000111000000000001101000011100",
			7176 => "0000001110000000000111010100010100",
			7177 => "0000001111000000000000010000010000",
			7178 => "0000001000000000000111110100001000",
			7179 => "0000000101000000000010110100000100",
			7180 => "00000000000000000111000011000101",
			7181 => "11111111100011110111000011000101",
			7182 => "0000001011000000000000011100000100",
			7183 => "00000000000000000111000011000101",
			7184 => "00000001001101100111000011000101",
			7185 => "11111111010001000111000011000101",
			7186 => "0000001010000000001000100100000100",
			7187 => "00000001101101000111000011000101",
			7188 => "00000000000000000111000011000101",
			7189 => "0000001111000000001111010100100000",
			7190 => "0000000111000000001000011000010000",
			7191 => "0000000110000000001101111100001000",
			7192 => "0000000101000000001110101000000100",
			7193 => "00000000000000000111000011000101",
			7194 => "11111111110001010111000011000101",
			7195 => "0000001101000000000101001000000100",
			7196 => "00000000000000000111000011000101",
			7197 => "00000001011100010111000011000101",
			7198 => "0000000000000000000001010100001000",
			7199 => "0000000011000000000110111100000100",
			7200 => "00000001011110010111000011000101",
			7201 => "11111110110100010111000011000101",
			7202 => "0000001110000000000010000100000100",
			7203 => "00000000000000000111000011000101",
			7204 => "00000001010111100111000011000101",
			7205 => "0000001110000000001011111000001100",
			7206 => "0000000000000000000110001000001000",
			7207 => "0000000110000000001101011000000100",
			7208 => "11111110110110100111000011000101",
			7209 => "00000001010101010111000011000101",
			7210 => "11111110000010100111000011000101",
			7211 => "0000001000000000000001010100001000",
			7212 => "0000000001000000000100110100000100",
			7213 => "00000000100010110111000011000101",
			7214 => "11111110101101110111000011000101",
			7215 => "00000001100000110111000011000101",
			7216 => "11111110011100110111000011000101",
			7217 => "0000000000000000001010101110000000",
			7218 => "0000000001000000000000111100111100",
			7219 => "0000000011000000001010000100101100",
			7220 => "0000000010000000001110110100011100",
			7221 => "0000000100000000001100010000001100",
			7222 => "0000000110000000001101111100001000",
			7223 => "0000000110000000000000111100000100",
			7224 => "00000000011111100111000111001011",
			7225 => "11111111001011010111000111001011",
			7226 => "00000001111000100111000111001011",
			7227 => "0000000110000000000100110100001000",
			7228 => "0000001000000000001000100100000100",
			7229 => "11111110000101010111000111001011",
			7230 => "11111111110010100111000111001011",
			7231 => "0000000011000000001100010000000100",
			7232 => "11111111101011010111000111001011",
			7233 => "00000000011101100111000111001011",
			7234 => "0000001011000000000010001000001100",
			7235 => "0000000110000000000100110100000100",
			7236 => "11111110100100110111000111001011",
			7237 => "0000000001000000001001011000000100",
			7238 => "11111111011011010111000111001011",
			7239 => "00000001110110000111000111001011",
			7240 => "00000010010011000111000111001011",
			7241 => "0000001001000000001111000000000100",
			7242 => "11111101111111000111000111001011",
			7243 => "0000000011000000000111010100000100",
			7244 => "00000001000000000111000111001011",
			7245 => "0000001011000000000100010000000100",
			7246 => "11111110011111110111000111001011",
			7247 => "00000000111100000111000111001011",
			7248 => "0000000111000000000001101000100000",
			7249 => "0000000001000000000101011100000100",
			7250 => "00000001011010000111000111001011",
			7251 => "0000001001000000001001111100001100",
			7252 => "0000000010000000000111011000001000",
			7253 => "0000001010000000001010100000000100",
			7254 => "11111110101100000111000111001011",
			7255 => "00000001001011000111000111001011",
			7256 => "11111101111010110111000111001011",
			7257 => "0000001110000000001100010000001000",
			7258 => "0000000100000000000111010100000100",
			7259 => "00000000011001010111000111001011",
			7260 => "11111110100011010111000111001011",
			7261 => "0000000100000000000001011100000100",
			7262 => "00000001010001110111000111001011",
			7263 => "11111111101011110111000111001011",
			7264 => "0000000101000000000111111100011000",
			7265 => "0000001001000000000100111100001000",
			7266 => "0000000100000000000111010100000100",
			7267 => "00000000100001000111000111001011",
			7268 => "11111111110011000111000111001011",
			7269 => "0000001011000000001011011100001000",
			7270 => "0000000100000000000001011100000100",
			7271 => "00000000111101010111000111001011",
			7272 => "11111111100111110111000111001011",
			7273 => "0000000111000000000111010000000100",
			7274 => "00000001101001100111000111001011",
			7275 => "00000000001101110111000111001011",
			7276 => "0000000111000000000101110100001000",
			7277 => "0000000101000000001110010000000100",
			7278 => "00000000000000000111000111001011",
			7279 => "11111110101111010111000111001011",
			7280 => "00000000001101000111000111001011",
			7281 => "11111110011010100111000111001011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(2358, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(4838, initial_addr_3'length));
	end generate gen_rom_2;

	gen_rom_3: if SELECT_ROM = 3 generate
		bank <= (
			0 => "00000000000000000000000000000101",
			1 => "00000000000000000000000000001001",
			2 => "00000000000000000000000000001101",
			3 => "00000000000000000000000000010001",
			4 => "00000000000000000000000000010101",
			5 => "00000000000000000000000000011001",
			6 => "00000000000000000000000000011101",
			7 => "00000000000000000000000000100001",
			8 => "00000000000000000000000000100101",
			9 => "00000000000000000000000000101001",
			10 => "00000000000000000000000000101101",
			11 => "00000000000000000000000000110001",
			12 => "00000000000000000000000000110101",
			13 => "00000000000000000000000000111001",
			14 => "00000000000000000000000000111101",
			15 => "00000000000000000000000001000001",
			16 => "00000000000000000000000001000101",
			17 => "00000000000000000000000001001001",
			18 => "00000000000000000000000001001101",
			19 => "00000000000000000000000001010001",
			20 => "00000000000000000000000001010101",
			21 => "00000000000000000000000001011001",
			22 => "0000000000000000000010101100000100",
			23 => "00000000000000000000000001100101",
			24 => "11111111111010110000000001100101",
			25 => "0000001100000000001100110000000100",
			26 => "11111111111100100000000001110001",
			27 => "00000000000000000000000001110001",
			28 => "0000000010000000001000000000000100",
			29 => "00000000001001010000000001111101",
			30 => "00000000000000000000000001111101",
			31 => "0000000100000000000111001000000100",
			32 => "00000000000000000000000010001001",
			33 => "11111111111111010000000010001001",
			34 => "0000001111000000001011000000000100",
			35 => "00000000000000000000000010010101",
			36 => "11111111111010100000000010010101",
			37 => "0000000100000000000110110100000100",
			38 => "00000000000010110000000010100001",
			39 => "00000000000000000000000010100001",
			40 => "0000000010000000001000000000000100",
			41 => "00000000001011100000000010101101",
			42 => "00000000000000000000000010101101",
			43 => "0000000100000000000111010000000100",
			44 => "00000000101111010000000011000001",
			45 => "0000001001000000001110010100000100",
			46 => "11111111110001100000000011000001",
			47 => "00000000000000000000000011000001",
			48 => "0000001001000000000000111100000100",
			49 => "11111111111001110000000011010101",
			50 => "0000001001000000001001100100000100",
			51 => "00000000000110100000000011010101",
			52 => "00000000000000000000000011010101",
			53 => "0000000000000000000010101100000100",
			54 => "00000000001101000000000011101001",
			55 => "0000001111000000001100010100000100",
			56 => "11111111111101100000000011101001",
			57 => "00000000000000000000000011101001",
			58 => "0000001111000000001001001000001000",
			59 => "0000000000000000000101000100000100",
			60 => "00000000001000100000000011111101",
			61 => "00000000000000000000000011111101",
			62 => "00000000000000000000000011111101",
			63 => "0000000000000000000110011000001000",
			64 => "0000001110000000000010001000000100",
			65 => "00000001110001000000000100010001",
			66 => "11010101110100010000000100010001",
			67 => "11000011110100010000000100010001",
			68 => "0000001010000000001101011000001000",
			69 => "0000001100000000000110000100000100",
			70 => "00000001001101100000000100101101",
			71 => "00000000000000000000000100101101",
			72 => "0000001001000000000101011100000100",
			73 => "11111111111100110000000100101101",
			74 => "00000000000000000000000100101101",
			75 => "0000000010000000001000000000001000",
			76 => "0000000110000000001101011100000100",
			77 => "00000000000000000000000101001001",
			78 => "00000000101010100000000101001001",
			79 => "0000000001000000000111100100000100",
			80 => "11111111110001010000000101001001",
			81 => "00000000000000000000000101001001",
			82 => "0000000010000000001000000000001000",
			83 => "0000001100000000000100000000000100",
			84 => "00000000000000000000000101100101",
			85 => "00000000010101010000000101100101",
			86 => "0000000111000000000111010000000100",
			87 => "11111111101010100000000101100101",
			88 => "00000000000000000000000101100101",
			89 => "0000001001000000000101011100001100",
			90 => "0000000010000000000100001000000100",
			91 => "00000000000000000000000110000001",
			92 => "0000000001000000000110101000000100",
			93 => "11111111100001010000000110000001",
			94 => "00000000000000000000000110000001",
			95 => "00000000000000000000000110000001",
			96 => "0000000001000000000110101000000100",
			97 => "00000000000000000000000110011101",
			98 => "0000001110000000000111110000001000",
			99 => "0000001000000000000111110100000100",
			100 => "00000000011001000000000110011101",
			101 => "00000000000000000000000110011101",
			102 => "00000000000000000000000110011101",
			103 => "0000001001000000000000111100001100",
			104 => "0000001110000000000100001000000100",
			105 => "00000000000000000000000110111001",
			106 => "0000000001000000000110101000000100",
			107 => "11111111110111010000000110111001",
			108 => "00000000000000000000000110111001",
			109 => "00000000000000000000000110111001",
			110 => "0000000100000000000111010000000100",
			111 => "00000000000000000000000111010101",
			112 => "0000000000000000000010101100000100",
			113 => "00000000000000000000000111010101",
			114 => "0000001111000000001010011100000100",
			115 => "00000000000000000000000111010101",
			116 => "11111111111110100000000111010101",
			117 => "0000000000000000000010101100001000",
			118 => "0000001100000000000110000100000100",
			119 => "00000000101110110000000111111001",
			120 => "00000000000000000000000111111001",
			121 => "0000000001000000000111100100001000",
			122 => "0000001100000000001110001100000100",
			123 => "11111111100000000000000111111001",
			124 => "00000000000000000000000111111001",
			125 => "00000000000000000000000111111001",
			126 => "0000000010000000000000110100010000",
			127 => "0000001001000000000000111100001000",
			128 => "0000001110000000000100001000000100",
			129 => "00000000000000000000001000011101",
			130 => "11111111101011100000001000011101",
			131 => "0000001111000000001011011100000100",
			132 => "00000000111001100000001000011101",
			133 => "00000000000000000000001000011101",
			134 => "11111111000011100000001000011101",
			135 => "0000001100000000000100000000001100",
			136 => "0000000100000000000111001000000100",
			137 => "00000000000000000000001001001001",
			138 => "0000000111000000001101100000000100",
			139 => "11111111010011100000001001001001",
			140 => "00000000000000000000001001001001",
			141 => "0000001011000000000100001000001000",
			142 => "0000000000000000000101000100000100",
			143 => "00000000011011100000001001001001",
			144 => "00000000000000000000001001001001",
			145 => "00000000000000000000001001001001",
			146 => "0000001001000000000000111100000100",
			147 => "00000000000000000000001001101101",
			148 => "0000001001000000001001100100001100",
			149 => "0000000111000000000101101100000100",
			150 => "00000000000000000000001001101101",
			151 => "0000000011000000001001100000000100",
			152 => "00000000001010000000001001101101",
			153 => "00000000000000000000001001101101",
			154 => "00000000000000000000001001101101",
			155 => "0000001001000000000000111100000100",
			156 => "00000000000000000000001010010001",
			157 => "0000001001000000001001100100001100",
			158 => "0000001101000000000010011100001000",
			159 => "0000001101000000000110100100000100",
			160 => "00000000000000000000001010010001",
			161 => "00000000001000100000001010010001",
			162 => "00000000000000000000001010010001",
			163 => "00000000000000000000001010010001",
			164 => "0000000100000000000110110100010000",
			165 => "0000001001000000000101011100001100",
			166 => "0000000011000000001010111100000100",
			167 => "00000000000000000000001010111101",
			168 => "0000000111000000001101100000000100",
			169 => "00000000000000000000001010111101",
			170 => "11111111110100100000001010111101",
			171 => "00000000011000100000001010111101",
			172 => "0000001001000000000111101000000100",
			173 => "11111111000111100000001010111101",
			174 => "00000000000000000000001010111101",
			175 => "0000000001000000000110101000010000",
			176 => "0000001111000000000001111100000100",
			177 => "00000000000000000000001011101001",
			178 => "0000001011000000000000001100001000",
			179 => "0000000111000000000110000100000100",
			180 => "11111111011100100000001011101001",
			181 => "00000000000000000000001011101001",
			182 => "00000000000000000000001011101001",
			183 => "0000001111000000001011011100000100",
			184 => "00000001001011110000001011101001",
			185 => "00000000000000000000001011101001",
			186 => "0000000010000000001000000000001000",
			187 => "0000000001000000000110101000000100",
			188 => "00000000000000000000001100010101",
			189 => "00000000101100010000001100010101",
			190 => "0000001001000000000111101000001100",
			191 => "0000000001000000001101101000001000",
			192 => "0000000100000000000001101000000100",
			193 => "00000000000000000000001100010101",
			194 => "11111111101011100000001100010101",
			195 => "00000000000000000000001100010101",
			196 => "00000000000000000000001100010101",
			197 => "0000001100000000001100110000001000",
			198 => "0000001001000000000101011100000100",
			199 => "11111111110100000000001101000001",
			200 => "00000000000000000000001101000001",
			201 => "0000001001000000001001100100001100",
			202 => "0000001100000000001000000000001000",
			203 => "0000001001000000001101011100000100",
			204 => "00000000000000000000001101000001",
			205 => "00000000001101000000001101000001",
			206 => "00000000000000000000001101000001",
			207 => "00000000000000000000001101000001",
			208 => "0000000010000000000000110100010100",
			209 => "0000001001000000000000111100001100",
			210 => "0000001110000000000100001000000100",
			211 => "00000000000000000000001101101101",
			212 => "0000000111000000001101100000000100",
			213 => "00000000000000000000001101101101",
			214 => "11111111100101010000001101101101",
			215 => "0000001111000000001011011100000100",
			216 => "00000000111101110000001101101101",
			217 => "00000000000000000000001101101101",
			218 => "11111111000001000000001101101101",
			219 => "0000001001000000000101011100001100",
			220 => "0000001110000000000100001000000100",
			221 => "00000000000000000000001110100001",
			222 => "0000000001000000000111100100000100",
			223 => "11111111110010100000001110100001",
			224 => "00000000000000000000001110100001",
			225 => "0000000001000000001001011000001100",
			226 => "0000001110000000001010001000001000",
			227 => "0000000111000000001101100000000100",
			228 => "00000000000000000000001110100001",
			229 => "00000000001011110000001110100001",
			230 => "00000000000000000000001110100001",
			231 => "00000000000000000000001110100001",
			232 => "0000000100000000000110110100010100",
			233 => "0000000001000000000110101000001100",
			234 => "0000000011000000001010111100000100",
			235 => "00000000000000000000001111011101",
			236 => "0000000111000000001101100000000100",
			237 => "00000000000000000000001111011101",
			238 => "11111111110101010000001111011101",
			239 => "0000000110000000001001011000000100",
			240 => "00000000000000000000001111011101",
			241 => "00000000010110010000001111011101",
			242 => "0000000111000000001100101000001000",
			243 => "0000001100000000001110001100000100",
			244 => "11111111001011010000001111011101",
			245 => "00000000000000000000001111011101",
			246 => "00000000000000000000001111011101",
			247 => "0000001001000000000000111100010000",
			248 => "0000000100000000000111001000000100",
			249 => "00000000000000000000010000011001",
			250 => "0000000001000000000110101000001000",
			251 => "0000000111000000001110001100000100",
			252 => "11111111100111100000010000011001",
			253 => "00000000000000000000010000011001",
			254 => "00000000000000000000010000011001",
			255 => "0000001010000000000111101100001100",
			256 => "0000001110000000001010001000001000",
			257 => "0000000001000000000111100100000100",
			258 => "00000000000000000000010000011001",
			259 => "00000000011001100000010000011001",
			260 => "00000000000000000000010000011001",
			261 => "00000000000000000000010000011001",
			262 => "0000001000000000000111110100011000",
			263 => "0000001001000000000000111100001100",
			264 => "0000001111000000001011000000001000",
			265 => "0000000111000000001001110000000100",
			266 => "00000000000000000000010001001101",
			267 => "00000000100000000000010001001101",
			268 => "11111111101101010000010001001101",
			269 => "0000000111000000000110000100000100",
			270 => "00000000000000000000010001001101",
			271 => "0000000011000000001001100000000100",
			272 => "00000000111000010000010001001101",
			273 => "00000000000000000000010001001101",
			274 => "11111111010000100000010001001101",
			275 => "0000001011000000000101101100001000",
			276 => "0000000100000000000111001000000100",
			277 => "00000000000000000000010010000001",
			278 => "11111111100110000000010010000001",
			279 => "0000000100000000001001100000010000",
			280 => "0000001001000000000000111100000100",
			281 => "00000000000000000000010010000001",
			282 => "0000001110000000001010001000001000",
			283 => "0000000001000000001001011000000100",
			284 => "00000000010011000000010010000001",
			285 => "00000000000000000000010010000001",
			286 => "00000000000000000000010010000001",
			287 => "00000000000000000000010010000001",
			288 => "0000001001000000000000111100001000",
			289 => "0000001100000000000110000100000100",
			290 => "11111111111010100000010010110101",
			291 => "00000000000000000000010010110101",
			292 => "0000001001000000001001100100010000",
			293 => "0000000101000000001110101000001100",
			294 => "0000000111000000001101100000000100",
			295 => "00000000000000000000010010110101",
			296 => "0000001100000000001000000000000100",
			297 => "00000000001001110000010010110101",
			298 => "00000000000000000000010010110101",
			299 => "00000000000000000000010010110101",
			300 => "00000000000000000000010010110101",
			301 => "0000000000000000000010101100000100",
			302 => "00000000011110000000010011100001",
			303 => "0000000001000000000111100100000100",
			304 => "11111111010111010000010011100001",
			305 => "0000000010000000001110010000001100",
			306 => "0000000110000000001101111100001000",
			307 => "0000000101000000001101000100000100",
			308 => "00000000001101100000010011100001",
			309 => "00000000000000000000010011100001",
			310 => "00000000000000000000010011100001",
			311 => "00000000000000000000010011100001",
			312 => "0000000000000000000110011000010100",
			313 => "0000001100000000000100000000000100",
			314 => "11111111110000100000010100011101",
			315 => "0000001111000000000001001000001100",
			316 => "0000000001000000000111100100001000",
			317 => "0000000011000000000110100100000100",
			318 => "00000001101100100000010100011101",
			319 => "11111101111011100000010100011101",
			320 => "00000001110000010000010100011101",
			321 => "11111111100011000000010100011101",
			322 => "0000000100000000001100010100001000",
			323 => "0000001010000000000100101100000100",
			324 => "11111110101001000000010100011101",
			325 => "00000011010010010000010100011101",
			326 => "11111110011001010000010100011101",
			327 => "0000001100000000001100110000001100",
			328 => "0000001010000000000100110100000100",
			329 => "00000000000000000000010101011001",
			330 => "0000000001000000000111100100000100",
			331 => "11111111101010100000010101011001",
			332 => "00000000000000000000010101011001",
			333 => "0000000001000000000110101000000100",
			334 => "00000000000000000000010101011001",
			335 => "0000000010000000001110010000001100",
			336 => "0000000001000000001001011000001000",
			337 => "0000000011000000001001100000000100",
			338 => "00000000100000110000010101011001",
			339 => "00000000000000000000010101011001",
			340 => "00000000000000000000010101011001",
			341 => "00000000000000000000010101011001",
			342 => "0000000000000000000110011000011000",
			343 => "0000001111000000001011000000001000",
			344 => "0000001011000000000101101100000100",
			345 => "00000000001100010000010110001101",
			346 => "00000001100110100000010110001101",
			347 => "0000001001000000000101011100000100",
			348 => "11111101100110100000010110001101",
			349 => "0000001111000000000010001000000100",
			350 => "00000001100110100000010110001101",
			351 => "0000001001000000001101111100000100",
			352 => "11111110000001010000010110001101",
			353 => "00000001010000000000010110001101",
			354 => "11111110011001110000010110001101",
			355 => "0000001010000000001001111100011000",
			356 => "0000000011000000000001001000010100",
			357 => "0000001100000000000100000000001000",
			358 => "0000000100000000000111001000000100",
			359 => "00000010100000100000010111010001",
			360 => "11111111010110110000010111010001",
			361 => "0000001111000000000010001000001000",
			362 => "0000000010000000000001101000000100",
			363 => "00000010100001110000010111010001",
			364 => "00000010010000110000010111010001",
			365 => "00000000100110100000010111010001",
			366 => "00000110101100000000010111010001",
			367 => "0000000100000000001100010100001000",
			368 => "0000000100000000001110010000000100",
			369 => "11111110011101000000010111010001",
			370 => "11111111110110010000010111010001",
			371 => "11111110010111110000010111010001",
			372 => "0000001100000000001100110000010000",
			373 => "0000000010000000000100001000000100",
			374 => "00000000000000000000011000010101",
			375 => "0000001001000000000101011100001000",
			376 => "0000001101000000001111011100000100",
			377 => "11111111101011110000011000010101",
			378 => "00000000000000000000011000010101",
			379 => "00000000000000000000011000010101",
			380 => "0000001001000000000000111100000100",
			381 => "00000000000000000000011000010101",
			382 => "0000000010000000001110010000001100",
			383 => "0000001001000000001001100100001000",
			384 => "0000000101000000001110101000000100",
			385 => "00000000011101000000011000010101",
			386 => "00000000000000000000011000010101",
			387 => "00000000000000000000011000010101",
			388 => "00000000000000000000011000010101",
			389 => "0000000000000000000110011000011000",
			390 => "0000000001000000001001111000000100",
			391 => "11111111001100100000011001100001",
			392 => "0000001111000000000010001000001100",
			393 => "0000001100000000001000111000001000",
			394 => "0000000011000000000011100000000100",
			395 => "00000001101101110000011001100001",
			396 => "11111111001100000000011001100001",
			397 => "00000001101001000000011001100001",
			398 => "0000000111000000000100001000000100",
			399 => "11111101101001010000011001100001",
			400 => "00000001111010010000011001100001",
			401 => "0000000100000000001001100000001100",
			402 => "0000001010000000000111101100000100",
			403 => "11111110011111100000011001100001",
			404 => "0000001000000000000111110100000100",
			405 => "00000100000100110000011001100001",
			406 => "11111111101110100000011001100001",
			407 => "11111110011001010000011001100001",
			408 => "0000000001000000000111100100011000",
			409 => "0000001111000000001011000000001100",
			410 => "0000001100000000000100000000000100",
			411 => "00000000000000000000011010110101",
			412 => "0000000110000000000111101000000100",
			413 => "00000000001010010000011010110101",
			414 => "00000000000000000000011010110101",
			415 => "0000001100000000001110001100001000",
			416 => "0000000110000000001001011000000100",
			417 => "00000000000000000000011010110101",
			418 => "11111111000101100000011010110101",
			419 => "00000000000000000000011010110101",
			420 => "0000000010000000001110010000010000",
			421 => "0000000110000000000000111100000100",
			422 => "00000000000000000000011010110101",
			423 => "0000000001000000001001011000001000",
			424 => "0000000101000000001110101000000100",
			425 => "00000000100101110000011010110101",
			426 => "00000000000000000000011010110101",
			427 => "00000000000000000000011010110101",
			428 => "00000000000000000000011010110101",
			429 => "0000000100000000001100010100100000",
			430 => "0000000001000000000111100100010000",
			431 => "0000000100000000001001001000001000",
			432 => "0000000110000000001111001100000100",
			433 => "00000000000000000000011011111001",
			434 => "00000001010011000000011011111001",
			435 => "0000000001000000000110101000000100",
			436 => "11111110101110010000011011111001",
			437 => "11111111110111110000011011111001",
			438 => "0000001111000000000010001000000100",
			439 => "00000001010111010000011011111001",
			440 => "0000001101000000000101110100000100",
			441 => "11111111110000010000011011111001",
			442 => "0000001111000000001010001000000100",
			443 => "00000000100101110000011011111001",
			444 => "00000000000000000000011011111001",
			445 => "11111110011100100000011011111001",
			446 => "0000001011000000000101101100001000",
			447 => "0000000100000000000111001000000100",
			448 => "00000000000000000000011100111101",
			449 => "11111111010010110000011100111101",
			450 => "0000000100000000000111010000000100",
			451 => "00000000011100010000011100111101",
			452 => "0000001100000000001000000000001100",
			453 => "0000001100000000001000111100000100",
			454 => "00000000000000000000011100111101",
			455 => "0000001100000000000110000100000100",
			456 => "11111111101001100000011100111101",
			457 => "00000000000000000000011100111101",
			458 => "0000001100000000001000000000001000",
			459 => "0000001011000000000101100100000100",
			460 => "00000000000000000000011100111101",
			461 => "00000000001111010000011100111101",
			462 => "00000000000000000000011100111101",
			463 => "0000001011000000000101101100001000",
			464 => "0000000100000000000111001000000100",
			465 => "00000000000000000000011110001001",
			466 => "11111111010000010000011110001001",
			467 => "0000001111000000001010011100001000",
			468 => "0000000000000000001100000100000100",
			469 => "00000000100000010000011110001001",
			470 => "00000000000000000000011110001001",
			471 => "0000000001000000000111100100001000",
			472 => "0000001100000000001110001100000100",
			473 => "11111111101010000000011110001001",
			474 => "00000000000000000000011110001001",
			475 => "0000001000000000000111110100001100",
			476 => "0000001110000000001010001000001000",
			477 => "0000001000000000000100101100000100",
			478 => "00000000000000000000011110001001",
			479 => "00000000010101100000011110001001",
			480 => "00000000000000000000011110001001",
			481 => "00000000000000000000011110001001",
			482 => "0000001000000000000111110100100100",
			483 => "0000000001000000000111100100010100",
			484 => "0000001000000000000101010000001100",
			485 => "0000001110000000000100001000000100",
			486 => "00000000011111010000011111010101",
			487 => "0000000111000000001101100000000100",
			488 => "11111111100110110000011111010101",
			489 => "00000000000000000000011111010101",
			490 => "0000001100000000000011011100000100",
			491 => "00000000000000000000011111010101",
			492 => "11111111001110000000011111010101",
			493 => "0000001110000000001010001000001100",
			494 => "0000000101000000001110101000001000",
			495 => "0000000010000000001110010000000100",
			496 => "00000000100101110000011111010101",
			497 => "00000000000000000000011111010101",
			498 => "00000000000000000000011111010101",
			499 => "00000000000000000000011111010101",
			500 => "11111110110100010000011111010101",
			501 => "0000000100000000001100010100011100",
			502 => "0000000001000000000010001100000100",
			503 => "11111110111111100000100000010001",
			504 => "0000001111000000001011000000000100",
			505 => "00000001100011010000100000010001",
			506 => "0000000111000000000110000100001100",
			507 => "0000000001000000000111100100000100",
			508 => "11111110100111010000100000010001",
			509 => "0000001100000000000011011100000100",
			510 => "00000000010010110000100000010001",
			511 => "11111111101111110000100000010001",
			512 => "0000001111000000001010001000000100",
			513 => "00000001010010000000100000010001",
			514 => "00000000000000000000100000010001",
			515 => "11111110011010100000100000010001",
			516 => "0000001000000000000111110100100100",
			517 => "0000000001000000000111100100010000",
			518 => "0000000000000000000010101100001100",
			519 => "0000000001000000001001111000000100",
			520 => "00000000000000000000100001011101",
			521 => "0000000001000000000110101000000100",
			522 => "00000000111101010000100001011101",
			523 => "00000000000000000000100001011101",
			524 => "11111111000110100000100001011101",
			525 => "0000001111000000000010001000000100",
			526 => "00000000111101110000100001011101",
			527 => "0000001100000000001000000000000100",
			528 => "11111111101110010000100001011101",
			529 => "0000000000000000001100011100000100",
			530 => "00000000000000000000100001011101",
			531 => "0000000010000000001100010100000100",
			532 => "00000000101001000000100001011101",
			533 => "00000000000000000000100001011101",
			534 => "11111110100111010000100001011101",
			535 => "0000001000000000000111110100101000",
			536 => "0000000001000000000111100100010100",
			537 => "0000001110000000000100001000001000",
			538 => "0000000110000000001001011000000100",
			539 => "00000000001011100000100010110001",
			540 => "00000000000000000000100010110001",
			541 => "0000000001000000000110101000000100",
			542 => "11111111010011110000100010110001",
			543 => "0000000110000000000000111100000100",
			544 => "00000000000001100000100010110001",
			545 => "11111111111111100000100010110001",
			546 => "0000001110000000001010001000010000",
			547 => "0000000110000000000000111100000100",
			548 => "00000000000000000000100010110001",
			549 => "0000001100000000001100110000000100",
			550 => "00000000000000000000100010110001",
			551 => "0000000101000000001101000100000100",
			552 => "00000000101010000000100010110001",
			553 => "00000000000000000000100010110001",
			554 => "00000000000000000000100010110001",
			555 => "11111111000001110000100010110001",
			556 => "0000000000000000000110011100011100",
			557 => "0000001100000000000100000000000100",
			558 => "11111111100000100000100011101101",
			559 => "0000000100000000000111010000000100",
			560 => "00000001000010010000100011101101",
			561 => "0000001100000000001100110000000100",
			562 => "11111111100011110000100011101101",
			563 => "0000001110000000001010001000001100",
			564 => "0000001001000000000111101000000100",
			565 => "00000000000000000000100011101101",
			566 => "0000000011000000001001100000000100",
			567 => "00000000111001000000100011101101",
			568 => "00000000000000000000100011101101",
			569 => "00000000000000000000100011101101",
			570 => "11111110100010010000100011101101",
			571 => "0000000000000000000110011100100100",
			572 => "0000000111000000000001101000011100",
			573 => "0000000010000000000000110100011000",
			574 => "0000001001000000000000111100001100",
			575 => "0000000100000000001001001000001000",
			576 => "0000001100000000000100000000000100",
			577 => "11111111111101110000100100111001",
			578 => "00000001011001000000100100111001",
			579 => "11111110010110100000100100111001",
			580 => "0000001111000000000010001000000100",
			581 => "00000001100001010000100100111001",
			582 => "0000000101000000001011011100000100",
			583 => "11111111011000110000100100111001",
			584 => "00000001001010100000100100111001",
			585 => "11111110111001010000100100111001",
			586 => "0000000010000000001110010000000100",
			587 => "00000011100001000000100100111001",
			588 => "00000000000000000000100100111001",
			589 => "11111110011011010000100100111001",
			590 => "0000000100000000001100010100100000",
			591 => "0000000001000000000010001100000100",
			592 => "11111110000000000000100101111101",
			593 => "0000000010000000000001001000010100",
			594 => "0000000001000000000110101000010000",
			595 => "0000001111000000000111001000001100",
			596 => "0000001110000000000100001000000100",
			597 => "00000001101101010000100101111101",
			598 => "0000001110000000000001111100000100",
			599 => "00000000000000000000100101111101",
			600 => "00000001001111000000100101111101",
			601 => "11111101110010110000100101111101",
			602 => "00000001100111000000100101111101",
			603 => "0000001001000000001101011000000100",
			604 => "11111110100010110000100101111101",
			605 => "00000100011100110000100101111101",
			606 => "11111110011001100000100101111101",
			607 => "0000000000000000000110011100101000",
			608 => "0000001100000000001000000000011100",
			609 => "0000000010000000000000110100011000",
			610 => "0000001001000000000000111100001100",
			611 => "0000000100000000001001001000001000",
			612 => "0000001100000000000100000000000100",
			613 => "00000000000000000000100111010001",
			614 => "00000001010111100000100111010001",
			615 => "11111110100010000000100111010001",
			616 => "0000001110000000000101100100000100",
			617 => "00000001100000000000100111010001",
			618 => "0000000111000000000001111100000100",
			619 => "11111110111010100000100111010001",
			620 => "00000001001111110000100111010001",
			621 => "11111110111101100000100111010001",
			622 => "0000001011000000000101100100000100",
			623 => "00000000000000000000100111010001",
			624 => "0000000101000000001110101000000100",
			625 => "00000010111100110000100111010001",
			626 => "00000000000000000000100111010001",
			627 => "11111110011011100000100111010001",
			628 => "0000000000000000000110011100100100",
			629 => "0000000111000000000001101000011100",
			630 => "0000001111000000000000110100011000",
			631 => "0000001100000000000100000000001000",
			632 => "0000000100000000000111001000000100",
			633 => "00000000111010110000101000011101",
			634 => "11111110101011000000101000011101",
			635 => "0000001100000000000011011100000100",
			636 => "00000001011100000000101000011101",
			637 => "0000000001000000000111100100001000",
			638 => "0000000011000000000110100100000100",
			639 => "00000000110010000000101000011101",
			640 => "11111111000100010000101000011101",
			641 => "00000001010111000000101000011101",
			642 => "11111111000010000000101000011101",
			643 => "0000000011000000001001100000000100",
			644 => "00000010100001110000101000011101",
			645 => "00000000000000000000101000011101",
			646 => "11111110011011110000101000011101",
			647 => "0000001000000000000111110100100100",
			648 => "0000000001000000001001111000001000",
			649 => "0000001111000000000000001100000100",
			650 => "00000000000000000000101001101001",
			651 => "11111111000010110000101001101001",
			652 => "0000001011000000000100001000000100",
			653 => "00000001010010110000101001101001",
			654 => "0000001100000000001100110000001000",
			655 => "0000001111000000001010011100000100",
			656 => "00000000000000000000101001101001",
			657 => "11111110111101110000101001101001",
			658 => "0000001110000000001010001000001100",
			659 => "0000000001000000000111100100000100",
			660 => "00000000000000000000101001101001",
			661 => "0000000110000000000000111100000100",
			662 => "00000000000000000000101001101001",
			663 => "00000000111111110000101001101001",
			664 => "00000000000000000000101001101001",
			665 => "11111110100001100000101001101001",
			666 => "0000000000000000000110011100101100",
			667 => "0000000001000000000111100100010100",
			668 => "0000000000000000000010101100001100",
			669 => "0000001100000000000100000000000100",
			670 => "11111111011111010000101011000101",
			671 => "0000001100000000000110000100000100",
			672 => "00000001010000110000101011000101",
			673 => "00000000000000000000101011000101",
			674 => "0000000001000000000111100100000100",
			675 => "11111110100010110000101011000101",
			676 => "00000000000000000000101011000101",
			677 => "0000000110000000000000111100000100",
			678 => "00000000000000000000101011000101",
			679 => "0000000010000000001110010000010000",
			680 => "0000001100000000001100110000000100",
			681 => "00000000000000000000101011000101",
			682 => "0000000001000000001001011000001000",
			683 => "0000000101000000001101000100000100",
			684 => "00000001010110010000101011000101",
			685 => "00000000000000000000101011000101",
			686 => "00000000000000000000101011000101",
			687 => "00000000000000000000101011000101",
			688 => "11111110011110110000101011000101",
			689 => "0000000000000000000110011100101000",
			690 => "0000001100000000000100000000000100",
			691 => "11111111101010000000101100011011",
			692 => "0000001111000000001010011100001100",
			693 => "0000001001000000000000111100001000",
			694 => "0000001001000000000000111100000100",
			695 => "00000000011011100000101100011011",
			696 => "00000000000000000000101100011011",
			697 => "00000001001100100000101100011011",
			698 => "0000001010000000001001100100001000",
			699 => "0000000001000000001101101000000100",
			700 => "11111111010100010000101100011011",
			701 => "00000000000000000000101100011011",
			702 => "0000001110000000001010001000001100",
			703 => "0000001100000000001100110000000100",
			704 => "00000000000000000000101100011011",
			705 => "0000000011000000001001100000000100",
			706 => "00000000101111000000101100011011",
			707 => "00000000000000000000101100011011",
			708 => "00000000000000000000101100011011",
			709 => "11111110100100000000101100011011",
			710 => "00000000000000000000101100011101",
			711 => "00000000000000000000101100100001",
			712 => "00000000000000000000101100100101",
			713 => "00000000000000000000101100101001",
			714 => "00000000000000000000101100101101",
			715 => "00000000000000000000101100110001",
			716 => "00000000000000000000101100110101",
			717 => "00000000000000000000101100111001",
			718 => "00000000000000000000101100111101",
			719 => "00000000000000000000101101000001",
			720 => "00000000000000000000101101000101",
			721 => "00000000000000000000101101001001",
			722 => "00000000000000000000101101001101",
			723 => "00000000000000000000101101010001",
			724 => "00000000000000000000101101010101",
			725 => "00000000000000000000101101011001",
			726 => "00000000000000000000101101011101",
			727 => "00000000000000000000101101100001",
			728 => "00000000000000000000101101100101",
			729 => "00000000000000000000101101101001",
			730 => "00000000000000000000101101101101",
			731 => "00000000000000000000101101110001",
			732 => "0000000000000000000010101100000100",
			733 => "00000000000000000000101101111101",
			734 => "11111111111101010000101101111101",
			735 => "0000001100000000001100110000000100",
			736 => "11111111111101100000101110001001",
			737 => "00000000000000000000101110001001",
			738 => "0000000010000000001000000000000100",
			739 => "00000000001001000000101110010101",
			740 => "00000000000000000000101110010101",
			741 => "0000000100000000000111001000000100",
			742 => "00000000000000000000101110100001",
			743 => "11111111111111100000101110100001",
			744 => "0000001111000000001011000000000100",
			745 => "00000000000000000000101110101101",
			746 => "11111111111011100000101110101101",
			747 => "0000000100000000000110110100000100",
			748 => "00000000000010000000101110111001",
			749 => "00000000000000000000101110111001",
			750 => "0000000010000000001000000000000100",
			751 => "00000000001010110000101111000101",
			752 => "00000000000000000000101111000101",
			753 => "0000000010000000000001101000000100",
			754 => "00000000101011100000101111011001",
			755 => "0000001001000000001110010100000100",
			756 => "11111111110011100000101111011001",
			757 => "00000000000000000000101111011001",
			758 => "0000001001000000000000111100000100",
			759 => "11111111111011000000101111101101",
			760 => "0000001001000000001001100100000100",
			761 => "00000000000101000000101111101101",
			762 => "00000000000000000000101111101101",
			763 => "0000000000000000000010101100000100",
			764 => "00000000001011110000110000000001",
			765 => "0000001111000000001100010100000100",
			766 => "11111111111111000000110000000001",
			767 => "00000000000000000000110000000001",
			768 => "0000001100000000001000000000001000",
			769 => "0000000011000000001100101100000100",
			770 => "00000000000000000000110000010101",
			771 => "11111111111101110000110000010101",
			772 => "00000000000000000000110000010101",
			773 => "0000001010000000001101011000001000",
			774 => "0000001100000000000110000100000100",
			775 => "00000001011011100000110000110001",
			776 => "00000000000000000000110000110001",
			777 => "0000001001000000000101011100000100",
			778 => "11111111111100000000110000110001",
			779 => "00000000000000000000110000110001",
			780 => "0000001001000000000000111100001000",
			781 => "0000000100000000000111001000000100",
			782 => "00000000000000000000110001001101",
			783 => "11111111100110000000110001001101",
			784 => "0000001111000000000111010000000100",
			785 => "00000000110001110000110001001101",
			786 => "00000000000000000000110001001101",
			787 => "0000000010000000001000000000001000",
			788 => "0000001100000000000100000000000100",
			789 => "00000000000000000000110001101001",
			790 => "00000000100101000000110001101001",
			791 => "0000001100000000001100110000000100",
			792 => "11111111111000110000110001101001",
			793 => "00000000000000000000110001101001",
			794 => "0000000010000000001000000000001000",
			795 => "0000001100000000000100000000000100",
			796 => "00000000000000000000110010000101",
			797 => "00000000010011100000110010000101",
			798 => "0000001001000000000111101000000100",
			799 => "11111111101011010000110010000101",
			800 => "00000000000000000000110010000101",
			801 => "0000001001000000000101011100001100",
			802 => "0000000010000000000100001000000100",
			803 => "00000000000000000000110010100001",
			804 => "0000000001000000000110101000000100",
			805 => "11111111100101000000110010100001",
			806 => "00000000000000000000110010100001",
			807 => "00000000000000000000110010100001",
			808 => "0000000001000000000110101000000100",
			809 => "00000000000000000000110010111101",
			810 => "0000001110000000000111110000001000",
			811 => "0000000111000000001101100000000100",
			812 => "00000000000000000000110010111101",
			813 => "00000000010100110000110010111101",
			814 => "00000000000000000000110010111101",
			815 => "0000000100000000000111010000000100",
			816 => "00000000000000000000110011011001",
			817 => "0000000000000000000010101100000100",
			818 => "00000000000000000000110011011001",
			819 => "0000001111000000001010011100000100",
			820 => "00000000000000000000110011011001",
			821 => "11111111111101110000110011011001",
			822 => "0000000000000000000010101100001000",
			823 => "0000001100000000000110000100000100",
			824 => "00000000101010100000110011111101",
			825 => "00000000000000000000110011111101",
			826 => "0000000001000000000111100100001000",
			827 => "0000001100000000001110001100000100",
			828 => "11111111001011100000110011111101",
			829 => "00000000000000000000110011111101",
			830 => "00000000000000000000110011111101",
			831 => "0000000000000000000010101100001000",
			832 => "0000001100000000000110000100000100",
			833 => "00000000101100100000110100100001",
			834 => "00000000000000000000110100100001",
			835 => "0000000001000000000111100100001000",
			836 => "0000001100000000001110001100000100",
			837 => "11111111100001110000110100100001",
			838 => "00000000000000000000110100100001",
			839 => "00000000000000000000110100100001",
			840 => "0000000010000000000000110100010000",
			841 => "0000000001000000000111100100001000",
			842 => "0000001000000000001001111100000100",
			843 => "00000000000000000000110101000101",
			844 => "11111111111001000000110101000101",
			845 => "0000001110000000001101010100000100",
			846 => "00000000000000000000110101000101",
			847 => "00000000010111100000110101000101",
			848 => "11111111100011010000110101000101",
			849 => "0000001111000000001001001000001100",
			850 => "0000001100000000000100000000000100",
			851 => "00000000000000000000110101110001",
			852 => "0000000000000000001010000000000100",
			853 => "00000000101000010000110101110001",
			854 => "00000000000000000000110101110001",
			855 => "0000001001000000000111101000001000",
			856 => "0000000001000000001101101000000100",
			857 => "11111111110100000000110101110001",
			858 => "00000000000000000000110101110001",
			859 => "00000000000000000000110101110001",
			860 => "0000001001000000000000111100000100",
			861 => "00000000000000000000110110010101",
			862 => "0000001001000000001001100100001100",
			863 => "0000001101000000000010011100001000",
			864 => "0000001101000000001001110100000100",
			865 => "00000000000000000000110110010101",
			866 => "00000000001010110000110110010101",
			867 => "00000000000000000000110110010101",
			868 => "00000000000000000000110110010101",
			869 => "0000001001000000000000111100000100",
			870 => "11111111111010010000110110111001",
			871 => "0000001001000000001001100100001100",
			872 => "0000001101000000000010011100001000",
			873 => "0000001101000000000110100100000100",
			874 => "00000000000000000000110110111001",
			875 => "00000000000101000000110110111001",
			876 => "00000000000000000000110110111001",
			877 => "00000000000000000000110110111001",
			878 => "0000001011000000000101101100001000",
			879 => "0000001010000000000100110100000100",
			880 => "00000000000000000000110111100101",
			881 => "11111111100111110000110111100101",
			882 => "0000000000000000000110011100001100",
			883 => "0000001001000000000000111100000100",
			884 => "00000000000000000000110111100101",
			885 => "0000001110000000001010001000000100",
			886 => "00000000010001000000110111100101",
			887 => "00000000000000000000110111100101",
			888 => "00000000000000000000110111100101",
			889 => "0000000001000000000110101000010000",
			890 => "0000000010000000000100001000000100",
			891 => "00000000000000000000111000010001",
			892 => "0000001011000000000000001100001000",
			893 => "0000000111000000000110000100000100",
			894 => "11111111011111110000111000010001",
			895 => "00000000000000000000111000010001",
			896 => "00000000000000000000111000010001",
			897 => "0000000100000000000110110100000100",
			898 => "00000001000110000000111000010001",
			899 => "00000000000000000000111000010001",
			900 => "0000001100000000001100110000001000",
			901 => "0000000001000000000111100100000100",
			902 => "11111111101111000000111000111101",
			903 => "00000000000000000000111000111101",
			904 => "0000000001000000001001011000001100",
			905 => "0000001100000000001000000000001000",
			906 => "0000001001000000001101011100000100",
			907 => "00000000000000000000111000111101",
			908 => "00000000010010110000111000111101",
			909 => "00000000000000000000111000111101",
			910 => "00000000000000000000111000111101",
			911 => "0000000001000000000110101000001000",
			912 => "0000001011000000000000001100000100",
			913 => "11111111110110000000111001101001",
			914 => "00000000000000000000111001101001",
			915 => "0000000001000000001001011000001100",
			916 => "0000000101000000001101000100001000",
			917 => "0000000101000000000011100000000100",
			918 => "00000000000000000000111001101001",
			919 => "00000000000011100000111001101001",
			920 => "00000000000000000000111001101001",
			921 => "00000000000000000000111001101001",
			922 => "0000000000000000000110011000010100",
			923 => "0000001001000000000000111100001100",
			924 => "0000001110000000000100001000000100",
			925 => "00000000000000000000111010010101",
			926 => "0000000111000000001101100000000100",
			927 => "00000000000000000000111010010101",
			928 => "11111111101101000000111010010101",
			929 => "0000001111000000001011011100000100",
			930 => "00000000110101100000111010010101",
			931 => "00000000000000000000111010010101",
			932 => "11111111000111010000111010010101",
			933 => "0000000001000000000110101000001100",
			934 => "0000000011000000000100001000000100",
			935 => "00000000000000000000111011001001",
			936 => "0000000111000000000110000100000100",
			937 => "11111111101110100000111011001001",
			938 => "00000000000000000000111011001001",
			939 => "0000000001000000001001011000001100",
			940 => "0000000011000000001001100000001000",
			941 => "0000000111000000001001110000000100",
			942 => "00000000000000000000111011001001",
			943 => "00000000000101110000111011001001",
			944 => "00000000000000000000111011001001",
			945 => "00000000000000000000111011001001",
			946 => "0000000000000000000110011000010100",
			947 => "0000001110000000000100010000010000",
			948 => "0000001100000000000100000000001000",
			949 => "0000001111000000001101111000000100",
			950 => "00000010001001010000111011110101",
			951 => "00000000001111110000111011110101",
			952 => "0000001111000000001011011100000100",
			953 => "00000010110010110000111011110101",
			954 => "00000001110010010000111011110101",
			955 => "00000110110000100000111011110101",
			956 => "11111110010111110000111011110101",
			957 => "0000000010000000000001001000010100",
			958 => "0000000100000000001001001000000100",
			959 => "00000000101000100000111100101001",
			960 => "0000000001000000000111100100001100",
			961 => "0000000111000000001110001100001000",
			962 => "0000000110000000001001011000000100",
			963 => "00000000000000000000111100101001",
			964 => "11111111001111100000111100101001",
			965 => "00000000000000000000111100101001",
			966 => "00000000100101000000111100101001",
			967 => "0000000111000000000111010000000100",
			968 => "11111110110111000000111100101001",
			969 => "00000000000000000000111100101001",
			970 => "0000000100000000000110110100010100",
			971 => "0000001001000000000101011100010000",
			972 => "0000000011000000001010111100000100",
			973 => "00000000000000000000111101011101",
			974 => "0000000001000000000110101000001000",
			975 => "0000000111000000001101100000000100",
			976 => "00000000000000000000111101011101",
			977 => "11111111101101100000111101011101",
			978 => "00000000000000000000111101011101",
			979 => "00000000011011000000111101011101",
			980 => "0000001001000000000111101000000100",
			981 => "11111111000100100000111101011101",
			982 => "00000000000000000000111101011101",
			983 => "0000000001000000000110101000001000",
			984 => "0000001011000000000000001100000100",
			985 => "11111111110110100000111110010001",
			986 => "00000000000000000000111110010001",
			987 => "0000000001000000001001011000010000",
			988 => "0000000101000000001110101000001100",
			989 => "0000001100000000001000000000001000",
			990 => "0000000101000000000011100000000100",
			991 => "00000000000000000000111110010001",
			992 => "00000000000100010000111110010001",
			993 => "00000000000000000000111110010001",
			994 => "00000000000000000000111110010001",
			995 => "00000000000000000000111110010001",
			996 => "0000000100000000001100010100010100",
			997 => "0000000100000000001001001000000100",
			998 => "00000000100101100000111110111101",
			999 => "0000001001000000000000111100000100",
			1000 => "11111111001110010000111110111101",
			1001 => "0000001111000000001010011100000100",
			1002 => "00000000101100110000111110111101",
			1003 => "0000000001000000000111100100000100",
			1004 => "11111111100000110000111110111101",
			1005 => "00000000000011000000111110111101",
			1006 => "11111110111011110000111110111101",
			1007 => "0000000000000000000110011000011000",
			1008 => "0000000100000000000110110100001100",
			1009 => "0000001110000000001011000000000100",
			1010 => "00000001110110000001000000000001",
			1011 => "0000001101000000001111011100000100",
			1012 => "11111111100001110001000000000001",
			1013 => "00000001101111100001000000000001",
			1014 => "0000001100000000000110000100000100",
			1015 => "11111100110001100001000000000001",
			1016 => "0000000001000000001011101000000100",
			1017 => "00000000111111110001000000000001",
			1018 => "00000010010100000001000000000001",
			1019 => "0000000100000000001100010100001000",
			1020 => "0000000000000000001100011100000100",
			1021 => "11111110100001010001000000000001",
			1022 => "00000101101101010001000000000001",
			1023 => "11111110011001000001000000000001",
			1024 => "0000000001000000000110101000001100",
			1025 => "0000001011000000000000001100001000",
			1026 => "0000000111000000000110000100000100",
			1027 => "11111111110100000001000000111101",
			1028 => "00000000000000000001000000111101",
			1029 => "00000000000000000001000000111101",
			1030 => "0000000001000000001001011000010000",
			1031 => "0000000101000000001110101000001100",
			1032 => "0000001100000000001000000000001000",
			1033 => "0000000111000000001001110000000100",
			1034 => "00000000000000000001000000111101",
			1035 => "00000000000101000001000000111101",
			1036 => "00000000000000000001000000111101",
			1037 => "00000000000000000001000000111101",
			1038 => "00000000000000000001000000111101",
			1039 => "0000000001000000000110101000001100",
			1040 => "0000001110000000000100001000000100",
			1041 => "00000000000000000001000001111001",
			1042 => "0000001011000000000000001100000100",
			1043 => "11111111101110110001000001111001",
			1044 => "00000000000000000001000001111001",
			1045 => "0000000001000000001001011000010000",
			1046 => "0000001110000000001010001000001100",
			1047 => "0000000101000000001101000100001000",
			1048 => "0000000101000000000011100000000100",
			1049 => "00000000000000000001000001111001",
			1050 => "00000000000110100001000001111001",
			1051 => "00000000000000000001000001111001",
			1052 => "00000000000000000001000001111001",
			1053 => "00000000000000000001000001111001",
			1054 => "0000000000000000000110011000011000",
			1055 => "0000001111000000001011000000001000",
			1056 => "0000000001000000001001111000000100",
			1057 => "00000000001010010001000010101101",
			1058 => "00000001100101000001000010101101",
			1059 => "0000001001000000000101011100000100",
			1060 => "11111110001011110001000010101101",
			1061 => "0000001111000000000010001000000100",
			1062 => "00000001100100110001000010101101",
			1063 => "0000000001000000001011101000000100",
			1064 => "11111110001111000001000010101101",
			1065 => "00000001010101000001000010101101",
			1066 => "11111110011010000001000010101101",
			1067 => "0000000000000000000110011000010100",
			1068 => "0000001100000000000100000000000100",
			1069 => "00000000000000000001000011110001",
			1070 => "0000000010000000000000110100001100",
			1071 => "0000000011000000001001010100001000",
			1072 => "0000001111000000001011011100000100",
			1073 => "00000010000001010001000011110001",
			1074 => "00000001010101110001000011110001",
			1075 => "00000100011001010001000011110001",
			1076 => "11111110011100010001000011110001",
			1077 => "0000000100000000001001100000001100",
			1078 => "0000001010000000000111101100000100",
			1079 => "11111110011011000001000011110001",
			1080 => "0000001000000000000111110100000100",
			1081 => "00000101101100010001000011110001",
			1082 => "11111111011011100001000011110001",
			1083 => "11111110011000100001000011110001",
			1084 => "0000001010000000001001111100011100",
			1085 => "0000000001000000000111100100010100",
			1086 => "0000000011000000000110100100001000",
			1087 => "0000001100000000000100000000000100",
			1088 => "11111111111101010001000100101101",
			1089 => "00000001100101110001000100101101",
			1090 => "0000000111000000001110001100001000",
			1091 => "0000000110000000001001011000000100",
			1092 => "11111101011110000001000100101101",
			1093 => "11111111000111010001000100101101",
			1094 => "00000000011101000001000100101101",
			1095 => "0000000010000000000001001000000100",
			1096 => "00000001100101000001000100101101",
			1097 => "11111111001101100001000100101101",
			1098 => "11111110011010000001000100101101",
			1099 => "0000000010000000000001101000000100",
			1100 => "00000000111111110001000101100001",
			1101 => "0000000001000000000111100100000100",
			1102 => "11111110100101000001000101100001",
			1103 => "0000000100000000001001100000010000",
			1104 => "0000000111000000000001101000001000",
			1105 => "0000001111000000000000110100000100",
			1106 => "00000000010001010001000101100001",
			1107 => "11111111100100100001000101100001",
			1108 => "0000001010000000000111101100000100",
			1109 => "00000000000000000001000101100001",
			1110 => "00000000100011000001000101100001",
			1111 => "11111111110001010001000101100001",
			1112 => "0000001010000000001001111100011000",
			1113 => "0000001111000000000000110100010100",
			1114 => "0000001100000000000100000000000100",
			1115 => "00000000000011110001000110100101",
			1116 => "0000001111000000000101110100001100",
			1117 => "0000001111000000000110110100001000",
			1118 => "0000001111000000001011011100000100",
			1119 => "00000001110100100001000110100101",
			1120 => "00000000111011100001000110100101",
			1121 => "11111111111101000001000110100101",
			1122 => "00000011010010100001000110100101",
			1123 => "11111110100100100001000110100101",
			1124 => "0000000100000000001100010100001000",
			1125 => "0000000100000000001110010000000100",
			1126 => "11111110100011100001000110100101",
			1127 => "00000000000111100001000110100101",
			1128 => "11111110011000110001000110100101",
			1129 => "0000000000000000000110011100100000",
			1130 => "0000000001000000000111100100010000",
			1131 => "0000001111000000001001001000001000",
			1132 => "0000001100000000000110000100000100",
			1133 => "00000001010011000001000111101001",
			1134 => "00000000000000000001000111101001",
			1135 => "0000000001000000000111100100000100",
			1136 => "11111110010100110001000111101001",
			1137 => "00000000000000000001000111101001",
			1138 => "0000001110000000001010001000001100",
			1139 => "0000001001000000001011001100001000",
			1140 => "0000001111000000000000110100000100",
			1141 => "00000001001010100001000111101001",
			1142 => "00000000000000000001000111101001",
			1143 => "00000010011010000001000111101001",
			1144 => "00000000000000000001000111101001",
			1145 => "11111110011101010001000111101001",
			1146 => "0000001011000000000101101100001000",
			1147 => "0000000100000000000111001000000100",
			1148 => "00000000000000000001001000101101",
			1149 => "11111111010101000001001000101101",
			1150 => "0000000010000000000001101000000100",
			1151 => "00000000011001010001001000101101",
			1152 => "0000001100000000001000000000001100",
			1153 => "0000001100000000001000111100000100",
			1154 => "00000000000000000001001000101101",
			1155 => "0000001100000000000110000100000100",
			1156 => "11111111101100010001001000101101",
			1157 => "00000000000000000001001000101101",
			1158 => "0000001100000000001000000000001000",
			1159 => "0000001011000000000101100100000100",
			1160 => "00000000000000000001001000101101",
			1161 => "00000000001010100001001000101101",
			1162 => "00000000000000000001001000101101",
			1163 => "0000000000000000000110011100100000",
			1164 => "0000000000000000000010101100001100",
			1165 => "0000001100000000000110000100000100",
			1166 => "00000001011010100001001001110001",
			1167 => "0000001100000000000110000100000100",
			1168 => "11111110111110000001001001110001",
			1169 => "00000000101111110001001001110001",
			1170 => "0000001001000000001011111100000100",
			1171 => "11111110110111110001001001110001",
			1172 => "0000001111000000001010001000001100",
			1173 => "0000001100000000001100110000000100",
			1174 => "00000000000000000001001001110001",
			1175 => "0000000111000000001101111000000100",
			1176 => "00000000000000000001001001110001",
			1177 => "00000001011110110001001001110001",
			1178 => "11111111101000000001001001110001",
			1179 => "11111110011011000001001001110001",
			1180 => "0000001010000000001001111100100100",
			1181 => "0000000100000000000110110100010100",
			1182 => "0000000111000000001001110000000100",
			1183 => "00000000010111110001001011010101",
			1184 => "0000001101000000001000011000000100",
			1185 => "00000001101010000001001011010101",
			1186 => "0000001101000000001010011100000100",
			1187 => "11111111011000100001001011010101",
			1188 => "0000001101000000001010011100000100",
			1189 => "00000000110110010001001011010101",
			1190 => "00000001101001000001001011010101",
			1191 => "0000001001000000000111101000001000",
			1192 => "0000000101000000001111011100000100",
			1193 => "11111101011001000001001011010101",
			1194 => "11111111001111000001001011010101",
			1195 => "0000001110000000000111110000000100",
			1196 => "00000001101100010001001011010101",
			1197 => "00000000000000000001001011010101",
			1198 => "0000000100000000001001100000001100",
			1199 => "0000001010000000000111101100000100",
			1200 => "11111110100100100001001011010101",
			1201 => "0000000100000000000110010000000100",
			1202 => "00000000000000000001001011010101",
			1203 => "00001101010111100001001011010101",
			1204 => "11111110011001100001001011010101",
			1205 => "0000000000000000000110011000100000",
			1206 => "0000000010000000000111010000010100",
			1207 => "0000000111000000001001110000000100",
			1208 => "00000000000111100001001100111001",
			1209 => "0000000011000000000110100100000100",
			1210 => "00000001101000000001001100111001",
			1211 => "0000001101000000001010011100000100",
			1212 => "11111110100011010001001100111001",
			1213 => "0000001101000000001010011100000100",
			1214 => "00000000011101100001001100111001",
			1215 => "00000001100110000001001100111001",
			1216 => "0000000001000000000111100100000100",
			1217 => "11111101110110110001001100111001",
			1218 => "0000001110000000000101110100000100",
			1219 => "00000001100100110001001100111001",
			1220 => "00000000010010010001001100111001",
			1221 => "0000001000000000000111110100010000",
			1222 => "0000001010000000000111101100000100",
			1223 => "11111110100111100001001100111001",
			1224 => "0000000000000000000110011100000100",
			1225 => "00000000000000000001001100111001",
			1226 => "0000001010000000000111101100000100",
			1227 => "00000110001110000001001100111001",
			1228 => "00000000000000000001001100111001",
			1229 => "11111110011001110001001100111001",
			1230 => "0000001000000000000111110100101000",
			1231 => "0000000001000000000111100100011000",
			1232 => "0000001110000000000100001000001000",
			1233 => "0000000001000000000010001100000100",
			1234 => "00000000000000000001001110001101",
			1235 => "00000000100001010001001110001101",
			1236 => "0000000001000000000110101000000100",
			1237 => "11111111000101000001001110001101",
			1238 => "0000000001000000000110101000000100",
			1239 => "00000000010001110001001110001101",
			1240 => "0000000111000000000110000100000100",
			1241 => "00000000000000000001001110001101",
			1242 => "11111111010011010001001110001101",
			1243 => "0000001110000000001010001000001100",
			1244 => "0000000101000000001110101000001000",
			1245 => "0000000010000000001110010000000100",
			1246 => "00000000101001110001001110001101",
			1247 => "00000000000000000001001110001101",
			1248 => "00000000000000000001001110001101",
			1249 => "00000000000000000001001110001101",
			1250 => "11111110110010010001001110001101",
			1251 => "0000000000000000000110011100100000",
			1252 => "0000001011000000000101100100011000",
			1253 => "0000001111000000001011000000000100",
			1254 => "00000001011000110001001111010001",
			1255 => "0000001001000000000101011100000100",
			1256 => "11111110101100110001001111010001",
			1257 => "0000001111000000000010001000000100",
			1258 => "00000001010010110001001111010001",
			1259 => "0000000110000000001011111100000100",
			1260 => "11111111011010100001001111010001",
			1261 => "0000000110000000001110010100000100",
			1262 => "00000000010111100001001111010001",
			1263 => "00000000000000000001001111010001",
			1264 => "0000001110000000001010001000000100",
			1265 => "00000010110011110001001111010001",
			1266 => "00000000000000000001001111010001",
			1267 => "11111110011100110001001111010001",
			1268 => "0000000100000000001001100000100100",
			1269 => "0000001100000000001000000000011100",
			1270 => "0000000010000000000000110100011000",
			1271 => "0000000001000000000111100100010000",
			1272 => "0000000100000000001001001000001000",
			1273 => "0000001100000000000100000000000100",
			1274 => "00000000000000000001010000011101",
			1275 => "00000001100010000001010000011101",
			1276 => "0000001001000000000000111100000100",
			1277 => "11111101110011100001010000011101",
			1278 => "11111111110111100001010000011101",
			1279 => "0000001111000000000010001000000100",
			1280 => "00000001100100000001010000011101",
			1281 => "00000000100010110001010000011101",
			1282 => "11111110110010000001010000011101",
			1283 => "0000001011000000000101100100000100",
			1284 => "00000000000000000001010000011101",
			1285 => "00000101011111010001010000011101",
			1286 => "11111110011010010001010000011101",
			1287 => "0000000100000000001001100000100100",
			1288 => "0000000100000000000111010000001000",
			1289 => "0000001100000000000100000000000100",
			1290 => "00000000000000000001010001101001",
			1291 => "00000001000001110001010001101001",
			1292 => "0000000001000000001101101000001000",
			1293 => "0000001100000000001000111100000100",
			1294 => "00000000000000000001010001101001",
			1295 => "11111111001001010001010001101001",
			1296 => "0000001110000000001010001000010000",
			1297 => "0000001100000000000110000100000100",
			1298 => "00000000000000000001010001101001",
			1299 => "0000000001000000001001011000001000",
			1300 => "0000000011000000001001100000000100",
			1301 => "00000000011100010001010001101001",
			1302 => "00000000000000000001010001101001",
			1303 => "00000000000000000001010001101001",
			1304 => "00000000000000000001010001101001",
			1305 => "11111110101011100001010001101001",
			1306 => "0000000100000000001100010100100000",
			1307 => "0000000001000000000010001100000100",
			1308 => "11111110001000100001010010101101",
			1309 => "0000000010000000000001001000010100",
			1310 => "0000000001000000000110101000010000",
			1311 => "0000001111000000000111001000001100",
			1312 => "0000001110000000000100001000000100",
			1313 => "00000001101011010001010010101101",
			1314 => "0000001110000000000001111100000100",
			1315 => "00000000000000000001010010101101",
			1316 => "00000001001010010001010010101101",
			1317 => "11111110000100010001010010101101",
			1318 => "00000001100100010001010010101101",
			1319 => "0000000111000000000110100100000100",
			1320 => "11111110100101010001010010101101",
			1321 => "00000011011100110001010010101101",
			1322 => "11111110011001100001010010101101",
			1323 => "0000001010000000000111101100101000",
			1324 => "0000000001000000000111100100010000",
			1325 => "0000001110000000000100001000001000",
			1326 => "0000000001000000000010001100000100",
			1327 => "00000000000000000001010100000001",
			1328 => "00000000001010010001010100000001",
			1329 => "0000000001000000000110101000000100",
			1330 => "11111111011000110001010100000001",
			1331 => "00000000000000000001010100000001",
			1332 => "0000000011000000001001100000010100",
			1333 => "0000001001000000001011111100000100",
			1334 => "00000000000000000001010100000001",
			1335 => "0000001100000000001100110000000100",
			1336 => "00000000000000000001010100000001",
			1337 => "0000000101000000001101000100001000",
			1338 => "0000000001000000001001011000000100",
			1339 => "00000000100110100001010100000001",
			1340 => "00000000000000000001010100000001",
			1341 => "00000000000000000001010100000001",
			1342 => "00000000000000000001010100000001",
			1343 => "11111111000100010001010100000001",
			1344 => "0000000100000000001001100000100100",
			1345 => "0000000001000000001001111000001000",
			1346 => "0000000010000000000100001000000100",
			1347 => "00000000000000000001010101001101",
			1348 => "11111110100010100001010101001101",
			1349 => "0000001011000000000100001000000100",
			1350 => "00000001010110000001010101001101",
			1351 => "0000001100000000001100110000001000",
			1352 => "0000000001000000000111100100000100",
			1353 => "11111110111100110001010101001101",
			1354 => "00000000000000000001010101001101",
			1355 => "0000000010000000001110010000001100",
			1356 => "0000000001000000000111100100000100",
			1357 => "00000000000000000001010101001101",
			1358 => "0000000110000000000000111100000100",
			1359 => "00000000000000000001010101001101",
			1360 => "00000001001001000001010101001101",
			1361 => "00000000000000000001010101001101",
			1362 => "11111110100000000001010101001101",
			1363 => "0000001000000000000111110100101000",
			1364 => "0000000001000000000111100100010000",
			1365 => "0000000000000000000010101100001100",
			1366 => "0000001100000000000100000000000100",
			1367 => "11111111100101000001010110100001",
			1368 => "0000001100000000000110000100000100",
			1369 => "00000001001110000001010110100001",
			1370 => "00000000000000000001010110100001",
			1371 => "11111110100111100001010110100001",
			1372 => "0000001110000000001010001000010100",
			1373 => "0000000110000000000000111100000100",
			1374 => "00000000000000000001010110100001",
			1375 => "0000000001000000000111100100000100",
			1376 => "00000000000000000001010110100001",
			1377 => "0000001100000000001100110000000100",
			1378 => "00000000000000000001010110100001",
			1379 => "0000000101000000001101000100000100",
			1380 => "00000001001111110001010110100001",
			1381 => "00000000000000000001010110100001",
			1382 => "00000000000000000001010110100001",
			1383 => "11111110011111010001010110100001",
			1384 => "0000000000000000000110011100100100",
			1385 => "0000001100000000000100000000000100",
			1386 => "11111111100101100001010111101101",
			1387 => "0000001111000000001010011100001100",
			1388 => "0000001001000000000000111100001000",
			1389 => "0000001001000000000000111100000100",
			1390 => "00000000011101110001010111101101",
			1391 => "00000000000000000001010111101101",
			1392 => "00000001001111000001010111101101",
			1393 => "0000001100000000001100110000000100",
			1394 => "11111111100011100001010111101101",
			1395 => "0000001110000000001010001000001100",
			1396 => "0000001001000000001110010100000100",
			1397 => "00000000000000000001010111101101",
			1398 => "0000000011000000001001100000000100",
			1399 => "00000000110100100001010111101101",
			1400 => "00000000000000000001010111101101",
			1401 => "00000000000000000001010111101101",
			1402 => "11111110100011000001010111101101",
			1403 => "0000000000000000000110011100110000",
			1404 => "0000000001000000000111100100011000",
			1405 => "0000000000000000000010101100010000",
			1406 => "0000001100000000000100000000000100",
			1407 => "11111111011010000001011001010011",
			1408 => "0000001100000000000110000100000100",
			1409 => "00000001010010110001011001010011",
			1410 => "0000001101000000001010011100000100",
			1411 => "11111111111111110001011001010011",
			1412 => "00000000000000000001011001010011",
			1413 => "0000000001000000000111100100000100",
			1414 => "11111110011101110001011001010011",
			1415 => "00000000000000000001011001010011",
			1416 => "0000001110000000001010001000010100",
			1417 => "0000000110000000000000111100000100",
			1418 => "00000000000000000001011001010011",
			1419 => "0000001100000000001100110000000100",
			1420 => "00000000000000000001011001010011",
			1421 => "0000000101000000001101000100001000",
			1422 => "0000000011000000001001100000000100",
			1423 => "00000001011100100001011001010011",
			1424 => "00000000000000000001011001010011",
			1425 => "00000000000000000001011001010011",
			1426 => "00000000000000000001011001010011",
			1427 => "11111110011110000001011001010011",
			1428 => "00000000000000000001011001010101",
			1429 => "00000000000000000001011001011001",
			1430 => "00000000000000000001011001011101",
			1431 => "00000000000000000001011001100001",
			1432 => "00000000000000000001011001100101",
			1433 => "00000000000000000001011001101001",
			1434 => "00000000000000000001011001101101",
			1435 => "00000000000000000001011001110001",
			1436 => "00000000000000000001011001110101",
			1437 => "00000000000000000001011001111001",
			1438 => "00000000000000000001011001111101",
			1439 => "00000000000000000001011010000001",
			1440 => "00000000000000000001011010000101",
			1441 => "00000000000000000001011010001001",
			1442 => "00000000000000000001011010001101",
			1443 => "00000000000000000001011010010001",
			1444 => "00000000000000000001011010010101",
			1445 => "00000000000000000001011010011001",
			1446 => "00000000000000000001011010011101",
			1447 => "00000000000000000001011010100001",
			1448 => "00000000000000000001011010100101",
			1449 => "0000000000000000000010101100000100",
			1450 => "00000000000000000001011010110001",
			1451 => "11111111111001110001011010110001",
			1452 => "0000000000000000000010101100000100",
			1453 => "00000000001010100001011010111101",
			1454 => "00000000000000000001011010111101",
			1455 => "0000001100000000001100110000000100",
			1456 => "11111111111110000001011011001001",
			1457 => "00000000000000000001011011001001",
			1458 => "0000000100000000000111001000000100",
			1459 => "00000000000000000001011011010101",
			1460 => "11111111111111000001011011010101",
			1461 => "0000001111000000001011000000000100",
			1462 => "00000000000000000001011011100001",
			1463 => "11111111111001010001011011100001",
			1464 => "0000000100000000000110110100000100",
			1465 => "00000000000011100001011011101101",
			1466 => "00000000000000000001011011101101",
			1467 => "0000000010000000001000000000000100",
			1468 => "00000000001100000001011011111001",
			1469 => "00000000000000000001011011111001",
			1470 => "0000000100000000000111010000000100",
			1471 => "00000000011001110001011100001101",
			1472 => "0000000111000000001100101000000100",
			1473 => "11111111100001110001011100001101",
			1474 => "00000000000000000001011100001101",
			1475 => "0000000100000000000111010000000100",
			1476 => "00000000101000110001011100100001",
			1477 => "0000001001000000001110010100000100",
			1478 => "11111111110011000001011100100001",
			1479 => "00000000000000000001011100100001",
			1480 => "0000001101000000001010011100000100",
			1481 => "11111111111110110001011100110101",
			1482 => "0000001101000000000010011100000100",
			1483 => "00000000000000010001011100110101",
			1484 => "00000000000000000001011100110101",
			1485 => "0000000010000000001000000000001000",
			1486 => "0000001111000000001010111100000100",
			1487 => "00000000000000000001011101001001",
			1488 => "00000000000000100001011101001001",
			1489 => "11111111111111110001011101001001",
			1490 => "0000001001000000000000111100000100",
			1491 => "11111111111100110001011101011101",
			1492 => "0000001001000000001001100100000100",
			1493 => "00000000000001100001011101011101",
			1494 => "00000000000000000001011101011101",
			1495 => "0000000010000000001000000000001000",
			1496 => "0000000001000000000110101000000100",
			1497 => "00000000000000000001011101111001",
			1498 => "00000001010000010001011101111001",
			1499 => "0000001001000000000101011100000100",
			1500 => "11111111111100100001011101111001",
			1501 => "00000000000000000001011101111001",
			1502 => "0000001001000000000000111100001000",
			1503 => "0000000100000000000111001000000100",
			1504 => "00000000000000000001011110010101",
			1505 => "11111111101001000001011110010101",
			1506 => "0000001111000000000111010000000100",
			1507 => "00000000101001100001011110010101",
			1508 => "00000000000000000001011110010101",
			1509 => "0000000010000000001000000000001000",
			1510 => "0000001100000000000100000000000100",
			1511 => "00000000000000000001011110110001",
			1512 => "00000000010111010001011110110001",
			1513 => "0000000111000000000111010000000100",
			1514 => "11111111101000000001011110110001",
			1515 => "00000000000000000001011110110001",
			1516 => "0000000100000000000111010000000100",
			1517 => "00000000011100000001011111001101",
			1518 => "0000000001000000000111100100001000",
			1519 => "0000000101000000001111011100000100",
			1520 => "11111111001111000001011111001101",
			1521 => "00000000000000000001011111001101",
			1522 => "00000000000000000001011111001101",
			1523 => "0000001001000000000101011100001100",
			1524 => "0000000010000000000100001000000100",
			1525 => "00000000000000000001011111101001",
			1526 => "0000000001000000000110101000000100",
			1527 => "11111111101000010001011111101001",
			1528 => "00000000000000000001011111101001",
			1529 => "00000000000000000001011111101001",
			1530 => "0000001001000000000000111100001100",
			1531 => "0000000100000000000111001000000100",
			1532 => "00000000000000000001100000000101",
			1533 => "0000000001000000000110101000000100",
			1534 => "11111111101100100001100000000101",
			1535 => "00000000000000000001100000000101",
			1536 => "00000000000000000001100000000101",
			1537 => "0000000100000000000111010000000100",
			1538 => "00000000000000000001100000100001",
			1539 => "0000000000000000000010101100000100",
			1540 => "00000000000000000001100000100001",
			1541 => "0000001111000000001010011100000100",
			1542 => "00000000000000000001100000100001",
			1543 => "11111111111110010001100000100001",
			1544 => "0000000000000000000010101100001000",
			1545 => "0000001100000000000110000100000100",
			1546 => "00000000110001100001100001000101",
			1547 => "00000000000000000001100001000101",
			1548 => "0000000001000000000111100100001000",
			1549 => "0000001100000000001110001100000100",
			1550 => "11111111011110010001100001000101",
			1551 => "00000000000000000001100001000101",
			1552 => "00000000000000000001100001000101",
			1553 => "0000000001000000000110101000001100",
			1554 => "0000001110000000000100001000000100",
			1555 => "00000000000000000001100001101001",
			1556 => "0000001011000000000000001100000100",
			1557 => "11111111110000110001100001101001",
			1558 => "00000000000000000001100001101001",
			1559 => "0000001110000000000110100100000100",
			1560 => "00000000000101110001100001101001",
			1561 => "00000000000000000001100001101001",
			1562 => "0000000010000000000000110100010000",
			1563 => "0000000001000000000111100100001000",
			1564 => "0000001000000000001001111100000100",
			1565 => "00000000000000000001100010001101",
			1566 => "11111111111010100001100010001101",
			1567 => "0000001110000000001101010100000100",
			1568 => "00000000000000000001100010001101",
			1569 => "00000000010101110001100010001101",
			1570 => "11111111100101010001100010001101",
			1571 => "0000001000000000000111110100010000",
			1572 => "0000001001000000001101101000000100",
			1573 => "00000000000000000001100010110001",
			1574 => "0000000011000000001001100000001000",
			1575 => "0000001001000000000000111100000100",
			1576 => "00000000000000000001100010110001",
			1577 => "00000000100101110001100010110001",
			1578 => "00000000000000000001100010110001",
			1579 => "11111111010011000001100010110001",
			1580 => "0000001001000000000000111100000100",
			1581 => "00000000000000000001100011010101",
			1582 => "0000001001000000001001100100001100",
			1583 => "0000001101000000000010011100001000",
			1584 => "0000001101000000001001110100000100",
			1585 => "00000000000000000001100011010101",
			1586 => "00000000001001110001100011010101",
			1587 => "00000000000000000001100011010101",
			1588 => "00000000000000000001100011010101",
			1589 => "0000001001000000000000111100000100",
			1590 => "11111111111011010001100011111001",
			1591 => "0000001001000000001001100100001100",
			1592 => "0000001101000000000010011100001000",
			1593 => "0000001101000000000110100100000100",
			1594 => "00000000000000000001100011111001",
			1595 => "00000000000011010001100011111001",
			1596 => "00000000000000000001100011111001",
			1597 => "00000000000000000001100011111001",
			1598 => "0000001001000000000101011100001000",
			1599 => "0000000001000000000111100100000100",
			1600 => "11111111110111010001100100100101",
			1601 => "00000000000000000001100100100101",
			1602 => "0000000001000000001001011000001100",
			1603 => "0000000101000000001110101000001000",
			1604 => "0000000111000000001101100000000100",
			1605 => "00000000000000000001100100100101",
			1606 => "00000000001001100001100100100101",
			1607 => "00000000000000000001100100100101",
			1608 => "00000000000000000001100100100101",
			1609 => "0000000001000000000110101000010000",
			1610 => "0000001111000000000001111100000100",
			1611 => "00000000000000000001100101010001",
			1612 => "0000001011000000000000001100001000",
			1613 => "0000000111000000000110000100000100",
			1614 => "11111111100010100001100101010001",
			1615 => "00000000000000000001100101010001",
			1616 => "00000000000000000001100101010001",
			1617 => "0000001111000000001011011100000100",
			1618 => "00000001000000100001100101010001",
			1619 => "00000000000000000001100101010001",
			1620 => "0000001100000000001100110000001000",
			1621 => "0000000001000000000111100100000100",
			1622 => "11111111110001000001100101111101",
			1623 => "00000000000000000001100101111101",
			1624 => "0000000001000000001001011000001100",
			1625 => "0000001100000000001000000000001000",
			1626 => "0000001001000000001101011100000100",
			1627 => "00000000000000000001100101111101",
			1628 => "00000000001111110001100101111101",
			1629 => "00000000000000000001100101111101",
			1630 => "00000000000000000001100101111101",
			1631 => "0000001001000000000000111100001100",
			1632 => "0000000010000000000100001000001000",
			1633 => "0000001000000000001000010000000100",
			1634 => "00000000011011110001100110110001",
			1635 => "00000000000000000001100110110001",
			1636 => "11111110100110110001100110110001",
			1637 => "0000000010000000000001001000001000",
			1638 => "0000001001000000000101011100000100",
			1639 => "00000000000000000001100110110001",
			1640 => "00000000110110010001100110110001",
			1641 => "0000000111000000000111010000000100",
			1642 => "11111111010001110001100110110001",
			1643 => "00000000000000000001100110110001",
			1644 => "0000001001000000000101011100001100",
			1645 => "0000001110000000000100001000000100",
			1646 => "00000000000000000001100111100101",
			1647 => "0000000001000000000111100100000100",
			1648 => "11111111101111110001100111100101",
			1649 => "00000000000000000001100111100101",
			1650 => "0000000001000000001001011000001100",
			1651 => "0000001110000000001010001000001000",
			1652 => "0000000111000000001101100000000100",
			1653 => "00000000000000000001100111100101",
			1654 => "00000000001101110001100111100101",
			1655 => "00000000000000000001100111100101",
			1656 => "00000000000000000001100111100101",
			1657 => "0000001100000000001100110000001100",
			1658 => "0000001111000000000001111100000100",
			1659 => "00000000000000000001101000011001",
			1660 => "0000000001000000000111100100000100",
			1661 => "11111111100110100001101000011001",
			1662 => "00000000000000000001101000011001",
			1663 => "0000000001000000000110101000000100",
			1664 => "00000000000000000001101000011001",
			1665 => "0000000010000000001110010000001000",
			1666 => "0000000001000000001001011000000100",
			1667 => "00000000100100110001101000011001",
			1668 => "00000000000000000001101000011001",
			1669 => "00000000000000000001101000011001",
			1670 => "0000000000000000000110011000010000",
			1671 => "0000001100000000000100000000000100",
			1672 => "00000000000000000001101001010101",
			1673 => "0000001111000000000000110100001000",
			1674 => "0000000010000000000101110100000100",
			1675 => "00000010001000000001101001010101",
			1676 => "00000110010110000001101001010101",
			1677 => "11111110011010010001101001010101",
			1678 => "0000000100000000001001100000001100",
			1679 => "0000001000000000000111110100000100",
			1680 => "11111110011010100001101001010101",
			1681 => "0000001000000000000111110100000100",
			1682 => "00001011100111010001101001010101",
			1683 => "11111111001010000001101001010101",
			1684 => "11111110011000010001101001010101",
			1685 => "0000000100000000001001100000011000",
			1686 => "0000001001000000000000111100001100",
			1687 => "0000001111000000001011000000001000",
			1688 => "0000000111000000001001110000000100",
			1689 => "00000000000000000001101010001001",
			1690 => "00000000100010010001101010001001",
			1691 => "11111111101011100001101010001001",
			1692 => "0000000111000000000110000100000100",
			1693 => "00000000000000000001101010001001",
			1694 => "0000001110000000001010001000000100",
			1695 => "00000000111100100001101010001001",
			1696 => "00000000000000000001101010001001",
			1697 => "11111111001110000001101010001001",
			1698 => "0000000001000000000111100100001000",
			1699 => "0000001000000000001001111100000100",
			1700 => "00000000000000000001101010111101",
			1701 => "11111111000111100001101010111101",
			1702 => "0000000010000000001110010000010000",
			1703 => "0000000110000000000000111100000100",
			1704 => "00000000000000000001101010111101",
			1705 => "0000000001000000001001011000001000",
			1706 => "0000000101000000001110101000000100",
			1707 => "00000000100001110001101010111101",
			1708 => "00000000000000000001101010111101",
			1709 => "00000000000000000001101010111101",
			1710 => "00000000000000000001101010111101",
			1711 => "0000001001000000000000111100001000",
			1712 => "0000000111000000001110001100000100",
			1713 => "11111111111001010001101011110001",
			1714 => "00000000000000000001101011110001",
			1715 => "0000001001000000001001100100010000",
			1716 => "0000000101000000001110101000001100",
			1717 => "0000000111000000001101100000000100",
			1718 => "00000000000000000001101011110001",
			1719 => "0000001100000000001000000000000100",
			1720 => "00000000001011000001101011110001",
			1721 => "00000000000000000001101011110001",
			1722 => "00000000000000000001101011110001",
			1723 => "00000000000000000001101011110001",
			1724 => "0000000000000000000010101100000100",
			1725 => "00000000011111110001101100011101",
			1726 => "0000000001000000000111100100000100",
			1727 => "11111111010101000001101100011101",
			1728 => "0000000010000000001110010000001100",
			1729 => "0000000110000000001101111100001000",
			1730 => "0000000101000000001101000100000100",
			1731 => "00000000010000000001101100011101",
			1732 => "00000000000000000001101100011101",
			1733 => "00000000000000000001101100011101",
			1734 => "00000000000000000001101100011101",
			1735 => "0000000000000000000110011000010100",
			1736 => "0000000100000000000110110100001100",
			1737 => "0000000100000000001001001000000100",
			1738 => "00000001101001000001101101100001",
			1739 => "0000001001000000000101011100000100",
			1740 => "11111110111011010001101101100001",
			1741 => "00000001101000010001101101100001",
			1742 => "0000001001000000000111101000000100",
			1743 => "11111110000000010001101101100001",
			1744 => "00000001011111110001101101100001",
			1745 => "0000000100000000001001100000001100",
			1746 => "0000001010000000000111101100000100",
			1747 => "11111110100110100001101101100001",
			1748 => "0000000100000000000110010000000100",
			1749 => "00000000000000000001101101100001",
			1750 => "00001000001010100001101101100001",
			1751 => "11111110011001110001101101100001",
			1752 => "0000001001000000000000111100001100",
			1753 => "0000000001000000000110101000001000",
			1754 => "0000000111000000001110001100000100",
			1755 => "11111111110110000001101110011101",
			1756 => "00000000000000000001101110011101",
			1757 => "00000000000000000001101110011101",
			1758 => "0000000001000000001001011000010000",
			1759 => "0000000101000000001110101000001100",
			1760 => "0000000111000000001101100000000100",
			1761 => "00000000000000000001101110011101",
			1762 => "0000001100000000001000000000000100",
			1763 => "00000000001100110001101110011101",
			1764 => "00000000000000000001101110011101",
			1765 => "00000000000000000001101110011101",
			1766 => "00000000000000000001101110011101",
			1767 => "0000001001000000000000111100010100",
			1768 => "0000000100000000001001001000001100",
			1769 => "0000000100000000000111001000000100",
			1770 => "00000000010110010001101111101001",
			1771 => "0000000110000000001101011100000100",
			1772 => "11111111100100100001101111101001",
			1773 => "00000000000000000001101111101001",
			1774 => "0000000001000000000110101000000100",
			1775 => "11111110100100100001101111101001",
			1776 => "00000000000000000001101111101001",
			1777 => "0000001110000000000111110000001100",
			1778 => "0000001001000000000101011100000100",
			1779 => "00000000000000000001101111101001",
			1780 => "0000000000000000000110011100000100",
			1781 => "00000000110001110001101111101001",
			1782 => "00000000000000000001101111101001",
			1783 => "0000000111000000000111010000000100",
			1784 => "11111111011010100001101111101001",
			1785 => "00000000000000000001101111101001",
			1786 => "0000000010000000000001001000011000",
			1787 => "0000000100000000001001001000000100",
			1788 => "00000000101101000001110000100101",
			1789 => "0000001001000000000000111100001000",
			1790 => "0000000110000000001001011000000100",
			1791 => "11111111000011100001110000100101",
			1792 => "00000000000000000001110000100101",
			1793 => "0000001111000000001010011100000100",
			1794 => "00000000101110100001110000100101",
			1795 => "0000001100000000000110000100000100",
			1796 => "11111111100111000001110000100101",
			1797 => "00000000000100100001110000100101",
			1798 => "0000000111000000000111010000000100",
			1799 => "11111110110100110001110000100101",
			1800 => "00000000000000000001110000100101",
			1801 => "0000000010000000000001001000011100",
			1802 => "0000001001000000000101011100010100",
			1803 => "0000001111000000000001111100001000",
			1804 => "0000000001000000000010001100000100",
			1805 => "00000000000000000001110001101001",
			1806 => "00000000100010000001110001101001",
			1807 => "0000001001000000000000111100001000",
			1808 => "0000000111000000001101100000000100",
			1809 => "00000000000000000001110001101001",
			1810 => "11111111000001110001110001101001",
			1811 => "00000000000000000001110001101001",
			1812 => "0000001111000000000010001000000100",
			1813 => "00000000110110110001110001101001",
			1814 => "00000000000000000001110001101001",
			1815 => "0000000111000000000111010000000100",
			1816 => "11111110101101110001110001101001",
			1817 => "00000000000000000001110001101001",
			1818 => "0000000100000000001100010100011100",
			1819 => "0000000001000000000111100100001100",
			1820 => "0000000100000000001001001000001000",
			1821 => "0000000110000000001111001100000100",
			1822 => "00000000000000000001110010100101",
			1823 => "00000001010111000001110010100101",
			1824 => "11111110111011010001110010100101",
			1825 => "0000001111000000000010001000000100",
			1826 => "00000001011010100001110010100101",
			1827 => "0000000011000000000001001000000100",
			1828 => "11111111100011010001110010100101",
			1829 => "0000001111000000001010001000000100",
			1830 => "00000000100101100001110010100101",
			1831 => "00000000000000000001110010100101",
			1832 => "11111110011011110001110010100101",
			1833 => "0000000001000000000111100100011000",
			1834 => "0000001111000000001011000000001100",
			1835 => "0000001100000000000100000000000100",
			1836 => "00000000000000000001110011111001",
			1837 => "0000000110000000000111101000000100",
			1838 => "00000000001011000001110011111001",
			1839 => "00000000000000000001110011111001",
			1840 => "0000001100000000001110001100001000",
			1841 => "0000000110000000001001011000000100",
			1842 => "00000000000000000001110011111001",
			1843 => "11111111000010000001110011111001",
			1844 => "00000000000000000001110011111001",
			1845 => "0000000010000000001110010000010000",
			1846 => "0000000110000000000000111100000100",
			1847 => "00000000000000000001110011111001",
			1848 => "0000000001000000001001011000001000",
			1849 => "0000001110000000001010001000000100",
			1850 => "00000000101010010001110011111001",
			1851 => "00000000000000000001110011111001",
			1852 => "00000000000000000001110011111001",
			1853 => "00000000000000000001110011111001",
			1854 => "0000000100000000001100010100100000",
			1855 => "0000000001000000000111100100010000",
			1856 => "0000000100000000001001001000001000",
			1857 => "0000000110000000001111001100000100",
			1858 => "00000000000000000001110100111101",
			1859 => "00000001010101010001110100111101",
			1860 => "0000000001000000000110101000000100",
			1861 => "11111110101000010001110100111101",
			1862 => "11111111110101010001110100111101",
			1863 => "0000001111000000000010001000000100",
			1864 => "00000001011001000001110100111101",
			1865 => "0000001101000000000101110100000100",
			1866 => "11111111101110110001110100111101",
			1867 => "0000001111000000001010001000000100",
			1868 => "00000000101000010001110100111101",
			1869 => "00000000000000000001110100111101",
			1870 => "11111110011100010001110100111101",
			1871 => "0000000000000000000110011100100000",
			1872 => "0000000001000000000111100100010000",
			1873 => "0000001111000000001001001000001000",
			1874 => "0000001100000000000110000100000100",
			1875 => "00000001001111000001110110000001",
			1876 => "00000000000000000001110110000001",
			1877 => "0000000001000000000111100100000100",
			1878 => "11111110011101000001110110000001",
			1879 => "00000000000000000001110110000001",
			1880 => "0000000011000000001001100000001100",
			1881 => "0000000110000000000000111100000100",
			1882 => "00000000000000000001110110000001",
			1883 => "0000000010000000001110010000000100",
			1884 => "00000001011111100001110110000001",
			1885 => "00000000000000000001110110000001",
			1886 => "00000000000000000001110110000001",
			1887 => "11111110011101110001110110000001",
			1888 => "0000000000000000000010101100000100",
			1889 => "00000000100001100001110110110101",
			1890 => "0000000001000000000111100100000100",
			1891 => "11111111010010100001110110110101",
			1892 => "0000000110000000001101111100010000",
			1893 => "0000001110000000001010001000001100",
			1894 => "0000000101000000001101000100001000",
			1895 => "0000001100000000001100110000000100",
			1896 => "00000000000000000001110110110101",
			1897 => "00000000010100010001110110110101",
			1898 => "00000000000000000001110110110101",
			1899 => "00000000000000000001110110110101",
			1900 => "00000000000000000001110110110101",
			1901 => "0000000000000000000110011000011100",
			1902 => "0000001111000000000000110100011000",
			1903 => "0000001111000000000101110100010100",
			1904 => "0000000100000000000110110100001100",
			1905 => "0000001111000000000111010000000100",
			1906 => "00000001111011010001111000000001",
			1907 => "0000001110000000001010001100000100",
			1908 => "00000000011001010001111000000001",
			1909 => "00000001110100100001111000000001",
			1910 => "0000000110000000000101011100000100",
			1911 => "11111101111011000001111000000001",
			1912 => "00000001111010110001111000000001",
			1913 => "00000011110110000001111000000001",
			1914 => "11111110100001000001111000000001",
			1915 => "0000000100000000001100010100001000",
			1916 => "0000000100000000001110010000000100",
			1917 => "11111110100001110001111000000001",
			1918 => "00000000000000010001111000000001",
			1919 => "11111110011000100001111000000001",
			1920 => "0000000000000000000110011000011000",
			1921 => "0000001001000000000100110100010100",
			1922 => "0000001111000000000001001000010000",
			1923 => "0000001100000000000100000000000100",
			1924 => "00000000000110010001111001010101",
			1925 => "0000001111000000000110110100001000",
			1926 => "0000001111000000001011011100000100",
			1927 => "00000010010011100001111001010101",
			1928 => "00000001100110110001111001010101",
			1929 => "00000011001000000001111001010101",
			1930 => "11111110010110110001111001010101",
			1931 => "00000101110010110001111001010101",
			1932 => "0000000000000000000110011100010000",
			1933 => "0000001000000000000111110100000100",
			1934 => "11111110011001110001111001010101",
			1935 => "0000001000000000000111110100001000",
			1936 => "0000001010000000000111101100000100",
			1937 => "11111111011000000001111001010101",
			1938 => "00000011011001000001111001010101",
			1939 => "11111111001000110001111001010101",
			1940 => "11111110011000000001111001010101",
			1941 => "0000000000000000000110011000100000",
			1942 => "0000000001000000001001111000000100",
			1943 => "11111111000010010001111010110001",
			1944 => "0000001111000000000010001000010100",
			1945 => "0000000001000000001001111000001000",
			1946 => "0000001110000000001100110000000100",
			1947 => "00000001101011110001111010110001",
			1948 => "11111111110001100001111010110001",
			1949 => "0000001110000000001011000000000100",
			1950 => "00000001110000000001111010110001",
			1951 => "0000001100000000001100110000000100",
			1952 => "11111111111110000001111010110001",
			1953 => "00000001110000000001111010110001",
			1954 => "0000000111000000000100001000000100",
			1955 => "11111101100001100001111010110001",
			1956 => "00000010000111010001111010110001",
			1957 => "0000000000000000000110011100001100",
			1958 => "0000001000000000000111110100000100",
			1959 => "11111110011101110001111010110001",
			1960 => "0000001000000000000111110100000100",
			1961 => "00000010110000010001111010110001",
			1962 => "11111111101101110001111010110001",
			1963 => "11111110011001010001111010110001",
			1964 => "0000001000000000000111110100101000",
			1965 => "0000000001000000000111100100010100",
			1966 => "0000001000000000000101010000001100",
			1967 => "0000001110000000000100001000000100",
			1968 => "00000000011101000001111100000101",
			1969 => "0000001111000000001101010100000100",
			1970 => "11111111101100010001111100000101",
			1971 => "00000000000000000001111100000101",
			1972 => "0000001001000000000000111100000100",
			1973 => "11111111001100000001111100000101",
			1974 => "00000000000000000001111100000101",
			1975 => "0000001110000000001010001000010000",
			1976 => "0000000101000000001110101000001100",
			1977 => "0000000011000000001001100000001000",
			1978 => "0000000010000000001110010000000100",
			1979 => "00000000100011110001111100000101",
			1980 => "00000000000000000001111100000101",
			1981 => "00000000000000000001111100000101",
			1982 => "00000000000000000001111100000101",
			1983 => "00000000000000000001111100000101",
			1984 => "11111110110110010001111100000101",
			1985 => "0000001000000000000111110100100000",
			1986 => "0000000001000000001001111000001000",
			1987 => "0000000010000000000100001000000100",
			1988 => "00000000000000000001111101001001",
			1989 => "11111111000001100001111101001001",
			1990 => "0000001111000000001010011100000100",
			1991 => "00000000111010010001111101001001",
			1992 => "0000000001000000000111100100000100",
			1993 => "11111111010101000001111101001001",
			1994 => "0000001110000000001010001000001100",
			1995 => "0000000110000000000101011100000100",
			1996 => "00000000000000000001111101001001",
			1997 => "0000000101000000001110101000000100",
			1998 => "00000000101100000001111101001001",
			1999 => "00000000000000000001111101001001",
			2000 => "00000000000000000001111101001001",
			2001 => "11111110100101000001111101001001",
			2002 => "0000000100000000001001100000100100",
			2003 => "0000001100000000001000000000011100",
			2004 => "0000000010000000000000110100011000",
			2005 => "0000000001000000000111100100010000",
			2006 => "0000000100000000001001001000001000",
			2007 => "0000001100000000000100000000000100",
			2008 => "00000000000000000001111110010101",
			2009 => "00000001100001000001111110010101",
			2010 => "0000001001000000000000111100000100",
			2011 => "11111101111110110001111110010101",
			2012 => "11111111111101010001111110010101",
			2013 => "0000001111000000000010001000000100",
			2014 => "00000001100011000001111110010101",
			2015 => "00000000011111010001111110010101",
			2016 => "11111110110110000001111110010101",
			2017 => "0000001011000000000101100100000100",
			2018 => "00000000000000000001111110010101",
			2019 => "00000011101011100001111110010101",
			2020 => "11111110011010100001111110010101",
			2021 => "0000001010000000001001111100011100",
			2022 => "0000000001000000001001111000000100",
			2023 => "11111110111010100001111111110001",
			2024 => "0000000010000000000000110100010100",
			2025 => "0000001111000000001011000000000100",
			2026 => "00000001110011000001111111110001",
			2027 => "0000000001000000000111100100000100",
			2028 => "11111101011001100001111111110001",
			2029 => "0000000111000000000110000100001000",
			2030 => "0000000110000000000000111100000100",
			2031 => "00000001101101000001111111110001",
			2032 => "11111111011100100001111111110001",
			2033 => "00000001110101110001111111110001",
			2034 => "11111110101110000001111111110001",
			2035 => "0000000100000000001001100000010000",
			2036 => "0000001010000000000111101100000100",
			2037 => "11111110011101100001111111110001",
			2038 => "0000001010000000000111101100001000",
			2039 => "0000001000000000000111110100000100",
			2040 => "00000000000000000001111111110001",
			2041 => "00001000000100110001111111110001",
			2042 => "11111111101010010001111111110001",
			2043 => "11111110011001000001111111110001",
			2044 => "0000001000000000000111110100100000",
			2045 => "0000000010000000000001101000000100",
			2046 => "00000000111100100010000000110101",
			2047 => "0000000001000000001101101000001000",
			2048 => "0000001100000000001000111100000100",
			2049 => "00000000000000000010000000110101",
			2050 => "11111111000101000010000000110101",
			2051 => "0000001110000000001010001000010000",
			2052 => "0000001100000000000110000100000100",
			2053 => "00000000000000000010000000110101",
			2054 => "0000000101000000001110101000001000",
			2055 => "0000000010000000001110010000000100",
			2056 => "00000000011111010010000000110101",
			2057 => "00000000000000000010000000110101",
			2058 => "00000000000000000010000000110101",
			2059 => "00000000000000000010000000110101",
			2060 => "11111110101010000010000000110101",
			2061 => "0000000001000000000110101000010000",
			2062 => "0000000010000000000100001000000100",
			2063 => "00000000000010110010000010011001",
			2064 => "0000000111000000000110000100001000",
			2065 => "0000001011000000000000001100000100",
			2066 => "11111110110110010010000010011001",
			2067 => "00000000000000000010000010011001",
			2068 => "00000000000000000010000010011001",
			2069 => "0000000000000000000010101100000100",
			2070 => "00000000100001000010000010011001",
			2071 => "0000000001000000000111100100001100",
			2072 => "0000001110000000000110100100000100",
			2073 => "00000000000000000010000010011001",
			2074 => "0000000111000000000101101100000100",
			2075 => "00000000000000000010000010011001",
			2076 => "11111111100000010010000010011001",
			2077 => "0000000010000000001110010000010000",
			2078 => "0000001100000000001100110000000100",
			2079 => "00000000000000000010000010011001",
			2080 => "0000001001000000001110010100000100",
			2081 => "00000000000000000010000010011001",
			2082 => "0000000001000000001001011000000100",
			2083 => "00000000101001110010000010011001",
			2084 => "00000000000000000010000010011001",
			2085 => "00000000000000000010000010011001",
			2086 => "0000000100000000001001100000100100",
			2087 => "0000000001000000001001111000001000",
			2088 => "0000000010000000000100001000000100",
			2089 => "00000000000000000010000011100101",
			2090 => "11111110100111110010000011100101",
			2091 => "0000001011000000000100001000000100",
			2092 => "00000001010011110010000011100101",
			2093 => "0000001100000000001100110000001000",
			2094 => "0000000001000000000111100100000100",
			2095 => "11111111000011110010000011100101",
			2096 => "00000000000000000010000011100101",
			2097 => "0000001110000000001010001000001100",
			2098 => "0000000001000000000111100100000100",
			2099 => "00000000000000000010000011100101",
			2100 => "0000000110000000000000111100000100",
			2101 => "00000000000000000010000011100101",
			2102 => "00000001000100100010000011100101",
			2103 => "00000000000000000010000011100101",
			2104 => "11111110100000110010000011100101",
			2105 => "0000001000000000000111110100101000",
			2106 => "0000000001000000001001111000001000",
			2107 => "0000001111000000000001111100000100",
			2108 => "00000000000000000010000100111001",
			2109 => "11111111000101000010000100111001",
			2110 => "0000001111000000001010011100001100",
			2111 => "0000001011000000000100001000000100",
			2112 => "00000001000101110010000100111001",
			2113 => "0000001011000000000001111100000100",
			2114 => "00000000000000000010000100111001",
			2115 => "00000000010110100010000100111001",
			2116 => "0000000001000000000111100100000100",
			2117 => "11111111011000010010000100111001",
			2118 => "0000001110000000001010001000001100",
			2119 => "0000000110000000000101011100000100",
			2120 => "00000000000000000010000100111001",
			2121 => "0000000101000000001110101000000100",
			2122 => "00000000100111110010000100111001",
			2123 => "00000000000000000010000100111001",
			2124 => "00000000000000000010000100111001",
			2125 => "11111110100110010010000100111001",
			2126 => "0000001000000000000111110100101000",
			2127 => "0000001100000000001000000000100000",
			2128 => "0000000010000000000000110100011100",
			2129 => "0000000001000000000111100100010000",
			2130 => "0000001000000000000101010000001000",
			2131 => "0000001100000000000100000000000100",
			2132 => "00000000000000000010000110001101",
			2133 => "00000001100011010010000110001101",
			2134 => "0000000000000000001010100000000100",
			2135 => "00000000011111100010000110001101",
			2136 => "11111110000011110010000110001101",
			2137 => "0000000111000000000110000100001000",
			2138 => "0000001111000000000110100100000100",
			2139 => "00000001010100000010000110001101",
			2140 => "00000000000000000010000110001101",
			2141 => "00000001100110010010000110001101",
			2142 => "11111110101101110010000110001101",
			2143 => "0000000011000000001001100000000100",
			2144 => "00001011001000000010000110001101",
			2145 => "00000000000000000010000110001101",
			2146 => "11111110011010010010000110001101",
			2147 => "0000000100000000001100010100100100",
			2148 => "0000001001000000001101101000000100",
			2149 => "11111111000010100010000111011011",
			2150 => "0000001111000000001011000000000100",
			2151 => "00000001100010010010000111011011",
			2152 => "0000000111000000000110000100001100",
			2153 => "0000001001000000000101011100000100",
			2154 => "11111110101111110010000111011011",
			2155 => "0000001100000000001100110000000100",
			2156 => "00000000001101110010000111011011",
			2157 => "11111111110000000010000111011011",
			2158 => "0000001111000000000000110100000100",
			2159 => "00000001010101000010000111011011",
			2160 => "0000000010000000000111111100000100",
			2161 => "11111111001111110010000111011011",
			2162 => "0000000010000000001001011100000100",
			2163 => "00000001100101010010000111011011",
			2164 => "00000000000000000010000111011011",
			2165 => "11111110011010110010000111011011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(710, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(1428, initial_addr_3'length));
	end generate gen_rom_3;

	gen_rom_4: if SELECT_ROM = 4 generate
		bank <= (
			0 => "00000000000000000000000000000101",
			1 => "00000000000000000000000000001001",
			2 => "00000000000000000000000000001101",
			3 => "00000000000000000000000000010001",
			4 => "00000000000000000000000000010101",
			5 => "00000000000000000000000000011001",
			6 => "00000000000000000000000000011101",
			7 => "00000000000000000000000000100001",
			8 => "00000000000000000000000000100101",
			9 => "0000001011000000000100010000001000",
			10 => "0000001011000000001011011100000100",
			11 => "00000000000000000000000001000001",
			12 => "00000000001000100000000001000001",
			13 => "0000001011000000000111111100000100",
			14 => "11111111111000000000000001000001",
			15 => "00000000000000000000000001000001",
			16 => "0000001010000000000000001000001000",
			17 => "0000001010000000001011001100000100",
			18 => "00000000000000000000000001011101",
			19 => "00000000001000100000000001011101",
			20 => "0000001010000000000110011000000100",
			21 => "11111111111101110000000001011101",
			22 => "00000000000000000000000001011101",
			23 => "0000000001000000000110101000000100",
			24 => "00000000000000000000000001111001",
			25 => "0000001101000000001010001000001000",
			26 => "0000000111000000001111011100000100",
			27 => "11111111110110010000000001111001",
			28 => "00000000000000000000000001111001",
			29 => "00000000000000000000000001111001",
			30 => "0000000101000000001111010000001100",
			31 => "0000000111000000000001101000000100",
			32 => "00000000000000000000000010011101",
			33 => "0000000101000000001101000100000100",
			34 => "00000000000000000000000010011101",
			35 => "11111111110010100000000010011101",
			36 => "0000000111000000000001001000000100",
			37 => "00000000001011000000000010011101",
			38 => "00000000000000000000000010011101",
			39 => "0000001001000000000101011100001100",
			40 => "0000001110000000000100001000000100",
			41 => "00000000000000000000000011000001",
			42 => "0000000000000000001100011100000100",
			43 => "00000000000100000000000011000001",
			44 => "00000000000000000000000011000001",
			45 => "0000000110000000001101111100000100",
			46 => "11111111101011110000000011000001",
			47 => "00000000000000000000000011000001",
			48 => "0000000111000000001000011000001000",
			49 => "0000000111000000000001101000000100",
			50 => "00000000000000000000000011100101",
			51 => "11111111111000000000000011100101",
			52 => "0000000011000000001010000100000100",
			53 => "00000000000000000000000011100101",
			54 => "0000000011000000000010100100000100",
			55 => "00000000000001110000000011100101",
			56 => "00000000000000000000000011100101",
			57 => "0000001011000000000101100100001100",
			58 => "0000001100000000001100110000000100",
			59 => "00000000000000000000000100010001",
			60 => "0000001100000000001000000000000100",
			61 => "11111111111010110000000100010001",
			62 => "00000000000000000000000100010001",
			63 => "0000000001000000000000111100001000",
			64 => "0000000111000000000111010000000100",
			65 => "00000000001100010000000100010001",
			66 => "00000000000000000000000100010001",
			67 => "00000000000000000000000100010001",
			68 => "0000001010000000000000001000001100",
			69 => "0000000000000000000010101100000100",
			70 => "00000000000000000000000100111101",
			71 => "0000000000000000000001110000000100",
			72 => "00000000001010110000000100111101",
			73 => "00000000000000000000000100111101",
			74 => "0000001010000000000110011000001000",
			75 => "0000000000000000000001010100000100",
			76 => "00000000000000000000000100111101",
			77 => "11111111111101100000000100111101",
			78 => "00000000000000000000000100111101",
			79 => "0000001011000000000100010000010000",
			80 => "0000001011000000001000011000000100",
			81 => "00000000000000000000000101100001",
			82 => "0000000001000000000000111100001000",
			83 => "0000000001000000001111001100000100",
			84 => "00000000000000000000000101100001",
			85 => "00000000001100010000000101100001",
			86 => "00000000000000000000000101100001",
			87 => "00000000000000000000000101100001",
			88 => "0000000100000000001111100100010000",
			89 => "0000000010000000001100010000000100",
			90 => "00000000000000000000000110000101",
			91 => "0000000010000000001010000100001000",
			92 => "0000001000000000001001000100000100",
			93 => "00000000001100100000000110000101",
			94 => "00000000000000000000000110000101",
			95 => "00000000000000000000000110000101",
			96 => "00000000000000000000000110000101",
			97 => "0000001100000000001100110000000100",
			98 => "00000000000000000000000110101001",
			99 => "0000000101000000001111010000001100",
			100 => "0000001101000000001010001000001000",
			101 => "0000000111000000001111011100000100",
			102 => "11111111101111010000000110101001",
			103 => "00000000000000000000000110101001",
			104 => "00000000000000000000000110101001",
			105 => "00000000000000000000000110101001",
			106 => "0000000101000000001110010000010000",
			107 => "0000000000000000001100011100001000",
			108 => "0000001010000000000100111100000100",
			109 => "11111111111101010000000111011101",
			110 => "00000000000000010000000111011101",
			111 => "0000001010000000000111101100000100",
			112 => "00000000000000000000000111011101",
			113 => "11111111101111110000000111011101",
			114 => "0000000110000000001000010000001000",
			115 => "0000000001000000001101111100000100",
			116 => "00000000000100100000000111011101",
			117 => "00000000000000000000000111011101",
			118 => "00000000000000000000000111011101",
			119 => "0000000111000000001000011000010000",
			120 => "0000001111000000001011000000000100",
			121 => "00000000000000000000001000010001",
			122 => "0000001111000000001010000100001000",
			123 => "0000001011000000000100010000000100",
			124 => "11111111110100110000001000010001",
			125 => "00000000000000000000001000010001",
			126 => "00000000000000000000001000010001",
			127 => "0000001111000000000110111100001000",
			128 => "0000001111000000000010000100000100",
			129 => "00000000000000000000001000010001",
			130 => "00000000001000100000001000010001",
			131 => "00000000000000000000001000010001",
			132 => "0000001010000000000000001000010000",
			133 => "0000001010000000000100110100000100",
			134 => "00000000000000000000001001000101",
			135 => "0000000000000000000001010100001000",
			136 => "0000001010000000000111101100000100",
			137 => "00000000000100000000001001000101",
			138 => "00000000000000000000001001000101",
			139 => "00000000000000000000001001000101",
			140 => "0000000000000000000101000100000100",
			141 => "00000000000000000000001001000101",
			142 => "0000001010000000000110011000000100",
			143 => "11111111111101000000001001000101",
			144 => "00000000000000000000001001000101",
			145 => "0000000011000000001110110100001100",
			146 => "0000001001000000000000111100000100",
			147 => "00000000000000000000001001111001",
			148 => "0000000001000000000110101000000100",
			149 => "00000000000000000000001001111001",
			150 => "11111111111010100000001001111001",
			151 => "0000000010000000000111010100001100",
			152 => "0000001011000000000101110100001000",
			153 => "0000000001000000000000111100000100",
			154 => "00000000001111110000001001111001",
			155 => "00000000000000000000001001111001",
			156 => "00000000000000000000001001111001",
			157 => "00000000000000000000001001111001",
			158 => "0000001010000000000000001000001100",
			159 => "0000001110000000000100001000000100",
			160 => "00000000000000000000001010110101",
			161 => "0000000111000000001101100000000100",
			162 => "00000000000000000000001010110101",
			163 => "00000000000111010000001010110101",
			164 => "0000000011000000001010000100001000",
			165 => "0000000101000000001111010000000100",
			166 => "11111111111011100000001010110101",
			167 => "00000000000000000000001010110101",
			168 => "0000000101000000001110000100000100",
			169 => "00000000000000000000001010110101",
			170 => "0000000101000000001000100000000100",
			171 => "00000000000010100000001010110101",
			172 => "00000000000000000000001010110101",
			173 => "0000000100000000001111100100010100",
			174 => "0000000010000000001100010000000100",
			175 => "00000000000000000000001011101001",
			176 => "0000001011000000000101110100001100",
			177 => "0000001001000000001000010000001000",
			178 => "0000000001000000000000111100000100",
			179 => "00000000011010000000001011101001",
			180 => "00000000000000000000001011101001",
			181 => "00000000000000000000001011101001",
			182 => "00000000000000000000001011101001",
			183 => "0000001011000000000111111100000100",
			184 => "11111111111110000000001011101001",
			185 => "00000000000000000000001011101001",
			186 => "0000001100000000001100110000000100",
			187 => "00000000000000000000001100010101",
			188 => "0000000101000000001111010000010000",
			189 => "0000001101000000001010001000001100",
			190 => "0000001100000000001001110100001000",
			191 => "0000000010000000000110101100000100",
			192 => "11111111101101100000001100010101",
			193 => "00000000000000000000001100010101",
			194 => "00000000000000000000001100010101",
			195 => "00000000000000000000001100010101",
			196 => "00000000000000000000001100010101",
			197 => "0000001000000000001001101000010100",
			198 => "0000001110000000000100001000000100",
			199 => "00000000000000000000001101000001",
			200 => "0000000001000000001001011000001100",
			201 => "0000001010000000001010100100001000",
			202 => "0000000111000000001101100000000100",
			203 => "00000000000000000000001101000001",
			204 => "00000000000111110000001101000001",
			205 => "00000000000000000000001101000001",
			206 => "00000000000000000000001101000001",
			207 => "00000000000000000000001101000001",
			208 => "0000001110000000000110100100000100",
			209 => "11111111011011100000001101110101",
			210 => "0000000101000000000101001000001000",
			211 => "0000001100000000001011000000000100",
			212 => "00000000000000000000001101110101",
			213 => "11111111101101100000001101110101",
			214 => "0000001100000000001011011100001100",
			215 => "0000000101000000001111010000000100",
			216 => "00000000000000000000001101110101",
			217 => "0000001100000000001011000000000100",
			218 => "00000000000000000000001101110101",
			219 => "00000000000100010000001101110101",
			220 => "00000000000000000000001101110101",
			221 => "0000000111000000000110000100010000",
			222 => "0000001100000000000100000000000100",
			223 => "00000000000000000000001110111001",
			224 => "0000001100000000000110000100001000",
			225 => "0000000001000000001101101000000100",
			226 => "11111111111010100000001110111001",
			227 => "00000000000000000000001110111001",
			228 => "00000000000000000000001110111001",
			229 => "0000000001000000000000111100010000",
			230 => "0000000111000000001111011100001100",
			231 => "0000001100000000000011011100000100",
			232 => "00000000000000000000001110111001",
			233 => "0000000001000000000110101000000100",
			234 => "00000000000000000000001110111001",
			235 => "00000000001001100000001110111001",
			236 => "00000000000000000000001110111001",
			237 => "00000000000000000000001110111001",
			238 => "0000000011000000001100010000010000",
			239 => "0000001111000000001011000000000100",
			240 => "00000000000000000000010000000101",
			241 => "0000001101000000000010011100001000",
			242 => "0000001100000000001000000000000100",
			243 => "11111111101111110000010000000101",
			244 => "00000000000000000000010000000101",
			245 => "00000000000000000000010000000101",
			246 => "0000001111000000001100000000001000",
			247 => "0000000110000000000100110100000100",
			248 => "00000000010011000000010000000101",
			249 => "00000000000000000000010000000101",
			250 => "0000001110000000001110111000001100",
			251 => "0000000000000000000001010100000100",
			252 => "00000000000000000000010000000101",
			253 => "0000001110000000000010000100000100",
			254 => "00000000000000000000010000000101",
			255 => "11111111101001100000010000000101",
			256 => "00000000000000000000010000000101",
			257 => "0000000000000000000001010100100000",
			258 => "0000001111000000000000011100001100",
			259 => "0000000001000000000110101000001000",
			260 => "0000001110000000000100001000000100",
			261 => "00000000000000000000010001010001",
			262 => "00000000010101010000010001010001",
			263 => "11111110111101010000010001010001",
			264 => "0000000111000000000001101000001100",
			265 => "0000001001000000001111000000001000",
			266 => "0000001010000000000100111100000100",
			267 => "00000000000000000000010001010001",
			268 => "00000000100110010000010001010001",
			269 => "00000000000000000000010001010001",
			270 => "0000000111000000001000011000000100",
			271 => "11111111101111110000010001010001",
			272 => "00000000000101100000010001010001",
			273 => "0000000110000000001101111100000100",
			274 => "00000000000000000000010001010001",
			275 => "11111111011101100000010001010001",
			276 => "0000000011000000001100010000011100",
			277 => "0000001001000000000000111100001100",
			278 => "0000001110000000000100001000000100",
			279 => "00000000000000000000010010100101",
			280 => "0000000000000000000101000100000100",
			281 => "00000000001011000000010010100101",
			282 => "00000000000000000000010010100101",
			283 => "0000000001000000000110101000000100",
			284 => "00000000000000000000010010100101",
			285 => "0000001101000000000010011100001000",
			286 => "0000001100000000001000000000000100",
			287 => "11111111101011110000010010100101",
			288 => "00000000000000000000010010100101",
			289 => "00000000000000000000010010100101",
			290 => "0000001010000000000001010000001100",
			291 => "0000000101000000001110101000000100",
			292 => "00000000000000000000010010100101",
			293 => "0000000001000000001101111100000100",
			294 => "00000000001100000000010010100101",
			295 => "00000000000000000000010010100101",
			296 => "00000000000000000000010010100101",
			297 => "0000001101000000001110101100001100",
			298 => "0000001000000000001001111100000100",
			299 => "00000000000000000000010011101001",
			300 => "0000001110000000001110101000000100",
			301 => "11111111110100010000010011101001",
			302 => "00000000000000000000010011101001",
			303 => "0000000001000000000101011100010100",
			304 => "0000001100000000001000011000010000",
			305 => "0000000110000000001011001100001100",
			306 => "0000001100000000001110001100000100",
			307 => "00000000000000000000010011101001",
			308 => "0000001101000000001110101000000100",
			309 => "00000000000000000000010011101001",
			310 => "00000000011001000000010011101001",
			311 => "00000000000000000000010011101001",
			312 => "00000000000000000000010011101001",
			313 => "00000000000000000000010011101001",
			314 => "0000001001000000001100011000011000",
			315 => "0000001100000000001100110000010000",
			316 => "0000000111000000001101100000000100",
			317 => "00000000000000000000010100111101",
			318 => "0000001110000000000100001000000100",
			319 => "00000000000000000000010100111101",
			320 => "0000000000000000000101000100000100",
			321 => "00000000001001010000010100111101",
			322 => "00000000000000000000010100111101",
			323 => "0000001001000000001100011000000100",
			324 => "11111111011010100000010100111101",
			325 => "00000000000000000000010100111101",
			326 => "0000000001000000000000111100010000",
			327 => "0000000111000000001111011100001100",
			328 => "0000000111000000000001111100000100",
			329 => "00000000000000000000010100111101",
			330 => "0000000110000000001011001100000100",
			331 => "00000000011100000000010100111101",
			332 => "00000000000000000000010100111101",
			333 => "00000000000000000000010100111101",
			334 => "00000000000000000000010100111101",
			335 => "0000000101000000000101001000000100",
			336 => "11111111101010100000010101110001",
			337 => "0000000111000000001000011000000100",
			338 => "00000000000000000000010101110001",
			339 => "0000000111000000001111011100010000",
			340 => "0000000010000000001010000100001100",
			341 => "0000001011000000000010001000000100",
			342 => "00000000000000000000010101110001",
			343 => "0000001001000000001000010000000100",
			344 => "00000000101001110000010101110001",
			345 => "00000000000000000000010101110001",
			346 => "00000000000000000000010101110001",
			347 => "00000000000000000000010101110001",
			348 => "0000000111000000001000011000011100",
			349 => "0000001111000000001011000000000100",
			350 => "00000000000000000000010110101101",
			351 => "0000000011000000001100010000001100",
			352 => "0000000111000000000001101000001000",
			353 => "0000001101000000000010011100000100",
			354 => "11111111101111000000010110101101",
			355 => "00000000000000000000010110101101",
			356 => "00000000000000000000010110101101",
			357 => "0000001111000000001100000000000100",
			358 => "00000000000000000000010110101101",
			359 => "0000001111000000001010000100000100",
			360 => "11111111111110100000010110101101",
			361 => "00000000000000000000010110101101",
			362 => "00000000000000000000010110101101",
			363 => "0000000101000000000110100100001100",
			364 => "0000001111000000001000000000000100",
			365 => "00000000000000000000011000000001",
			366 => "0000001110000000001000011000000100",
			367 => "11111111010101000000011000000001",
			368 => "00000000000000000000011000000001",
			369 => "0000001001000000001001100100010100",
			370 => "0000001110000000001011000000000100",
			371 => "00000000000000000000011000000001",
			372 => "0000001101000000000111111100001100",
			373 => "0000001010000000000111110100001000",
			374 => "0000001011000000000100001000000100",
			375 => "00000000000000000000011000000001",
			376 => "00000000011110000000011000000001",
			377 => "00000000000000000000011000000001",
			378 => "00000000000000000000011000000001",
			379 => "0000001101000000001001011100001000",
			380 => "0000000011000000001010000100000100",
			381 => "11111111111001000000011000000001",
			382 => "00000000000000000000011000000001",
			383 => "00000000000000000000011000000001",
			384 => "0000000000000000000001010100100100",
			385 => "0000000101000000001100100100011000",
			386 => "0000000111000000001100101000001100",
			387 => "0000000010000000000100001000000100",
			388 => "00000000000000000000011001011101",
			389 => "0000001100000000001110001100000100",
			390 => "00000000001011000000011001011101",
			391 => "00000000000000000000011001011101",
			392 => "0000001100000000001000000000001000",
			393 => "0000000010000000000110010000000100",
			394 => "11111111110110000000011001011101",
			395 => "00000000000000000000011001011101",
			396 => "00000000000000000000011001011101",
			397 => "0000000110000000000100110100001000",
			398 => "0000001100000000001011000000000100",
			399 => "00000000000000000000011001011101",
			400 => "00000000010100010000011001011101",
			401 => "00000000000000000000011001011101",
			402 => "0000001111000000000110001100001000",
			403 => "0000001010000000000000001000000100",
			404 => "00000000000000000000011001011101",
			405 => "11111111101111010000011001011101",
			406 => "00000000000000000000011001011101",
			407 => "0000000101000000000110100100001100",
			408 => "0000001100000000000110000100001000",
			409 => "0000000110000000001101011100000100",
			410 => "00000000000000000000011011000001",
			411 => "11111110100100110000011011000001",
			412 => "00000000000000000000011011000001",
			413 => "0000000001000000001001011000010000",
			414 => "0000001101000000000010110100000100",
			415 => "00000000000000000000011011000001",
			416 => "0000000101000000000010011100001000",
			417 => "0000000001000000001111001100000100",
			418 => "00000000000000000000011011000001",
			419 => "00000000011110010000011011000001",
			420 => "00000000000000000000011011000001",
			421 => "0000001101000000001010001000001100",
			422 => "0000000101000000001111010000001000",
			423 => "0000001001000000001011001100000100",
			424 => "00000000000000000000011011000001",
			425 => "11111111101111100000011011000001",
			426 => "00000000000000000000011011000001",
			427 => "0000000001000000001101111100001000",
			428 => "0000001001000000001111000000000100",
			429 => "00000000000000000000011011000001",
			430 => "00000000000100100000011011000001",
			431 => "00000000000000000000011011000001",
			432 => "0000001010000000000000001000011000",
			433 => "0000001001000000000101011100010000",
			434 => "0000000001000000000110101000001100",
			435 => "0000000010000000000100001000000100",
			436 => "00000000000000000000011100101101",
			437 => "0000000000000000000011101000000100",
			438 => "00000000011101000000011100101101",
			439 => "00000000000000000000011100101101",
			440 => "00000000000000000000011100101101",
			441 => "0000000010000000001101000100000100",
			442 => "11111111111101010000011100101101",
			443 => "00000000000001010000011100101101",
			444 => "0000000011000000001010000100001100",
			445 => "0000001111000000001111010100001000",
			446 => "0000000001000000000000111100000100",
			447 => "11111111101101110000011100101101",
			448 => "00000000000000000000011100101101",
			449 => "00000000000000000000011100101101",
			450 => "0000001100000000001011000000000100",
			451 => "00000000000000000000011100101101",
			452 => "0000000101000000000010011100001100",
			453 => "0000000001000000000000111100001000",
			454 => "0000000111000000001111011100000100",
			455 => "00000000010110100000011100101101",
			456 => "00000000000000000000011100101101",
			457 => "00000000000000000000011100101101",
			458 => "00000000000000000000011100101101",
			459 => "0000000011000000001100010000011100",
			460 => "0000001001000000000000111100010000",
			461 => "0000000000000000000011101000001100",
			462 => "0000000010000000000100001000000100",
			463 => "00000000000000000000011110010001",
			464 => "0000000100000000000111001000000100",
			465 => "00000000000000000000011110010001",
			466 => "00000000001100100000011110010001",
			467 => "00000000000000000000011110010001",
			468 => "0000001100000000001100110000000100",
			469 => "00000000000000000000011110010001",
			470 => "0000000011000000001001100000000100",
			471 => "11111111101000110000011110010001",
			472 => "00000000000000000000011110010001",
			473 => "0000001001000000001100011000000100",
			474 => "00000000000000000000011110010001",
			475 => "0000000001000000001101111100010000",
			476 => "0000001101000000001111010000000100",
			477 => "00000000000000000000011110010001",
			478 => "0000001010000000000001010000001000",
			479 => "0000001100000000000111001000000100",
			480 => "00000000000000000000011110010001",
			481 => "00000000010001110000011110010001",
			482 => "00000000000000000000011110010001",
			483 => "00000000000000000000011110010001",
			484 => "0000001101000000000111111100011100",
			485 => "0000000011000000001001001000000100",
			486 => "00000000000000000000011111011101",
			487 => "0000001010000000001010100000010100",
			488 => "0000001001000000000100111100010000",
			489 => "0000001100000000000011011100000100",
			490 => "00000000000000000000011111011101",
			491 => "0000001111000000001011000000000100",
			492 => "00000000000000000000011111011101",
			493 => "0000001100000000001011000000000100",
			494 => "00000000011011010000011111011101",
			495 => "00000000000000000000011111011101",
			496 => "00000000000000000000011111011101",
			497 => "00000000000000000000011111011101",
			498 => "0000001010000000001010100000001000",
			499 => "0000000010000000001100000000000100",
			500 => "11111111110000100000011111011101",
			501 => "00000000000000000000011111011101",
			502 => "00000000000000000000011111011101",
			503 => "0000000111000000001000000000010100",
			504 => "0000000010000000000000110100001100",
			505 => "0000000001000000000110101000001000",
			506 => "0000001110000000000100001000000100",
			507 => "00000000000000000000100001010001",
			508 => "00000000010100110000100001010001",
			509 => "00000000000000000000100001010001",
			510 => "0000001100000000000100011000000100",
			511 => "11111111100110010000100001010001",
			512 => "00000000000000000000100001010001",
			513 => "0000001100000000001011000000010000",
			514 => "0000001001000000001111000000001100",
			515 => "0000000111000000001000011000001000",
			516 => "0000000100000000001000001000000100",
			517 => "00000000101010110000100001010001",
			518 => "00000000000000000000100001010001",
			519 => "00000000000000000000100001010001",
			520 => "00000000000000000000100001010001",
			521 => "0000000011000000000110111100001000",
			522 => "0000000101000000001101000100000100",
			523 => "00000000000000000000100001010001",
			524 => "11111111110111110000100001010001",
			525 => "0000000101000000000111100000000100",
			526 => "00000000000000000000100001010001",
			527 => "0000000011000000000010100100001000",
			528 => "0000000011000000001111010100000100",
			529 => "00000000000000000000100001010001",
			530 => "00000000000111100000100001010001",
			531 => "00000000000000000000100001010001",
			532 => "0000000110000000001001011000001100",
			533 => "0000000001000000000110101000001000",
			534 => "0000001110000000000100001000000100",
			535 => "00000000000000000000100010110101",
			536 => "00000000010101000000100010110101",
			537 => "00000000000000000000100010110101",
			538 => "0000000101000000000101001000011000",
			539 => "0000001010000000000111101100000100",
			540 => "00000000000000000000100010110101",
			541 => "0000000011000000001100010000001000",
			542 => "0000001000000000000111110100000100",
			543 => "00000000000000000000100010110101",
			544 => "11111111010011110000100010110101",
			545 => "0000001000000000001000100100000100",
			546 => "00000000000000000000100010110101",
			547 => "0000001000000000000001010000000100",
			548 => "11111111111010100000100010110101",
			549 => "00000000000000000000100010110101",
			550 => "0000001100000000001001110100001100",
			551 => "0000000001000000000101011100001000",
			552 => "0000000011000000001010000100000100",
			553 => "00000000000000000000100010110101",
			554 => "00000000011011010000100010110101",
			555 => "00000000000000000000100010110101",
			556 => "00000000000000000000100010110101",
			557 => "0000001010000000000010101100100000",
			558 => "0000001111000000001001001000001000",
			559 => "0000001100000000000110000100000100",
			560 => "11111111111100100000100011111001",
			561 => "00000000000000000000100011111001",
			562 => "0000000001000000000000111100010100",
			563 => "0000000111000000001000011000010000",
			564 => "0000001100000000001001110100001100",
			565 => "0000001100000000000011011100000100",
			566 => "00000000000000000000100011111001",
			567 => "0000001001000000000100111100000100",
			568 => "00000000011111000000100011111001",
			569 => "00000000000000000000100011111001",
			570 => "00000000000000000000100011111001",
			571 => "00000000000000000000100011111001",
			572 => "00000000000000000000100011111001",
			573 => "00000000000000000000100011111001",
			574 => "0000001010000000000000001000100100",
			575 => "0000000011000000000000110100010100",
			576 => "0000001001000000000101011100010000",
			577 => "0000001100000000001100110000001100",
			578 => "0000001111000000000001111100000100",
			579 => "00000000000000000000100101111101",
			580 => "0000001100000000000100000000000100",
			581 => "00000000000000000000100101111101",
			582 => "00000000001101100000100101111101",
			583 => "00000000000000000000100101111101",
			584 => "11111111101100110000100101111101",
			585 => "0000000110000000000100110100001100",
			586 => "0000001100000000001000000000001000",
			587 => "0000001001000000000100111100000100",
			588 => "00000000100001110000100101111101",
			589 => "00000000000000000000100101111101",
			590 => "00000000000000000000100101111101",
			591 => "00000000000000000000100101111101",
			592 => "0000000011000000001010000100001000",
			593 => "0000001111000000000110111100000100",
			594 => "11111111010011000000100101111101",
			595 => "00000000000000000000100101111101",
			596 => "0000001001000000001111000000001100",
			597 => "0000001001000000001100011000000100",
			598 => "00000000000000000000100101111101",
			599 => "0000000110000000001011001100000100",
			600 => "00000000100000000000100101111101",
			601 => "00000000000000000000100101111101",
			602 => "0000000111000000000001001000001000",
			603 => "0000000000000000000001010100000100",
			604 => "00000000000000000000100101111101",
			605 => "11111111111000000000100101111101",
			606 => "00000000000000000000100101111101",
			607 => "0000000101000000000110100100001100",
			608 => "0000001100000000000110000100001000",
			609 => "0000000110000000001101011100000100",
			610 => "00000000000000000000100111110001",
			611 => "11111110101100100000100111110001",
			612 => "00000000000000000000100111110001",
			613 => "0000000011000000001111010100011100",
			614 => "0000000001000000001001011000010000",
			615 => "0000000011000000000000110100000100",
			616 => "00000000000000000000100111110001",
			617 => "0000001100000000001000000000001000",
			618 => "0000001100000000000011011100000100",
			619 => "00000000000000000000100111110001",
			620 => "00000000001010100000100111110001",
			621 => "00000000000000000000100111110001",
			622 => "0000001100000000000100011000000100",
			623 => "00000000000000000000100111110001",
			624 => "0000001100000000001001110100000100",
			625 => "11111111101011010000100111110001",
			626 => "00000000000000000000100111110001",
			627 => "0000001100000000001000000000000100",
			628 => "00000000000000000000100111110001",
			629 => "0000000001000000001101111100001100",
			630 => "0000001100000000001011011100001000",
			631 => "0000000001000000001111001100000100",
			632 => "00000000000000000000100111110001",
			633 => "00000000010011100000100111110001",
			634 => "00000000000000000000100111110001",
			635 => "00000000000000000000100111110001",
			636 => "0000001110000000001010001000011100",
			637 => "0000000000000000001100011100011000",
			638 => "0000001010000000000100111100010000",
			639 => "0000000101000000000001101000001100",
			640 => "0000000011000000000110100100000100",
			641 => "00000000000000000000101001110101",
			642 => "0000000110000000000000111100000100",
			643 => "00000000001101100000101001110101",
			644 => "00000000000000000000101001110101",
			645 => "11111111011100110000101001110101",
			646 => "0000001111000000000010001000000100",
			647 => "00000000000000000000101001110101",
			648 => "00000000010110110000101001110101",
			649 => "11111110110000010000101001110101",
			650 => "0000000001000000000000111100011100",
			651 => "0000000011000000001010000100010100",
			652 => "0000000110000000000100110100001100",
			653 => "0000001101000000000111111100001000",
			654 => "0000001010000000000000001000000100",
			655 => "00000000110110010000101001110101",
			656 => "00000000000000000000101001110101",
			657 => "00000000000000000000101001110101",
			658 => "0000000001000000001001011000000100",
			659 => "00000000000000000000101001110101",
			660 => "11111111011101000000101001110101",
			661 => "0000000110000000001011001100000100",
			662 => "00000000111000010000101001110101",
			663 => "00000000000000000000101001110101",
			664 => "0000000101000000001110010000000100",
			665 => "11111111100111110000101001110101",
			666 => "0000001010000000000110011000000100",
			667 => "00000000001011100000101001110101",
			668 => "00000000000000000000101001110101",
			669 => "0000000000000000000001010100110000",
			670 => "0000000101000000001100100100011100",
			671 => "0000001100000000000100011000010000",
			672 => "0000000111000000001101100000000100",
			673 => "00000000000000000000101100001001",
			674 => "0000001110000000000100001000000100",
			675 => "00000000000000000000101100001001",
			676 => "0000001010000000000111101100000100",
			677 => "00000000011011100000101100001001",
			678 => "00000000000000000000101100001001",
			679 => "0000000100000000001100000000001000",
			680 => "0000001001000000001111000000000100",
			681 => "00000000000000000000101100001001",
			682 => "11111111100110000000101100001001",
			683 => "00000000000000000000101100001001",
			684 => "0000000001000000001001011000000100",
			685 => "00000000000000000000101100001001",
			686 => "0000001001000000000100111100001100",
			687 => "0000001101000000000010011100000100",
			688 => "00000000000000000000101100001001",
			689 => "0000001100000000000100011000000100",
			690 => "00000000000000000000101100001001",
			691 => "00000001000010000000101100001001",
			692 => "00000000000000000000101100001001",
			693 => "0000001011000000000101100100001000",
			694 => "0000000000000000000001110000000100",
			695 => "00000000000000000000101100001001",
			696 => "11111110111010100000101100001001",
			697 => "0000001011000000000110110100001000",
			698 => "0000001001000000000100111100000100",
			699 => "00000000010000000000101100001001",
			700 => "00000000000000000000101100001001",
			701 => "0000000101000000001110010000001000",
			702 => "0000001100000000000100011000000100",
			703 => "00000000000000000000101100001001",
			704 => "11111111100110100000101100001001",
			705 => "00000000000000000000101100001001",
			706 => "0000000000000000000001010100101000",
			707 => "0000000011000000000110111100100100",
			708 => "0000000110000000001101111100011000",
			709 => "0000000111000000001101100000000100",
			710 => "00000000000000000000101101111101",
			711 => "0000001010000000000100111100001100",
			712 => "0000000101000000000001101000001000",
			713 => "0000001110000000000100001000000100",
			714 => "00000000000000000000101101111101",
			715 => "00000000011000010000101101111101",
			716 => "11111111110110010000101101111101",
			717 => "0000001111000000000000110100000100",
			718 => "00000000000000000000101101111101",
			719 => "00000000110000000000101101111101",
			720 => "0000000110000000001101111100001000",
			721 => "0000001010000000000000001000000100",
			722 => "00000000000000000000101101111101",
			723 => "11111111100001100000101101111101",
			724 => "00000000000000000000101101111101",
			725 => "00000000111011000000101101111101",
			726 => "0000000011000000001000001100001000",
			727 => "0000000010000000000110101100000100",
			728 => "11111111000101100000101101111101",
			729 => "00000000000000000000101101111101",
			730 => "0000000001000000000101011100001000",
			731 => "0000001011000000000101110100000100",
			732 => "00000000010111110000101101111101",
			733 => "00000000000000000000101101111101",
			734 => "11111111101100100000101101111101",
			735 => "0000000011000000001000001100101100",
			736 => "0000001000000000001000100100101000",
			737 => "0000001100000000001100110000010000",
			738 => "0000000001000000000111100100001100",
			739 => "0000000010000000000100001000000100",
			740 => "00000000000000000000101111110001",
			741 => "0000000001000000000010001100000100",
			742 => "00000000000000000000101111110001",
			743 => "00000000010111010000101111110001",
			744 => "00000000000000000000101111110001",
			745 => "0000000011000000001100010000010000",
			746 => "0000000001000000000110101000000100",
			747 => "00000000000000000000101111110001",
			748 => "0000001100000000001000000000001000",
			749 => "0000001101000000000010011100000100",
			750 => "11111111100011110000101111110001",
			751 => "00000000000000000000101111110001",
			752 => "00000000000000000000101111110001",
			753 => "0000000001000000001001011000000100",
			754 => "00000000011000100000101111110001",
			755 => "00000000000000000000101111110001",
			756 => "11111111101101010000101111110001",
			757 => "0000000110000000001000010000001100",
			758 => "0000001100000000001011000000000100",
			759 => "00000000000000000000101111110001",
			760 => "0000000001000000001101111100000100",
			761 => "00000000011100100000101111110001",
			762 => "00000000000000000000101111110001",
			763 => "00000000000000000000101111110001",
			764 => "0000001010000000001010100000110000",
			765 => "0000001110000000000101110100010100",
			766 => "0000001100000000000100000000001000",
			767 => "0000000111000000001001110000000100",
			768 => "11111110101000010000110010011101",
			769 => "00000101000111100000110010011101",
			770 => "0000000010000000000001101000000100",
			771 => "11111110011010010000110010011101",
			772 => "0000001001000000001011111100000100",
			773 => "00000010011111010000110010011101",
			774 => "11111110010110000000110010011101",
			775 => "0000001001000000000100111100011000",
			776 => "0000000011000000000111010100010100",
			777 => "0000000101000000001111010000001100",
			778 => "0000001110000000001110101000000100",
			779 => "00000001110001110000110010011101",
			780 => "0000000010000000000010000100000100",
			781 => "00000010110011010000110010011101",
			782 => "00000011110110000000110010011101",
			783 => "0000000010000000000010000100000100",
			784 => "00000010110010110000110010011101",
			785 => "11111110000001010000110010011101",
			786 => "00000101000101010000110010011101",
			787 => "11111110011110110000110010011101",
			788 => "0000001010000000000010101100010100",
			789 => "0000000010000000001010000100001100",
			790 => "0000000011000000001000001100000100",
			791 => "11111110010111110000110010011101",
			792 => "0000000111000000001000011000000100",
			793 => "00000010110110000000110010011101",
			794 => "11111110011101100000110010011101",
			795 => "0000000001000000000101011100000100",
			796 => "00000101010100100000110010011101",
			797 => "11111110100110100000110010011101",
			798 => "0000001010000000000010101100001000",
			799 => "0000001101000000000100101000000100",
			800 => "11111110011110110000110010011101",
			801 => "00000001010111100000110010011101",
			802 => "0000001101000000000011000000000100",
			803 => "11111110010111000000110010011101",
			804 => "0000001011000000000111111100000100",
			805 => "00000010110011110000110010011101",
			806 => "11111110011000100000110010011101",
			807 => "0000000100000000001111100100111000",
			808 => "0000000011000000001111010100101000",
			809 => "0000001010000000000000001000011100",
			810 => "0000001011000000000100001000001100",
			811 => "0000000001000000000110101000001000",
			812 => "0000001110000000000100001000000100",
			813 => "00000000000000000000110100011001",
			814 => "00000000001001000000110100011001",
			815 => "11111111101011000000110100011001",
			816 => "0000000001000000000000111100001100",
			817 => "0000001110000000001110101000000100",
			818 => "00000000000000000000110100011001",
			819 => "0000001111000000000010000100000100",
			820 => "00000000100011010000110100011001",
			821 => "00000000000000000000110100011001",
			822 => "00000000000000000000110100011001",
			823 => "0000000000000000000101000100000100",
			824 => "00000000000000000000110100011001",
			825 => "0000000110000000001101111100000100",
			826 => "00000000000000000000110100011001",
			827 => "11111111010101100000110100011001",
			828 => "0000001011000000000101110100001100",
			829 => "0000001001000000001000010000001000",
			830 => "0000000001000000000000111100000100",
			831 => "00000000010100110000110100011001",
			832 => "00000000000000000000110100011001",
			833 => "00000000000000000000110100011001",
			834 => "00000000000000000000110100011001",
			835 => "0000001101000000001111101000000100",
			836 => "11111111011011010000110100011001",
			837 => "00000000000000000000110100011001",
			838 => "0000000100000000001111100100111000",
			839 => "0000000111000000001100101000010000",
			840 => "0000000111000000001101100000000100",
			841 => "00000000000000000000110110011101",
			842 => "0000000001000000000111100100001000",
			843 => "0000001111000000000001111100000100",
			844 => "00000000000000000000110110011101",
			845 => "00000000100000100000110110011101",
			846 => "00000000000000000000110110011101",
			847 => "0000000011000000001001100000001000",
			848 => "0000001111000000000010000000000100",
			849 => "11111111010011010000110110011101",
			850 => "00000000000000000000110110011101",
			851 => "0000000110000000001101111100001000",
			852 => "0000001101000000000111111100000100",
			853 => "00000000100101010000110110011101",
			854 => "00000000000000000000110110011101",
			855 => "0000000011000000000110111100001100",
			856 => "0000001010000000000000001000000100",
			857 => "00000000000000000000110110011101",
			858 => "0000000111000000000110100100000100",
			859 => "00000000000000000000110110011101",
			860 => "11111111011111010000110110011101",
			861 => "0000001001000000001111000000000100",
			862 => "00000000011010000000110110011101",
			863 => "0000000011000000001000001100000100",
			864 => "11111111110000110000110110011101",
			865 => "00000000000000000000110110011101",
			866 => "0000001111000000000110001100001000",
			867 => "0000000100000000000110111000000100",
			868 => "00000000000000000000110110011101",
			869 => "11111111000000000000110110011101",
			870 => "00000000000000000000110110011101",
			871 => "0000000011000000001100000000101000",
			872 => "0000000110000000001101111100100000",
			873 => "0000001110000000000110100100001000",
			874 => "0000000110000000001111001100000100",
			875 => "00000000000000000000111000110001",
			876 => "11111111101000100000111000110001",
			877 => "0000001100000000001110001100010000",
			878 => "0000001011000000000100001000000100",
			879 => "00000000000000000000111000110001",
			880 => "0000001111000000001010011100000100",
			881 => "00000000000000000000111000110001",
			882 => "0000000111000000001100101000000100",
			883 => "00000000100010000000111000110001",
			884 => "00000000000000000000111000110001",
			885 => "0000001011000000000110100100000100",
			886 => "11111111101100010000111000110001",
			887 => "00000000001010010000111000110001",
			888 => "0000001010000000000111101100000100",
			889 => "00000000000000000000111000110001",
			890 => "11111110111101110000111000110001",
			891 => "0000001001000000001100011000000100",
			892 => "00000000000000000000111000110001",
			893 => "0000001001000000000100111100011000",
			894 => "0000000111000000001000011000001100",
			895 => "0000000110000000001101111100000100",
			896 => "00000000000000000000111000110001",
			897 => "0000000011000000000111011000000100",
			898 => "00000000000000000000111000110001",
			899 => "00000000110011000000111000110001",
			900 => "0000001011000000000100010000001000",
			901 => "0000001011000000000010001000000100",
			902 => "00000000000000000000111000110001",
			903 => "00000000001101000000111000110001",
			904 => "00000000000000000000111000110001",
			905 => "0000000011000000001000100000000100",
			906 => "00000000000000000000111000110001",
			907 => "00000000000001000000111000110001",
			908 => "0000001100000000000011011100001000",
			909 => "0000000110000000001101011100000100",
			910 => "00000000000000000000111010110101",
			911 => "11111111000001100000111010110101",
			912 => "0000000011000000001000100000101100",
			913 => "0000001000000000001000100100100000",
			914 => "0000001011000000000010001000010100",
			915 => "0000000010000000001101000100001100",
			916 => "0000001100000000000110000100001000",
			917 => "0000000110000000001001011000000100",
			918 => "00000000000000000000111010110101",
			919 => "00000000011100100000111010110101",
			920 => "11111111100000010000111010110101",
			921 => "0000000001000000001001011000000100",
			922 => "00000000110100100000111010110101",
			923 => "00000000000000000000111010110101",
			924 => "0000000011000000001010000100001000",
			925 => "0000000010000000001110110100000100",
			926 => "00000000000000000000111010110101",
			927 => "11111111101000110000111010110101",
			928 => "00000000000000000000111010110101",
			929 => "0000000011000000001011111000001000",
			930 => "0000000010000000001000100000000100",
			931 => "11111111011110000000111010110101",
			932 => "00000000000000000000111010110101",
			933 => "00000000000000000000111010110101",
			934 => "0000000110000000001000010000001100",
			935 => "0000001100000000001000000000000100",
			936 => "00000000000000000000111010110101",
			937 => "0000000001000000001101111100000100",
			938 => "00000000101000010000111010110101",
			939 => "00000000000000000000111010110101",
			940 => "00000000000000000000111010110101",
			941 => "0000000111000000001101100000000100",
			942 => "11111111000000000000111100111001",
			943 => "0000000011000000001010000100101000",
			944 => "0000001000000000001000100100011100",
			945 => "0000000010000000001101000100010000",
			946 => "0000001001000000000000111100001000",
			947 => "0000001110000000000100001000000100",
			948 => "00000000000000000000111100111001",
			949 => "00000000010101110000111100111001",
			950 => "0000001001000000001110010100000100",
			951 => "11111111011001110000111100111001",
			952 => "00000000000000000000111100111001",
			953 => "0000001001000000001111000000001000",
			954 => "0000000110000000001101111100000100",
			955 => "00000000110011010000111100111001",
			956 => "00000000000000000000111100111001",
			957 => "00000000000000000000111100111001",
			958 => "0000001100000000001001110100001000",
			959 => "0000001100000000001011000000000100",
			960 => "00000000000000000000111100111001",
			961 => "11111111001100110000111100111001",
			962 => "00000000000000000000111100111001",
			963 => "0000000111000000001111011100001000",
			964 => "0000001001000000001000010000000100",
			965 => "00000000110011110000111100111001",
			966 => "00000000000000000000111100111001",
			967 => "0000000101000000001110010000000100",
			968 => "11111111101011000000111100111001",
			969 => "0000000110000000001000010000001000",
			970 => "0000001001000000001010100000000100",
			971 => "00000000010100110000111100111001",
			972 => "00000000000000000000111100111001",
			973 => "00000000000000000000111100111001",
			974 => "0000000000000000001011010101000000",
			975 => "0000001001000000001111000000011000",
			976 => "0000000111000000001101100000000100",
			977 => "00000000000000000000111111001101",
			978 => "0000001100000000001000000000010000",
			979 => "0000000111000000001000011000001100",
			980 => "0000001110000000001110101000001000",
			981 => "0000001111000000001001110100000100",
			982 => "00000000111100010000111111001101",
			983 => "11111111111000010000111111001101",
			984 => "00000000111101110000111111001101",
			985 => "00000000000000000000111111001101",
			986 => "00000000000000000000111111001101",
			987 => "0000001011000000000010001000001100",
			988 => "0000000001000000001001011000000100",
			989 => "00000000000000000000111111001101",
			990 => "0000001000000000000111110100000100",
			991 => "00000000000000000000111111001101",
			992 => "11111111000100100000111111001101",
			993 => "0000001011000000000100010000010000",
			994 => "0000001010000000001010100000001000",
			995 => "0000000110000000000100110100000100",
			996 => "00000000111110110000111111001101",
			997 => "00000000000000000000111111001101",
			998 => "0000000010000000000111011000000100",
			999 => "11111111100010010000111111001101",
			1000 => "00000000000000000000111111001101",
			1001 => "0000000110000000001010011000000100",
			1002 => "11111111000101000000111111001101",
			1003 => "0000001010000000001010100100000100",
			1004 => "00000000101001100000111111001101",
			1005 => "00000000000000000000111111001101",
			1006 => "0000001111000000000110001100000100",
			1007 => "11111110101001110000111111001101",
			1008 => "0000000110000000001000010000000100",
			1009 => "00000000100011000000111111001101",
			1010 => "00000000000000000000111111001101",
			1011 => "0000001000000000001000100100101100",
			1012 => "0000001111000000000001001000011100",
			1013 => "0000001111000000000010001000011000",
			1014 => "0000001100000000001000111100001000",
			1015 => "0000001110000000000100001000000100",
			1016 => "11001110010101000001000010001001",
			1017 => "11011000100000110001000010001001",
			1018 => "0000001111000000001011011100001100",
			1019 => "0000001110000000001011000000000100",
			1020 => "11001110001111000001000010001001",
			1021 => "0000001001000000000001000100000100",
			1022 => "11010101111010000001000010001001",
			1023 => "11001110010000010001000010001001",
			1024 => "11010000111001110001000010001001",
			1025 => "11010100011110000001000010001001",
			1026 => "0000001001000000001111000000001000",
			1027 => "0000000010000000000111100000000100",
			1028 => "11100011100110010001000010001001",
			1029 => "11101111111101110001000010001001",
			1030 => "0000001101000000000100101000000100",
			1031 => "11001110010011110001000010001001",
			1032 => "11100011100110010001000010001001",
			1033 => "0000001000000000001000100100001100",
			1034 => "0000001001000000001111000000000100",
			1035 => "11101001110000000001000010001001",
			1036 => "0000001111000000001100000000000100",
			1037 => "11001110010110010001000010001001",
			1038 => "11010110000110010001000010001001",
			1039 => "0000001000000000001001000100010100",
			1040 => "0000000010000000001010000100010000",
			1041 => "0000001001000000001111000000001000",
			1042 => "0000000010000000000111100000000100",
			1043 => "11001110100111010001000010001001",
			1044 => "11010111010011000001000010001001",
			1045 => "0000000011000000000000010000000100",
			1046 => "11001110001111100001000010001001",
			1047 => "11010010000111000001000010001001",
			1048 => "11011011101010010001000010001001",
			1049 => "0000001010000000000010101100010000",
			1050 => "0000000100000000001101101100001000",
			1051 => "0000001010000000001010100100000100",
			1052 => "11010000001111000001000010001001",
			1053 => "11001110001111100001000010001001",
			1054 => "0000001000000000001010110000000100",
			1055 => "11010011110001110001000010001001",
			1056 => "11001110011001010001000010001001",
			1057 => "11001110001110010001000010001001",
			1058 => "0000000000000000001011010101001000",
			1059 => "0000000110000000000100110100101000",
			1060 => "0000001110000000001110101000010100",
			1061 => "0000000110000000000001000100010000",
			1062 => "0000001100000000000110000100001100",
			1063 => "0000001110000000000100001000000100",
			1064 => "11111111111001010001000100110101",
			1065 => "0000001001000000000101011100000100",
			1066 => "00000001010011000001000100110101",
			1067 => "00000000011010010001000100110101",
			1068 => "11111111101111010001000100110101",
			1069 => "11111110011110100001000100110101",
			1070 => "0000001001000000000100111100010000",
			1071 => "0000000111000000001111011100001100",
			1072 => "0000001001000000001111000000000100",
			1073 => "00000001100000100001000100110101",
			1074 => "0000000111000000001000011000000100",
			1075 => "11111111111110110001000100110101",
			1076 => "00000001101011110001000100110101",
			1077 => "00000000000000000001000100110101",
			1078 => "11111111101001110001000100110101",
			1079 => "0000000011000000001000001100010100",
			1080 => "0000000010000000000010000100001100",
			1081 => "0000000101000000000001000000001000",
			1082 => "0000001000000000001000100100000100",
			1083 => "00000000000000000001000100110101",
			1084 => "11111110111111110001000100110101",
			1085 => "00000000110101010001000100110101",
			1086 => "0000000001000000001001011000000100",
			1087 => "00000000000000000001000100110101",
			1088 => "11111110100101010001000100110101",
			1089 => "0000000001000000000101011100001000",
			1090 => "0000001100000000001001110100000100",
			1091 => "00000001010010100001000100110101",
			1092 => "00000000000000000001000100110101",
			1093 => "00000000000000000001000100110101",
			1094 => "0000001111000000000110001100000100",
			1095 => "11111110011011010001000100110101",
			1096 => "0000000110000000000101010000001000",
			1097 => "0000000001000000000100110100000100",
			1098 => "00000001100110110001000100110101",
			1099 => "00000000000000000001000100110101",
			1100 => "11111110111100110001000100110101",
			1101 => "0000000100000000001111100101000100",
			1102 => "0000001001000000000101011100010000",
			1103 => "0000000000000000000011101000001100",
			1104 => "0000001111000000000001111100000100",
			1105 => "00000000000000000001000111010001",
			1106 => "0000000001000000000111100100000100",
			1107 => "00000000011011010001000111010001",
			1108 => "00000000000000000001000111010001",
			1109 => "00000000000000000001000111010001",
			1110 => "0000000011000000001001100000010100",
			1111 => "0000000001000000001101011100001000",
			1112 => "0000001001000000001110010100000100",
			1113 => "11111111111100010001000111010001",
			1114 => "00000000000000000001000111010001",
			1115 => "0000001001000000001101011000000100",
			1116 => "00000000000000000001000111010001",
			1117 => "0000000010000000001110010000000100",
			1118 => "11111111001110010001000111010001",
			1119 => "00000000000000000001000111010001",
			1120 => "0000000110000000001101111100001000",
			1121 => "0000001101000000000111111100000100",
			1122 => "00000000100011110001000111010001",
			1123 => "00000000000000000001000111010001",
			1124 => "0000000011000000000110111100001100",
			1125 => "0000001010000000000000001000000100",
			1126 => "00000000000000000001000111010001",
			1127 => "0000001100000000001010111000000100",
			1128 => "00000000000000000001000111010001",
			1129 => "11111111100110110001000111010001",
			1130 => "0000001011000000000101110100001000",
			1131 => "0000000101000000000111100000000100",
			1132 => "00000000000000000001000111010001",
			1133 => "00000000001110100001000111010001",
			1134 => "00000000000000000001000111010001",
			1135 => "0000001111000000000110001100001000",
			1136 => "0000000100000000000110111000000100",
			1137 => "00000000000000000001000111010001",
			1138 => "11111111000011000001000111010001",
			1139 => "00000000000000000001000111010001",
			1140 => "0000000000000000001101010001000000",
			1141 => "0000001100000000000001111100011100",
			1142 => "0000000110000000000001000100010100",
			1143 => "0000000001000000000111100100010000",
			1144 => "0000001110000000000100001000000100",
			1145 => "00000000000000000001001001010101",
			1146 => "0000001100000000001100110000001000",
			1147 => "0000000111000000001101100000000100",
			1148 => "00000000000000000001001001010101",
			1149 => "00000000010001000001001001010101",
			1150 => "00000000000000000001001001010101",
			1151 => "00000000000000000001001001010101",
			1152 => "0000000111000000001000000000000100",
			1153 => "11111111011111110001001001010101",
			1154 => "00000000000000000001001001010101",
			1155 => "0000000001000000001001011000001000",
			1156 => "0000001001000000001100011000000100",
			1157 => "00000000000000000001001001010101",
			1158 => "00000000101100000001001001010101",
			1159 => "0000000011000000001111010100001100",
			1160 => "0000000001000000001001011000001000",
			1161 => "0000000101000000001101000100000100",
			1162 => "00000000000000000001001001010101",
			1163 => "11111111110011110001001001010101",
			1164 => "00000000000000000001001001010101",
			1165 => "0000000001000000000000111100001000",
			1166 => "0000000101000000001111010000000100",
			1167 => "00000000010001100001001001010101",
			1168 => "00000000000000000001001001010101",
			1169 => "0000000101000000001100010000000100",
			1170 => "11111111111100100001001001010101",
			1171 => "00000000000000000001001001010101",
			1172 => "11111111100111010001001001010101",
			1173 => "0000000111000000001101100000000100",
			1174 => "11111110111011100001001011101001",
			1175 => "0000000011000000001010000100101000",
			1176 => "0000000000000000000101000100011000",
			1177 => "0000000010000000001101000100010000",
			1178 => "0000001001000000000000111100001000",
			1179 => "0000001110000000000100001000000100",
			1180 => "00000000000000000001001011101001",
			1181 => "00000000100101000001001011101001",
			1182 => "0000001001000000001110010100000100",
			1183 => "11111111010000010001001011101001",
			1184 => "00000000000000000001001011101001",
			1185 => "0000000110000000001101111100000100",
			1186 => "00000000110000010001001011101001",
			1187 => "00000000000000000001001011101001",
			1188 => "0000001000000000001000100100000100",
			1189 => "00000000000000000001001011101001",
			1190 => "0000001011000000000110110100000100",
			1191 => "00000000000000000001001011101001",
			1192 => "0000000010000000000111011000000100",
			1193 => "11111111000010010001001011101001",
			1194 => "00000000000000000001001011101001",
			1195 => "0000000111000000001111011100010000",
			1196 => "0000001001000000001000010000001100",
			1197 => "0000000001000000000000111100001000",
			1198 => "0000000110000000000100110100000100",
			1199 => "00000000000000000001001011101001",
			1200 => "00000001000010000001001011101001",
			1201 => "00000000000000000001001011101001",
			1202 => "00000000000000000001001011101001",
			1203 => "0000001101000000000110010000000100",
			1204 => "11111111100101010001001011101001",
			1205 => "0000000110000000001000010000001000",
			1206 => "0000000001000000001101111100000100",
			1207 => "00000000010100010001001011101001",
			1208 => "00000000000000000001001011101001",
			1209 => "00000000000000000001001011101001",
			1210 => "0000000000000000001011010101010100",
			1211 => "0000001001000000001111000000100100",
			1212 => "0000000000000000001010100100010000",
			1213 => "0000001001000000000000111100001100",
			1214 => "0000001111000000000001111100000100",
			1215 => "00000000000000000001001110100101",
			1216 => "0000000111000000001101100000000100",
			1217 => "00000000000000000001001110100101",
			1218 => "00000001011101100001001110100101",
			1219 => "00000000000000000001001110100101",
			1220 => "0000000011000000000000110100001000",
			1221 => "0000001001000000000101011100000100",
			1222 => "00000000000000000001001110100101",
			1223 => "11111111001101100001001110100101",
			1224 => "0000001100000000001000000000001000",
			1225 => "0000000111000000001000011000000100",
			1226 => "00000001000000000001001110100101",
			1227 => "00000000000000000001001110100101",
			1228 => "00000000000000000001001110100101",
			1229 => "0000000011000000000111010100011000",
			1230 => "0000000000000000000101000100001100",
			1231 => "0000001101000000000101110000001000",
			1232 => "0000001100000000000100011000000100",
			1233 => "00000000000000000001001110100101",
			1234 => "11111111101101000001001110100101",
			1235 => "00000000110010110001001110100101",
			1236 => "0000000111000000001111011100001000",
			1237 => "0000001100000000001011000000000100",
			1238 => "00000000000000000001001110100101",
			1239 => "11111110100011110001001110100101",
			1240 => "00000000000000000001001110100101",
			1241 => "0000001100000000001001110100001100",
			1242 => "0000001011000000000010001000000100",
			1243 => "00000000000000000001001110100101",
			1244 => "0000000001000000000101011100000100",
			1245 => "00000000111111110001001110100101",
			1246 => "00000000000000000001001110100101",
			1247 => "0000000110000000001010011000000100",
			1248 => "11111111001010100001001110100101",
			1249 => "0000001101000000001110010000000100",
			1250 => "00000000010001010001001110100101",
			1251 => "00000000000000000001001110100101",
			1252 => "0000001111000000000110001100000100",
			1253 => "11111110100100110001001110100101",
			1254 => "0000000110000000001000010000000100",
			1255 => "00000000101011110001001110100101",
			1256 => "00000000000000000001001110100101",
			1257 => "0000001000000000001000100100110100",
			1258 => "0000001110000000000101110100011100",
			1259 => "0000000110000000001101011100001000",
			1260 => "0000000011000000001010111100000100",
			1261 => "11111110101101010001010001110001",
			1262 => "00000110001111100001010001110001",
			1263 => "0000001100000000000100000000000100",
			1264 => "00000000110011110001010001110001",
			1265 => "0000001011000000000100001000000100",
			1266 => "11111110010001110001010001110001",
			1267 => "0000001001000000000001000100001000",
			1268 => "0000001100000000001100110000000100",
			1269 => "00000100001001100001010001110001",
			1270 => "11111111000110010001010001110001",
			1271 => "11111110011011110001010001110001",
			1272 => "0000001001000000000100111100010100",
			1273 => "0000000011000000000111010100010000",
			1274 => "0000001110000000000010000100001100",
			1275 => "0000000111000000000100001000000100",
			1276 => "00000100010110110001010001110001",
			1277 => "0000001111000000001111010000000100",
			1278 => "00000000111010000001010001110001",
			1279 => "00000011001111110001010001110001",
			1280 => "00000001011011110001010001110001",
			1281 => "00000111100111010001010001110001",
			1282 => "11111110011100100001010001110001",
			1283 => "0000001010000000000010101100100000",
			1284 => "0000000011000000001000100000011100",
			1285 => "0000000010000000001010000100010100",
			1286 => "0000000011000000001000001100001100",
			1287 => "0000001010000000001010100000001000",
			1288 => "0000001111000000000111011000000100",
			1289 => "11111110100010010001010001110001",
			1290 => "00000001011000100001010001110001",
			1291 => "11111110010111100001010001110001",
			1292 => "0000001110000000000111011000000100",
			1293 => "00000100001100110001010001110001",
			1294 => "11111110011101000001010001110001",
			1295 => "0000000010000000000111010100000100",
			1296 => "00000100010010010001010001110001",
			1297 => "11111110100010010001010001110001",
			1298 => "00001001011001100001010001110001",
			1299 => "0000001010000000000010101100001000",
			1300 => "0000001101000000000100101000000100",
			1301 => "11111110011101100001010001110001",
			1302 => "00000001100100010001010001110001",
			1303 => "0000001101000000000011000000000100",
			1304 => "11111110010110100001010001110001",
			1305 => "0000001011000000000111111100000100",
			1306 => "00000011100111010001010001110001",
			1307 => "11111110010111110001010001110001",
			1308 => "0000000000000000001011010100111100",
			1309 => "0000001100000000000001101000111000",
			1310 => "0000001000000000000111110100011100",
			1311 => "0000000010000000001100100100010100",
			1312 => "0000000001000000000111100100001100",
			1313 => "0000001110000000001011000000001000",
			1314 => "0000001100000000000110000100000100",
			1315 => "11111111011111000001010100001101",
			1316 => "00000000010001000001010100001101",
			1317 => "00000001011001100001010100001101",
			1318 => "0000001100000000001100110000000100",
			1319 => "00000000000000000001010100001101",
			1320 => "11111110110011110001010100001101",
			1321 => "0000001001000000001001100100000100",
			1322 => "00000001011010110001010100001101",
			1323 => "00000000000000000001010100001101",
			1324 => "0000000011000000001100010000001000",
			1325 => "0000001010000000000111101100000100",
			1326 => "00000000000000000001010100001101",
			1327 => "11111110001101000001010100001101",
			1328 => "0000001010000000000000001000000100",
			1329 => "00000001010010110001010100001101",
			1330 => "0000000011000000001010000100001000",
			1331 => "0000001011000000000010001000000100",
			1332 => "00000000001101010001010100001101",
			1333 => "11111110010010000001010100001101",
			1334 => "0000000000000000000001010100000100",
			1335 => "00000001011001000001010100001101",
			1336 => "00000000000000000001010100001101",
			1337 => "00000010110011000001010100001101",
			1338 => "0000001011000000000101100100000100",
			1339 => "11111110011010000001010100001101",
			1340 => "0000001011000000001011011100001000",
			1341 => "0000001110000000000110111100000100",
			1342 => "00000001000001100001010100001101",
			1343 => "00000000000000000001010100001101",
			1344 => "0000000101000000001111100100000100",
			1345 => "11111110101100110001010100001101",
			1346 => "00000000000000000001010100001101",
			1347 => "0000001001000000000100111101000100",
			1348 => "0000001110000000001010001000100000",
			1349 => "0000000000000000001100011100011000",
			1350 => "0000000111000000000000001100010000",
			1351 => "0000001100000000000011011100000100",
			1352 => "00000000000000000001010110100001",
			1353 => "0000001101000000001000011000000100",
			1354 => "00000000000000000001010110100001",
			1355 => "0000001100000000000110000100000100",
			1356 => "00000000010100100001010110100001",
			1357 => "00000000000000000001010110100001",
			1358 => "0000001101000000000000110100000100",
			1359 => "11111111111101000001010110100001",
			1360 => "00000000000000000001010110100001",
			1361 => "0000001000000000000011101000000100",
			1362 => "00000000000000000001010110100001",
			1363 => "11111111001101000001010110100001",
			1364 => "0000000111000000001111011100100000",
			1365 => "0000000111000000001000011000011000",
			1366 => "0000001011000000000110110100001100",
			1367 => "0000000111000000000001101000001000",
			1368 => "0000000000000000000010101000000100",
			1369 => "00000000100001010001010110100001",
			1370 => "00000000000000000001010110100001",
			1371 => "00000000000000000001010110100001",
			1372 => "0000000000000000000101000100000100",
			1373 => "00000000000000000001010110100001",
			1374 => "0000001100000000001011000000000100",
			1375 => "00000000000000000001010110100001",
			1376 => "11111111011110010001010110100001",
			1377 => "0000000011000000001100000000000100",
			1378 => "00000000000000000001010110100001",
			1379 => "00000000101110000001010110100001",
			1380 => "00000000000000000001010110100001",
			1381 => "0000000001000000000000111100000100",
			1382 => "00000000000000000001010110100001",
			1383 => "11111111011110010001010110100001",
			1384 => "0000000000000000000011101000001100",
			1385 => "0000000001000000000111100100001000",
			1386 => "0000001110000000000100001000000100",
			1387 => "00000000000000000001011000111101",
			1388 => "00000000100110010001011000111101",
			1389 => "00000000000000000001011000111101",
			1390 => "0000000111000000001000000000001100",
			1391 => "0000000110000000000001000100000100",
			1392 => "00000000000000000001011000111101",
			1393 => "0000001100000000001010111100000100",
			1394 => "11111110110110010001011000111101",
			1395 => "00000000000000000001011000111101",
			1396 => "0000000001000000001001011000001100",
			1397 => "0000000110000000001011001100001000",
			1398 => "0000001110000000001110101000000100",
			1399 => "00000000000000000001011000111101",
			1400 => "00000000110110100001011000111101",
			1401 => "00000000000000000001011000111101",
			1402 => "0000000011000000001100000000010000",
			1403 => "0000000110000000001101111100000100",
			1404 => "00000000000000000001011000111101",
			1405 => "0000000111000000001001001000000100",
			1406 => "00000000000000000001011000111101",
			1407 => "0000001100000000000100011000000100",
			1408 => "00000000000000000001011000111101",
			1409 => "11111111001011110001011000111101",
			1410 => "0000001100000000001000000000010000",
			1411 => "0000000110000000000100110100001000",
			1412 => "0000001011000000000101100100000100",
			1413 => "00000000000000000001011000111101",
			1414 => "00000000101000100001011000111101",
			1415 => "0000001101000000001010001000000100",
			1416 => "11111111111110000001011000111101",
			1417 => "00000000000000000001011000111101",
			1418 => "0000000010000000001110110100000100",
			1419 => "00000000000000000001011000111101",
			1420 => "0000000100000000000000010000000100",
			1421 => "11111111011001110001011000111101",
			1422 => "00000000000000000001011000111101",
			1423 => "0000000000000000001101010001000000",
			1424 => "0000000111000000001000000000010100",
			1425 => "0000000000000000000110011100010000",
			1426 => "0000001111000000001011000000000100",
			1427 => "00000000000000000001011011000001",
			1428 => "0000000001000000000111100100001000",
			1429 => "0000001100000000000011011100000100",
			1430 => "00000000000000000001011011000001",
			1431 => "00000000101101110001011011000001",
			1432 => "00000000000000000001011011000001",
			1433 => "11111111001001000001011011000001",
			1434 => "0000000001000000001001011000001100",
			1435 => "0000000111000000001111011100001000",
			1436 => "0000001101000000000111111100000100",
			1437 => "00000001000001000001011011000001",
			1438 => "00000000000000000001011011000001",
			1439 => "00000000000000000001011011000001",
			1440 => "0000001101000000000100101000000100",
			1441 => "11111111011101110001011011000001",
			1442 => "0000000111000000001000011000010000",
			1443 => "0000001100000000001000000000001000",
			1444 => "0000001011000000000100010000000100",
			1445 => "00000000101000000001011011000001",
			1446 => "00000000000000000001011011000001",
			1447 => "0000000111000000000001101000000100",
			1448 => "00000000000000000001011011000001",
			1449 => "11111111010001010001011011000001",
			1450 => "0000001011000000000010001000000100",
			1451 => "00000000000000000001011011000001",
			1452 => "0000000001000000001101111100000100",
			1453 => "00000000101001000001011011000001",
			1454 => "00000000000000000001011011000001",
			1455 => "11111110110001110001011011000001",
			1456 => "0000000111000000001101100000000100",
			1457 => "11111110011101010001011101000101",
			1458 => "0000001010000000000111101100010000",
			1459 => "0000000010000000001101000100001100",
			1460 => "0000001011000000001110110000001000",
			1461 => "0000000010000000000100001000000100",
			1462 => "00000000000000000001011101000101",
			1463 => "00000001000011000001011101000101",
			1464 => "11111110110111100001011101000101",
			1465 => "00000001010110110001011101000101",
			1466 => "0000000101000000001110101000001100",
			1467 => "0000001000000000000111110100000100",
			1468 => "00000000000000000001011101000101",
			1469 => "0000001011000000001011011100000100",
			1470 => "11111110100100100001011101000101",
			1471 => "00000000000000000001011101000101",
			1472 => "0000001001000000001100011000000100",
			1473 => "11111110110101000001011101000101",
			1474 => "0000000111000000001000011000010000",
			1475 => "0000001001000000001111000000001000",
			1476 => "0000000011000000001111010100000100",
			1477 => "00000000000100000001011101000101",
			1478 => "00000001100101010001011101000101",
			1479 => "0000001101000000001010001000000100",
			1480 => "11111111011100000001011101000101",
			1481 => "00000000010100000001011101000101",
			1482 => "0000000011000000001000100000001000",
			1483 => "0000001000000000001000100100000100",
			1484 => "00000000000000000001011101000101",
			1485 => "11111110101000100001011101000101",
			1486 => "0000001001000000001010100000000100",
			1487 => "00000001010010000001011101000101",
			1488 => "11111111010000010001011101000101",
			1489 => "0000001010000000001010100101100000",
			1490 => "0000001000000000001000100100110000",
			1491 => "0000000010000000001101000100011100",
			1492 => "0000000001000000000111100100010000",
			1493 => "0000001110000000001010111000001000",
			1494 => "0000000110000000001111001100000100",
			1495 => "00000001000111010001100000110001",
			1496 => "11111110101011110001100000110001",
			1497 => "0000001111000000001011000000000100",
			1498 => "00001100100111110001100000110001",
			1499 => "00000010000000000001100000110001",
			1500 => "0000001000000000000000001000000100",
			1501 => "11111110011100100001100000110001",
			1502 => "0000000110000000000001000100000100",
			1503 => "00000000111101000001100000110001",
			1504 => "11111110111110010001100000110001",
			1505 => "0000000001000000000000111100010000",
			1506 => "0000000111000000001000011000001100",
			1507 => "0000001010000000000000001000000100",
			1508 => "00000001101110100001100000110001",
			1509 => "0000001110000000000110010000000100",
			1510 => "00000000010010100001100000110001",
			1511 => "00000010001011110001100000110001",
			1512 => "00000000001001110001100000110001",
			1513 => "11111110110111000001100000110001",
			1514 => "0000000011000000001010000100100000",
			1515 => "0000001010000000000000001000001000",
			1516 => "0000000010000000000110010000000100",
			1517 => "11111110011001010001100000110001",
			1518 => "00000001110111110001100000110001",
			1519 => "0000000110000000001101111100001000",
			1520 => "0000000001000000001111001100000100",
			1521 => "11111111000110000001100000110001",
			1522 => "00000001110101110001100000110001",
			1523 => "0000001111000000001100010000001000",
			1524 => "0000000101000000000001000000000100",
			1525 => "11111110100001000001100000110001",
			1526 => "00000010000100100001100000110001",
			1527 => "0000000111000000000001101000000100",
			1528 => "11111111110110110001100000110001",
			1529 => "11111101001011110001100000110001",
			1530 => "0000000111000000001111011100001100",
			1531 => "0000001001000000000100111100001000",
			1532 => "0000000011000000000111010100000100",
			1533 => "00000001010110110001100000110001",
			1534 => "00000011000000110001100000110001",
			1535 => "11111111000100000001100000110001",
			1536 => "11111110011110110001100000110001",
			1537 => "0000001010000000000111110100001100",
			1538 => "0000000010000000000110101100000100",
			1539 => "11111110011100110001100000110001",
			1540 => "0000000001000000001110010100000100",
			1541 => "00000011100110000001100000110001",
			1542 => "11111111111001100001100000110001",
			1543 => "0000000101000000001111100100000100",
			1544 => "11111110011010010001100000110001",
			1545 => "0000001111000000001011100100000100",
			1546 => "00000001100100000001100000110001",
			1547 => "11111110100011100001100000110001",
			1548 => "0000000000000000001001101001001100",
			1549 => "0000001110000000001110101000011100",
			1550 => "0000000110000000000001000100011000",
			1551 => "0000000011000000001001001000000100",
			1552 => "11111111000010010001100011111101",
			1553 => "0000001100000000000110000100010000",
			1554 => "0000001100000000001100110000001000",
			1555 => "0000000100000000000111010000000100",
			1556 => "11111111110100010001100011111101",
			1557 => "00000000111000100001100011111101",
			1558 => "0000000001000000000111100100000100",
			1559 => "00000001101100010001100011111101",
			1560 => "00000000000000000001100011111101",
			1561 => "11111111000100000001100011111101",
			1562 => "11111110011010010001100011111101",
			1563 => "0000000110000000001101111100001000",
			1564 => "0000001100000000001000000000000100",
			1565 => "00000001100100100001100011111101",
			1566 => "00000000000000000001100011111101",
			1567 => "0000000011000000001100000000001000",
			1568 => "0000001100000000000100011000000100",
			1569 => "00000000000000000001100011111101",
			1570 => "11111110000100110001100011111101",
			1571 => "0000001100000000001000000000010000",
			1572 => "0000000110000000000100110100001000",
			1573 => "0000001001000000000100111100000100",
			1574 => "00000001101101110001100011111101",
			1575 => "00000000000000000001100011111101",
			1576 => "0000000011000000000111010100000100",
			1577 => "11111111011010000001100011111101",
			1578 => "00000001010001110001100011111101",
			1579 => "0000001101000000001010001000001000",
			1580 => "0000000000000000000101000100000100",
			1581 => "00000001001010110001100011111101",
			1582 => "11111101111000100001100011111101",
			1583 => "0000001100000000001001001000000100",
			1584 => "00000001101101010001100011111101",
			1585 => "00000000000000000001100011111101",
			1586 => "0000000010000000000010110000010000",
			1587 => "0000001000000000000110011100001100",
			1588 => "0000001101000000001111010000000100",
			1589 => "11111110101111110001100011111101",
			1590 => "0000001110000000000110111100000100",
			1591 => "00000000111110000001100011111101",
			1592 => "11111111001011110001100011111101",
			1593 => "11111110011010010001100011111101",
			1594 => "0000001010000000000001010000001000",
			1595 => "0000000110000000000101010000000100",
			1596 => "00000010101110010001100011111101",
			1597 => "00000000000000000001100011111101",
			1598 => "11111110101001000001100011111101",
			1599 => "0000001010000000000010101101000100",
			1600 => "0000000001000000000000111101000000",
			1601 => "0000001110000000001110101000100000",
			1602 => "0000000000000000000110011000011100",
			1603 => "0000001100000000001100110000010000",
			1604 => "0000001111000000001011000000001000",
			1605 => "0000000110000000001111001100000100",
			1606 => "00000001111010110001100110110001",
			1607 => "11111110100110010001100110110001",
			1608 => "0000000001000000000111100100000100",
			1609 => "00000011110011110001100110110001",
			1610 => "00000001001011000001100110110001",
			1611 => "0000000001000000000111100100001000",
			1612 => "0000001100000000000110000100000100",
			1613 => "00000000011000010001100110110001",
			1614 => "00000000000000000001100110110001",
			1615 => "11111110011100010001100110110001",
			1616 => "11111101111110010001100110110001",
			1617 => "0000000011000000001000001100011000",
			1618 => "0000000110000000001101111100001100",
			1619 => "0000001011000000000010001000000100",
			1620 => "00000001110100110001100110110001",
			1621 => "0000001100000000001011000000000100",
			1622 => "00000001001011000001100110110001",
			1623 => "00000000100001100001100110110001",
			1624 => "0000000011000000001100010000000100",
			1625 => "11111100001001000001100110110001",
			1626 => "0000000001000000001001011000000100",
			1627 => "00000001110011000001100110110001",
			1628 => "11111111101111100001100110110001",
			1629 => "0000001011000000000101110100000100",
			1630 => "00000011101111000001100110110001",
			1631 => "00000001011011000001100110110001",
			1632 => "11111110011100110001100110110001",
			1633 => "0000001010000000000011101000001100",
			1634 => "0000000100000000001111101000000100",
			1635 => "11111110011111000001100110110001",
			1636 => "0000001000000000000110011100000100",
			1637 => "00000100000010110001100110110001",
			1638 => "11111111011001100001100110110001",
			1639 => "0000000101000000001111100100000100",
			1640 => "11111110011000110001100110110001",
			1641 => "0000001011000000000111111100000100",
			1642 => "00000001010110010001100110110001",
			1643 => "11111110011110110001100110110001",
			1644 => "0000000000000000001100000101011000",
			1645 => "0000001000000000000111110100011100",
			1646 => "0000000010000000001101000100010100",
			1647 => "0000000111000000001100101000010000",
			1648 => "0000001110000000000100001000000100",
			1649 => "11111111101111010001101010010101",
			1650 => "0000001001000000000000111100000100",
			1651 => "00000010000010000001101010010101",
			1652 => "0000001101000000000100000100000100",
			1653 => "11111110110100100001101010010101",
			1654 => "00000001100000000001101010010101",
			1655 => "11111110010001000001101010010101",
			1656 => "0000000110000000001101111100000100",
			1657 => "00000001100011110001101010010101",
			1658 => "00000000000000000001101010010101",
			1659 => "0000000011000000001110110100001100",
			1660 => "0000001011000000000101100100001000",
			1661 => "0000000010000000000011001000000100",
			1662 => "11111110100001010001101010010101",
			1663 => "00000000000000000001101010010101",
			1664 => "11111100111100110001101010010101",
			1665 => "0000000010000000001110110100010000",
			1666 => "0000001010000000000000001000001000",
			1667 => "0000001001000000000100111100000100",
			1668 => "00000001110001000001101010010101",
			1669 => "00000000000000000001101010010101",
			1670 => "0000000011000000000110111100000100",
			1671 => "11111110110110000001101010010101",
			1672 => "00000000000000000001101010010101",
			1673 => "0000000011000000001010000100010000",
			1674 => "0000001011000000000110110100001000",
			1675 => "0000001001000000001111000000000100",
			1676 => "00000000101011000001101010010101",
			1677 => "00000000000000000001101010010101",
			1678 => "0000000000000000000001010100000100",
			1679 => "11111110000101010001101010010101",
			1680 => "00000000000000000001101010010101",
			1681 => "0000001101000000001001011100001000",
			1682 => "0000000000000000000001110000000100",
			1683 => "00000010000111000001101010010101",
			1684 => "11111111101011110001101010010101",
			1685 => "0000000010000000000110111100000100",
			1686 => "11111110111010000001101010010101",
			1687 => "00000001001011000001101010010101",
			1688 => "0000000010000000000010110000010000",
			1689 => "0000001010000000000011101000001100",
			1690 => "0000000100000000001101101100000100",
			1691 => "11111110110010110001101010010101",
			1692 => "0000000101000000001101000100000100",
			1693 => "00000000000000000001101010010101",
			1694 => "00000000101111010001101010010101",
			1695 => "11111110011010010001101010010101",
			1696 => "0000000110000000001000010000000100",
			1697 => "00000010101010100001101010010101",
			1698 => "0000001000000000001001101000000100",
			1699 => "00000000000000000001101010010101",
			1700 => "11111110101100000001101010010101",
			1701 => "0000000000000000001100000101010000",
			1702 => "0000001000000000000111110100011000",
			1703 => "0000001110000000000100001000000100",
			1704 => "11111111001001110001101101100001",
			1705 => "0000000001000000000000111100010000",
			1706 => "0000000001000000000110101000000100",
			1707 => "00000010100100010001101101100001",
			1708 => "0000001011000000000100001000000100",
			1709 => "11111110110010100001101101100001",
			1710 => "0000001111000000000010001000000100",
			1711 => "00000000010101100001101101100001",
			1712 => "00000001100110010001101101100001",
			1713 => "11111111100110100001101101100001",
			1714 => "0000000011000000001100010000001000",
			1715 => "0000000100000000001100000000000100",
			1716 => "11111101110110100001101101100001",
			1717 => "00000000000000000001101101100001",
			1718 => "0000001100000000001000000000100000",
			1719 => "0000001111000000000111011000010000",
			1720 => "0000001000000000001000100100001000",
			1721 => "0000000011000000001100000000000100",
			1722 => "00000000000000000001101101100001",
			1723 => "00000001100110110001101101100001",
			1724 => "0000001110000000000010000100000100",
			1725 => "00000000000000000001101101100001",
			1726 => "11111110101110010001101101100001",
			1727 => "0000000000000000000001110000001000",
			1728 => "0000001011000000000010001000000100",
			1729 => "00000000110001110001101101100001",
			1730 => "00000010110011100001101101100001",
			1731 => "0000001100000000001011000000000100",
			1732 => "00000000001001100001101101100001",
			1733 => "00000000000000000001101101100001",
			1734 => "0000000000000000000101000100000100",
			1735 => "00000001011100110001101101100001",
			1736 => "0000000101000000001001010000000100",
			1737 => "11111101010110110001101101100001",
			1738 => "0000001100000000001001001000000100",
			1739 => "00000001101100100001101101100001",
			1740 => "11111111000110110001101101100001",
			1741 => "0000000001000000001111001100000100",
			1742 => "11111110011000110001101101100001",
			1743 => "0000001001000000000100111100001100",
			1744 => "0000001101000000001111010000000100",
			1745 => "11111110111101000001101101100001",
			1746 => "0000000011000000000010010100000100",
			1747 => "00000010100000110001101101100001",
			1748 => "11111111101110000001101101100001",
			1749 => "0000000101000000000000010000000100",
			1750 => "11111110011011100001101101100001",
			1751 => "00000001111001100001101101100001",
			1752 => "0000000000000000001100000101011000",
			1753 => "0000001100000000001000000000110100",
			1754 => "0000001111000000001100100100010100",
			1755 => "0000000110000000000001000100010000",
			1756 => "0000001100000000000110000100001100",
			1757 => "0000001110000000000100001000000100",
			1758 => "11111111110100000001110001000101",
			1759 => "0000001001000000000000111100000100",
			1760 => "00000001101011000001110001000101",
			1761 => "00000000011100000001110001000101",
			1762 => "11111111001100110001110001000101",
			1763 => "11111110010001010001110001000101",
			1764 => "0000001001000000001111000000000100",
			1765 => "00000001100011000001110001000101",
			1766 => "0000000111000000001000011000010000",
			1767 => "0000001100000000001011000000001000",
			1768 => "0000000101000000001110101000000100",
			1769 => "11111111010001110001110001000101",
			1770 => "00000001001110110001110001000101",
			1771 => "0000001010000000000000001000000100",
			1772 => "11111111111001110001110001000101",
			1773 => "11111110011001000001110001000101",
			1774 => "0000000111000000001000011000001000",
			1775 => "0000001001000000000100111100000100",
			1776 => "00000001111101000001110001000101",
			1777 => "00000000000000000001110001000101",
			1778 => "11111111110011100001110001000101",
			1779 => "0000001110000000001010001000000100",
			1780 => "11111110000111000001110001000101",
			1781 => "0000001111000000001100010000001000",
			1782 => "0000001010000000000000001000000100",
			1783 => "00000001100010010001110001000101",
			1784 => "00000000000000000001110001000101",
			1785 => "0000001100000000001000000000001000",
			1786 => "0000001000000000001000100100000100",
			1787 => "00000001000110010001110001000101",
			1788 => "00000000000000000001110001000101",
			1789 => "0000001000000000001000010100001000",
			1790 => "0000001100000000001001110100000100",
			1791 => "11111110001111010001110001000101",
			1792 => "00000000000000000001110001000101",
			1793 => "0000001100000000001001110100000100",
			1794 => "00000001001000100001110001000101",
			1795 => "00000000000000000001110001000101",
			1796 => "0000001111000000000110001100010000",
			1797 => "0000001010000000000011101000001100",
			1798 => "0000000100000000001101101100000100",
			1799 => "11111110110111110001110001000101",
			1800 => "0000000101000000001101000100000100",
			1801 => "00000000000000000001110001000101",
			1802 => "00000000100101010001110001000101",
			1803 => "11111110011010110001110001000101",
			1804 => "0000000110000000000101010000001000",
			1805 => "0000000000000000001101010000000100",
			1806 => "00000000000000000001110001000101",
			1807 => "00000010001111100001110001000101",
			1808 => "11111110110001000001110001000101",
			1809 => "0000000101000000001110110000000100",
			1810 => "11111110011110000001110011110001",
			1811 => "0000000000000000000001010100110100",
			1812 => "0000000011000000000110111100101100",
			1813 => "0000001100000000000100011000011000",
			1814 => "0000001111000000001100100100001100",
			1815 => "0000000110000000000001000100001000",
			1816 => "0000001011000000000100001000000100",
			1817 => "00000000000000000001110011110001",
			1818 => "00000000111100000001110011110001",
			1819 => "11111110111111000001110011110001",
			1820 => "0000000110000000000100110100001000",
			1821 => "0000001001000000000100111100000100",
			1822 => "00000001011000110001110011110001",
			1823 => "00000000000000000001110011110001",
			1824 => "00000000000000000001110011110001",
			1825 => "0000000110000000001101111100000100",
			1826 => "00000000100001100001110011110001",
			1827 => "0000000101000000001100100100001000",
			1828 => "0000001001000000001001100100000100",
			1829 => "00000000000000000001110011110001",
			1830 => "11111110011000000001110011110001",
			1831 => "0000000000000000000101000100000100",
			1832 => "00000000110100000001110011110001",
			1833 => "11111110111010010001110011110001",
			1834 => "0000000101000000001110000100000100",
			1835 => "00000000000000000001110011110001",
			1836 => "00000001011110110001110011110001",
			1837 => "0000000011000000001000001100001000",
			1838 => "0000001111000000000000010000000100",
			1839 => "11111110111000100001110011110001",
			1840 => "00000000000000000001110011110001",
			1841 => "0000000110000000001011001100001100",
			1842 => "0000001001000000001000010000001000",
			1843 => "0000000101000000000010011100000100",
			1844 => "00000001110110110001110011110001",
			1845 => "00000000000000000001110011110001",
			1846 => "00000000000000000001110011110001",
			1847 => "0000001101000000000011000000000100",
			1848 => "11111110110100100001110011110001",
			1849 => "0000000000000000001010111000000100",
			1850 => "00000000111001010001110011110001",
			1851 => "00000000000000000001110011110001",
			1852 => "0000000111000000001101100000000100",
			1853 => "11111110100000000001110110110101",
			1854 => "0000000111000000001000011000111000",
			1855 => "0000001010000000000000001000100100",
			1856 => "0000000011000000001100010000011100",
			1857 => "0000001000000000000111110100010000",
			1858 => "0000000010000000001101000100001000",
			1859 => "0000001001000000000000111100000100",
			1860 => "00000000111111100001110110110101",
			1861 => "11111111101100110001110110110101",
			1862 => "0000001001000000001001100100000100",
			1863 => "00000001001101110001110110110101",
			1864 => "00000000000000000001110110110101",
			1865 => "0000000000000000000110011100000100",
			1866 => "00000000000000000001110110110101",
			1867 => "0000001101000000000010011100000100",
			1868 => "11111110110110100001110110110101",
			1869 => "00000000000000000001110110110101",
			1870 => "0000001001000000000100111100000100",
			1871 => "00000001001010100001110110110101",
			1872 => "00000000000000000001110110110101",
			1873 => "0000000011000000001010000100001000",
			1874 => "0000001111000000001010000100000100",
			1875 => "11111110111000000001110110110101",
			1876 => "00000000000000000001110110110101",
			1877 => "0000000010000000001100000000000100",
			1878 => "00000000101010110001110110110101",
			1879 => "0000001100000000000100011000000100",
			1880 => "11111111001100010001110110110101",
			1881 => "00000000000000000001110110110101",
			1882 => "0000000111000000001111011100010000",
			1883 => "0000001001000000001000010000001100",
			1884 => "0000000010000000000110010000000100",
			1885 => "00000000000000000001110110110101",
			1886 => "0000001101000000000101110000000100",
			1887 => "00000000000000000001110110110101",
			1888 => "00000001010011000001110110110101",
			1889 => "11111111111101100001110110110101",
			1890 => "0000001101000000001100010100001000",
			1891 => "0000001100000000001011000000000100",
			1892 => "00000000000000000001110110110101",
			1893 => "11111111010000000001110110110101",
			1894 => "0000001001000000001010100000001100",
			1895 => "0000001000000000001001101000001000",
			1896 => "0000000110000000000101010000000100",
			1897 => "00000000110100010001110110110101",
			1898 => "00000000000000000001110110110101",
			1899 => "00000000000000000001110110110101",
			1900 => "11111111110010110001110110110101",
			1901 => "0000000111000000001101100000000100",
			1902 => "11111110110100110001111001010011",
			1903 => "0000001010000000000111101100001000",
			1904 => "0000001110000000000100001000000100",
			1905 => "00000000000000000001111001010011",
			1906 => "00000000110010010001111001010011",
			1907 => "0000000011000000001010000100101000",
			1908 => "0000000011000000001100010000010000",
			1909 => "0000000000000000001100011100000100",
			1910 => "00000000000000000001111001010011",
			1911 => "0000000111000000000001101000001000",
			1912 => "0000001101000000000010011100000100",
			1913 => "11111110111101010001111001010011",
			1914 => "00000000000000000001111001010011",
			1915 => "00000000000000000001111001010011",
			1916 => "0000001101000000000111111100001100",
			1917 => "0000000001000000000000111100001000",
			1918 => "0000000111000000001111011100000100",
			1919 => "00000000110001110001111001010011",
			1920 => "00000000000000000001111001010011",
			1921 => "00000000000000000001111001010011",
			1922 => "0000000111000000001111011100001000",
			1923 => "0000001100000000001001001000000100",
			1924 => "11111110110100000001111001010011",
			1925 => "00000000000000000001111001010011",
			1926 => "00000000000000000001111001010011",
			1927 => "0000001100000000000100011000000100",
			1928 => "11111111111001100001111001010011",
			1929 => "0000001001000000000100111100001000",
			1930 => "0000000111000000001111011100000100",
			1931 => "00000001000110000001111001010011",
			1932 => "00000000000000000001111001010011",
			1933 => "0000000011000000001000100000001000",
			1934 => "0000000111000000000001101000000100",
			1935 => "00000000000000000001111001010011",
			1936 => "11111111101111100001111001010011",
			1937 => "0000000001000000001101111100000100",
			1938 => "00000000100011100001111001010011",
			1939 => "00000000000000000001111001010011",
			1940 => "00000000000000000001111001010101",
			1941 => "00000000000000000001111001011001",
			1942 => "00000000000000000001111001011101",
			1943 => "00000000000000000001111001100001",
			1944 => "00000000000000000001111001100101",
			1945 => "00000000000000000001111001101001",
			1946 => "00000000000000000001111001101101",
			1947 => "00000000000000000001111001110001",
			1948 => "0000001100000000001100110000000100",
			1949 => "00000000000000000001111010000101",
			1950 => "0000001100000000000001101000000100",
			1951 => "11111111111011110001111010000101",
			1952 => "00000000000000000001111010000101",
			1953 => "0000000011000000000111010100001000",
			1954 => "0000000011000000001101010100000100",
			1955 => "00000000000000000001111010100001",
			1956 => "11111111111001100001111010100001",
			1957 => "0000000011000000000010100100000100",
			1958 => "00000000000001010001111010100001",
			1959 => "00000000000000000001111010100001",
			1960 => "0000000000000000000001010100001100",
			1961 => "0000000111000000001101100000000100",
			1962 => "00000000000000000001111010111101",
			1963 => "0000000100000000000111001000000100",
			1964 => "00000000000000000001111010111101",
			1965 => "00000000000100110001111010111101",
			1966 => "00000000000000000001111010111101",
			1967 => "0000000011000000000111010100001100",
			1968 => "0000001001000000000000111100000100",
			1969 => "00000000000000000001111011011001",
			1970 => "0000000010000000001010000100000100",
			1971 => "11111111101111110001111011011001",
			1972 => "00000000000000000001111011011001",
			1973 => "00000000000000000001111011011001",
			1974 => "0000000101000000001111010000001100",
			1975 => "0000000111000000000001101000000100",
			1976 => "00000000000000000001111011111101",
			1977 => "0000000101000000001101000100000100",
			1978 => "00000000000000000001111011111101",
			1979 => "11111111110100010001111011111101",
			1980 => "0000000111000000000001001000000100",
			1981 => "00000000001010010001111011111101",
			1982 => "00000000000000000001111011111101",
			1983 => "0000001001000000000101011100001100",
			1984 => "0000001110000000000100001000000100",
			1985 => "00000000000000000001111100100001",
			1986 => "0000000000000000001100011100000100",
			1987 => "00000000000011110001111100100001",
			1988 => "00000000000000000001111100100001",
			1989 => "0000000110000000001101111100000100",
			1990 => "11111111101110100001111100100001",
			1991 => "00000000000000000001111100100001",
			1992 => "0000001011000000000101100100001100",
			1993 => "0000001100000000001100110000000100",
			1994 => "00000000000000000001111101001101",
			1995 => "0000001100000000001000000000000100",
			1996 => "11111111111001100001111101001101",
			1997 => "00000000000000000001111101001101",
			1998 => "0000000001000000000000111100001000",
			1999 => "0000000111000000000111010000000100",
			2000 => "00000000010000100001111101001101",
			2001 => "00000000000000000001111101001101",
			2002 => "00000000000000000001111101001101",
			2003 => "0000000011000000001010000100001100",
			2004 => "0000000111000000000001101000001000",
			2005 => "0000000111000000000110000100000100",
			2006 => "00000000000000000001111101111001",
			2007 => "00000000000000110001111101111001",
			2008 => "11111111110110010001111101111001",
			2009 => "0000000111000000001000011000000100",
			2010 => "00000000000000000001111101111001",
			2011 => "0000000111000000001111011100000100",
			2012 => "00000000000010110001111101111001",
			2013 => "00000000000000000001111101111001",
			2014 => "0000001010000000000010101100010000",
			2015 => "0000001110000000001110101000000100",
			2016 => "00000000000000000001111110011101",
			2017 => "0000001011000000000101110100001000",
			2018 => "0000000001000000000000111100000100",
			2019 => "00000000010110110001111110011101",
			2020 => "00000000000000000001111110011101",
			2021 => "00000000000000000001111110011101",
			2022 => "00000000000000000001111110011101",
			2023 => "0000001011000000000100010000010000",
			2024 => "0000001011000000001000011000000100",
			2025 => "00000000000000000001111111000001",
			2026 => "0000000001000000000000111100001000",
			2027 => "0000000001000000001111001100000100",
			2028 => "00000000000000000001111111000001",
			2029 => "00000000001011010001111111000001",
			2030 => "00000000000000000001111111000001",
			2031 => "00000000000000000001111111000001",
			2032 => "0000000000000000000001010100010000",
			2033 => "0000000001000000000000111100001100",
			2034 => "0000000111000000001101100000000100",
			2035 => "00000000000000000001111111100101",
			2036 => "0000000100000000000111001000000100",
			2037 => "00000000000000000001111111100101",
			2038 => "00000000000111100001111111100101",
			2039 => "00000000000000000001111111100101",
			2040 => "00000000000000000001111111100101",
			2041 => "0000000110000000000100110100010000",
			2042 => "0000001010000000001010100000001100",
			2043 => "0000000110000000000111101000000100",
			2044 => "00000000000000000010000000010001",
			2045 => "0000001010000000000000001000000100",
			2046 => "00000000010001000010000000010001",
			2047 => "00000000000000000010000000010001",
			2048 => "00000000000000000010000000010001",
			2049 => "0000001010000000000000001000000100",
			2050 => "00000000000000000010000000010001",
			2051 => "11111111110111100010000000010001",
			2052 => "0000001110000000000110100100000100",
			2053 => "11111111010111100010000000111101",
			2054 => "0000000101000000001111010000001100",
			2055 => "0000000101000000000100000100000100",
			2056 => "00000000000000000010000000111101",
			2057 => "0000000101000000000101001000000100",
			2058 => "11111111110110100010000000111101",
			2059 => "00000000000000000010000000111101",
			2060 => "0000000101000000001111100100000100",
			2061 => "00000000000001110010000000111101",
			2062 => "00000000000000000010000000111101",
			2063 => "0000000000000000000110011100010000",
			2064 => "0000001101000000001010011100001100",
			2065 => "0000000100000000000111001000000100",
			2066 => "00000000000000000010000001110001",
			2067 => "0000000111000000001110001100000100",
			2068 => "00000000001000000010000001110001",
			2069 => "00000000000000000010000001110001",
			2070 => "00000000000000000010000001110001",
			2071 => "0000000111000000001000011000001000",
			2072 => "0000001101000000001110010000000100",
			2073 => "11111111110101100010000001110001",
			2074 => "00000000000000000010000001110001",
			2075 => "00000000000000000010000001110001",
			2076 => "0000000110000000000100110100010000",
			2077 => "0000001010000000001010100000001100",
			2078 => "0000000010000000000111100000000100",
			2079 => "00000000000000000010000010100101",
			2080 => "0000001010000000000000001000000100",
			2081 => "00000000010101000010000010100101",
			2082 => "00000000000000000010000010100101",
			2083 => "00000000000000000010000010100101",
			2084 => "0000000010000000001110111000001000",
			2085 => "0000001010000000000000001000000100",
			2086 => "00000000000000000010000010100101",
			2087 => "11111111110011100010000010100101",
			2088 => "00000000000000000010000010100101",
			2089 => "0000000101000000001110010000010100",
			2090 => "0000001000000000000111110100001100",
			2091 => "0000001010000000000100111100000100",
			2092 => "11111111111011110010000011100001",
			2093 => "0000000000000000000110011100000100",
			2094 => "00000000000011010010000011100001",
			2095 => "00000000000000000010000011100001",
			2096 => "0000001010000000000111101100000100",
			2097 => "00000000000000000010000011100001",
			2098 => "11111111101100110010000011100001",
			2099 => "0000000110000000001000010000001000",
			2100 => "0000000001000000001101111100000100",
			2101 => "00000000000110010010000011100001",
			2102 => "00000000000000000010000011100001",
			2103 => "00000000000000000010000011100001",
			2104 => "0000001110000000000110100100001000",
			2105 => "0000000110000000001101011100000100",
			2106 => "00000000000000000010000100010101",
			2107 => "11111111110011100010000100010101",
			2108 => "0000001010000000000000001000010000",
			2109 => "0000000110000000000100110100001100",
			2110 => "0000001001000000000100111100001000",
			2111 => "0000001111000000001010011100000100",
			2112 => "00000000000000000010000100010101",
			2113 => "00000000010111100010000100010101",
			2114 => "00000000000000000010000100010101",
			2115 => "00000000000000000010000100010101",
			2116 => "00000000000000000010000100010101",
			2117 => "0000001110000000001110101000001000",
			2118 => "0000001000000000001001111100000100",
			2119 => "00000000000000000010000101001001",
			2120 => "11111111110101010010000101001001",
			2121 => "0000000001000000000101011100010000",
			2122 => "0000000111000000000111010000001100",
			2123 => "0000000110000000001010011000001000",
			2124 => "0000001100000000000110000100000100",
			2125 => "00000000000000000010000101001001",
			2126 => "00000000011000000010000101001001",
			2127 => "00000000000000000010000101001001",
			2128 => "00000000000000000010000101001001",
			2129 => "00000000000000000010000101001001",
			2130 => "0000000000000000000001010100010100",
			2131 => "0000000001000000000000111100010000",
			2132 => "0000000111000000001101100000000100",
			2133 => "00000000000000000010000101110101",
			2134 => "0000001100000000001000000000001000",
			2135 => "0000000100000000000111001000000100",
			2136 => "00000000000000000010000101110101",
			2137 => "00000000001001100010000101110101",
			2138 => "00000000000000000010000101110101",
			2139 => "00000000000000000010000101110101",
			2140 => "00000000000000000010000101110101",
			2141 => "0000001100000000001100110000001100",
			2142 => "0000000000000000001010110000001000",
			2143 => "0000000010000000000100001000000100",
			2144 => "00000000000000000010000110111001",
			2145 => "00000000010101010010000110111001",
			2146 => "00000000000000000010000110111001",
			2147 => "0000000111000000001000000000001100",
			2148 => "0000001100000000001100110000000100",
			2149 => "00000000000000000010000110111001",
			2150 => "0000001100000000000100011000000100",
			2151 => "11111111101010000010000110111001",
			2152 => "00000000000000000010000110111001",
			2153 => "0000000110000000000100110100001000",
			2154 => "0000001100000000001000000000000100",
			2155 => "00000000001011100010000110111001",
			2156 => "00000000000000000010000110111001",
			2157 => "00000000000000000010000110111001",
			2158 => "0000000011000000001100010000011000",
			2159 => "0000001001000000000000111100001100",
			2160 => "0000001110000000000100001000000100",
			2161 => "00000000000000000010001000000101",
			2162 => "0000000000000000000101000100000100",
			2163 => "00000000001001110010001000000101",
			2164 => "00000000000000000010001000000101",
			2165 => "0000000001000000000110101000000100",
			2166 => "00000000000000000010001000000101",
			2167 => "0000001101000000000010011100000100",
			2168 => "11111111101101110010001000000101",
			2169 => "00000000000000000010001000000101",
			2170 => "0000001010000000000001010000001100",
			2171 => "0000000101000000001110101000000100",
			2172 => "00000000000000000010001000000101",
			2173 => "0000000001000000001101111100000100",
			2174 => "00000000001010110010001000000101",
			2175 => "00000000000000000010001000000101",
			2176 => "00000000000000000010001000000101",
			2177 => "0000001100000000001100110000001100",
			2178 => "0000000010000000001101000100001000",
			2179 => "0000001110000000000100001000000100",
			2180 => "00000000000000000010001001010001",
			2181 => "00000000011000100010001001010001",
			2182 => "00000000000000000010001001010001",
			2183 => "0000000011000000001010000100010000",
			2184 => "0000001100000000001001110100001100",
			2185 => "0000000010000000001010000100001000",
			2186 => "0000001110000000001100010000000100",
			2187 => "11111111100111100010001001010001",
			2188 => "00000000000000000010001001010001",
			2189 => "00000000000000000010001001010001",
			2190 => "00000000000000000010001001010001",
			2191 => "0000001001000000001000010000001000",
			2192 => "0000000010000000001101001000000100",
			2193 => "00000000010001100010001001010001",
			2194 => "00000000000000000010001001010001",
			2195 => "00000000000000000010001001010001",
			2196 => "0000001001000000001100011000001100",
			2197 => "0000001001000000000000111100000100",
			2198 => "00000000000000000010001010011101",
			2199 => "0000000001000000000110101000000100",
			2200 => "00000000000000000010001010011101",
			2201 => "11111111110111000010001010011101",
			2202 => "0000000100000000000110111100001100",
			2203 => "0000001100000000000100011000000100",
			2204 => "00000000000000000010001010011101",
			2205 => "0000001100000000001001001000000100",
			2206 => "11111111110111110010001010011101",
			2207 => "00000000000000000010001010011101",
			2208 => "0000000001000000000000111100001100",
			2209 => "0000001100000000001001110100001000",
			2210 => "0000001100000000000111001000000100",
			2211 => "00000000000000000010001010011101",
			2212 => "00000000010110000010001010011101",
			2213 => "00000000000000000010001010011101",
			2214 => "00000000000000000010001010011101",
			2215 => "0000000101000000000111100000011100",
			2216 => "0000000000000000000110011100001100",
			2217 => "0000001111000000001010011100000100",
			2218 => "11111111111110000010001011110001",
			2219 => "0000000011000000001001010100000100",
			2220 => "00000000001100110010001011110001",
			2221 => "00000000000000000010001011110001",
			2222 => "0000001011000000000010001000001100",
			2223 => "0000001010000000000111101100000100",
			2224 => "00000000000000000010001011110001",
			2225 => "0000001100000000001001110100000100",
			2226 => "11111111001011000010001011110001",
			2227 => "00000000000000000010001011110001",
			2228 => "00000000000000000010001011110001",
			2229 => "0000000110000000001000010000001100",
			2230 => "0000000001000000001101111100001000",
			2231 => "0000001011000000000101100100000100",
			2232 => "00000000000000000010001011110001",
			2233 => "00000000011100110010001011110001",
			2234 => "00000000000000000010001011110001",
			2235 => "00000000000000000010001011110001",
			2236 => "0000000011000000001100010000011000",
			2237 => "0000001001000000000000111100001100",
			2238 => "0000001110000000000100001000000100",
			2239 => "00000000000000000010001101000101",
			2240 => "0000000000000000000101000100000100",
			2241 => "00000000001000110010001101000101",
			2242 => "00000000000000000010001101000101",
			2243 => "0000000111000000000101101100000100",
			2244 => "00000000000000000010001101000101",
			2245 => "0000001101000000000010011100000100",
			2246 => "11111111101111100010001101000101",
			2247 => "00000000000000000010001101000101",
			2248 => "0000001010000000000001010000010000",
			2249 => "0000001001000000001010100000001100",
			2250 => "0000001101000000001111010000000100",
			2251 => "00000000000000000010001101000101",
			2252 => "0000001110000000001100010100000100",
			2253 => "00000000000000000010001101000101",
			2254 => "00000000001001100010001101000101",
			2255 => "00000000000000000010001101000101",
			2256 => "00000000000000000010001101000101",
			2257 => "0000001001000000001100011000010100",
			2258 => "0000000110000000001101011100000100",
			2259 => "00000000000000000010001110010001",
			2260 => "0000000101000000000110100100000100",
			2261 => "11111111010101000010001110010001",
			2262 => "0000000111000000001100101000001000",
			2263 => "0000000111000000000110000100000100",
			2264 => "00000000000000000010001110010001",
			2265 => "00000000000110100010001110010001",
			2266 => "11111111111001100010001110010001",
			2267 => "0000000001000000000000111100010000",
			2268 => "0000000111000000001111011100001100",
			2269 => "0000000111000000000001111100000100",
			2270 => "00000000000000000010001110010001",
			2271 => "0000000110000000001011001100000100",
			2272 => "00000000011110100010001110010001",
			2273 => "00000000000000000010001110010001",
			2274 => "00000000000000000010001110010001",
			2275 => "00000000000000000010001110010001",
			2276 => "0000000101000000001111010000011000",
			2277 => "0000000000000000000101000100010000",
			2278 => "0000001100000000001100110000001100",
			2279 => "0000000000000000000110011000001000",
			2280 => "0000001100000000001100110000000100",
			2281 => "00000000000100110010001111100101",
			2282 => "00000000000000000010001111100101",
			2283 => "00000000000000000010001111100101",
			2284 => "00000000000000000010001111100101",
			2285 => "0000001000000000001000100100000100",
			2286 => "00000000000000000010001111100101",
			2287 => "11111111111100000010001111100101",
			2288 => "0000000110000000000101010000010000",
			2289 => "0000001100000000001011000000000100",
			2290 => "00000000000000000010001111100101",
			2291 => "0000000001000000001101011100000100",
			2292 => "00000000000000000010001111100101",
			2293 => "0000000001000000001101111100000100",
			2294 => "00000000001111000010001111100101",
			2295 => "00000000000000000010001111100101",
			2296 => "00000000000000000010001111100101",
			2297 => "0000001000000000001001101000011000",
			2298 => "0000001110000000000100001000000100",
			2299 => "00000000000000000010010000011001",
			2300 => "0000001001000000001111000000010000",
			2301 => "0000000111000000001000011000001100",
			2302 => "0000000111000000001101100000000100",
			2303 => "00000000000000000010010000011001",
			2304 => "0000000110000000001011001100000100",
			2305 => "00000000000111110010010000011001",
			2306 => "00000000000000000010010000011001",
			2307 => "00000000000000000010010000011001",
			2308 => "00000000000000000010010000011001",
			2309 => "00000000000000000010010000011001",
			2310 => "0000000000000000000001010100100000",
			2311 => "0000001111000000000000011100001100",
			2312 => "0000000001000000000110101000001000",
			2313 => "0000001110000000000100001000000100",
			2314 => "00000000000000000010010001100101",
			2315 => "00000000010001110010010001100101",
			2316 => "11111111000011010010010001100101",
			2317 => "0000001100000000001000000000010000",
			2318 => "0000000110000000000100110100001100",
			2319 => "0000000001000000000000111100001000",
			2320 => "0000001010000000000100111100000100",
			2321 => "00000000000000000010010001100101",
			2322 => "00000000011001110010010001100101",
			2323 => "00000000000000000010010001100101",
			2324 => "00000000000000000010010001100101",
			2325 => "00000000000000000010010001100101",
			2326 => "0000000110000000001101111100000100",
			2327 => "00000000000000000010010001100101",
			2328 => "11111111100001000010010001100101",
			2329 => "0000000101000000001100100100011100",
			2330 => "0000000000000000000110011100001100",
			2331 => "0000001111000000001010011100000100",
			2332 => "00000000000000000010010011000001",
			2333 => "0000000010000000001010010100000100",
			2334 => "00000000000110100010010011000001",
			2335 => "00000000000000000010010011000001",
			2336 => "0000001111000000001100010000001100",
			2337 => "0000001101000000000101110000001000",
			2338 => "0000001000000000000111110100000100",
			2339 => "00000000000000000010010011000001",
			2340 => "11111111001000110010010011000001",
			2341 => "00000000000000000010010011000001",
			2342 => "00000000000000000010010011000001",
			2343 => "0000000110000000001000010000010000",
			2344 => "0000000101000000000111100000000100",
			2345 => "00000000000000000010010011000001",
			2346 => "0000000001000000001101111100001000",
			2347 => "0000001011000000000101100100000100",
			2348 => "00000000000000000010010011000001",
			2349 => "00000000011001110010010011000001",
			2350 => "00000000000000000010010011000001",
			2351 => "00000000000000000010010011000001",
			2352 => "0000000011000000001100010000011000",
			2353 => "0000001001000000000000111100001100",
			2354 => "0000000100000000000110110100001000",
			2355 => "0000001110000000000100001000000100",
			2356 => "00000000000000000010010100011101",
			2357 => "00000000001100010010010100011101",
			2358 => "00000000000000000010010100011101",
			2359 => "0000001100000000001100110000000100",
			2360 => "00000000000000000010010100011101",
			2361 => "0000001110000000001010001000000100",
			2362 => "11111111101001110010010100011101",
			2363 => "00000000000000000010010100011101",
			2364 => "0000001001000000001100011000000100",
			2365 => "00000000000000000010010100011101",
			2366 => "0000001001000000001010100000010000",
			2367 => "0000001010000000000001010000001100",
			2368 => "0000001101000000001111010000000100",
			2369 => "00000000000000000010010100011101",
			2370 => "0000001100000000000111001000000100",
			2371 => "00000000000000000010010100011101",
			2372 => "00000000001111000010010100011101",
			2373 => "00000000000000000010010100011101",
			2374 => "00000000000000000010010100011101",
			2375 => "0000001001000000001100011000001000",
			2376 => "0000001001000000000000111100000100",
			2377 => "00000000000000000010010101110001",
			2378 => "11111111111001110010010101110001",
			2379 => "0000000100000000000110111100010100",
			2380 => "0000001100000000000100011000000100",
			2381 => "00000000000000000010010101110001",
			2382 => "0000001100000000001001001000001100",
			2383 => "0000001001000000001001100100000100",
			2384 => "00000000000000000010010101110001",
			2385 => "0000001010000000000111101100000100",
			2386 => "00000000000000000010010101110001",
			2387 => "11111111101111110010010101110001",
			2388 => "00000000000000000010010101110001",
			2389 => "0000001010000000000001010000001100",
			2390 => "0000001100000000000111001000000100",
			2391 => "00000000000000000010010101110001",
			2392 => "0000001001000000001010100000000100",
			2393 => "00000000001101010010010101110001",
			2394 => "00000000000000000010010101110001",
			2395 => "00000000000000000010010101110001",
			2396 => "0000001010000000000000001000011000",
			2397 => "0000001001000000000101011100010000",
			2398 => "0000000001000000000110101000001100",
			2399 => "0000000010000000000100001000000100",
			2400 => "00000000000000000010010111011101",
			2401 => "0000000000000000000011101000000100",
			2402 => "00000000011001000010010111011101",
			2403 => "00000000000000000010010111011101",
			2404 => "00000000000000000010010111011101",
			2405 => "0000000010000000001101000100000100",
			2406 => "11111111111101100010010111011101",
			2407 => "00000000000001100010010111011101",
			2408 => "0000000011000000001010000100001100",
			2409 => "0000001111000000001111010100001000",
			2410 => "0000000001000000000000111100000100",
			2411 => "11111111101111110010010111011101",
			2412 => "00000000000000000010010111011101",
			2413 => "00000000000000000010010111011101",
			2414 => "0000001100000000001011000000000100",
			2415 => "00000000000000000010010111011101",
			2416 => "0000000101000000000010011100001100",
			2417 => "0000000001000000000000111100001000",
			2418 => "0000000111000000001111011100000100",
			2419 => "00000000010100100010010111011101",
			2420 => "00000000000000000010010111011101",
			2421 => "00000000000000000010010111011101",
			2422 => "00000000000000000010010111011101",
			2423 => "0000001110000000001100010000100000",
			2424 => "0000001100000000000100011000010100",
			2425 => "0000001100000000000110000100000100",
			2426 => "00000000000000000010011001000001",
			2427 => "0000001001000000000100111100001100",
			2428 => "0000001001000000001001011000000100",
			2429 => "00000000000000000010011001000001",
			2430 => "0000000000000000000110001000000100",
			2431 => "00000000010100110010011001000001",
			2432 => "00000000000000000010011001000001",
			2433 => "00000000000000000010011001000001",
			2434 => "0000000111000000000001101000000100",
			2435 => "00000000000000000010011001000001",
			2436 => "0000000000000000000110011100000100",
			2437 => "00000000000000000010011001000001",
			2438 => "11111111101011110010011001000001",
			2439 => "0000001011000000000101100100000100",
			2440 => "00000000000000000010011001000001",
			2441 => "0000001010000000000001010000001100",
			2442 => "0000000001000000001101111100001000",
			2443 => "0000000101000000000111100000000100",
			2444 => "00000000000000000010011001000001",
			2445 => "00000000010000010010011001000001",
			2446 => "00000000000000000010011001000001",
			2447 => "00000000000000000010011001000001",
			2448 => "0000001101000000000111111100011100",
			2449 => "0000000011000000001001001000000100",
			2450 => "00000000000000000010011010001101",
			2451 => "0000001010000000001010100000010100",
			2452 => "0000001100000000000011011100000100",
			2453 => "00000000000000000010011010001101",
			2454 => "0000000001000000000000111100001100",
			2455 => "0000000111000000000110000100000100",
			2456 => "00000000000000000010011010001101",
			2457 => "0000000111000000001000011000000100",
			2458 => "00000000010101110010011010001101",
			2459 => "00000000000000000010011010001101",
			2460 => "00000000000000000010011010001101",
			2461 => "00000000000000000010011010001101",
			2462 => "0000001010000000001010100000001000",
			2463 => "0000000010000000001100000000000100",
			2464 => "11111111110001000010011010001101",
			2465 => "00000000000000000010011010001101",
			2466 => "00000000000000000010011010001101",
			2467 => "0000000011000000001000011000001000",
			2468 => "0000000110000000001101011100000100",
			2469 => "00000000000000000010011011010001",
			2470 => "11111111110110010010011011010001",
			2471 => "0000001010000000000000001000011000",
			2472 => "0000000110000000000100110100010100",
			2473 => "0000000110000000000000111100000100",
			2474 => "00000000000000000010011011010001",
			2475 => "0000001011000000000100001000000100",
			2476 => "00000000000000000010011011010001",
			2477 => "0000001001000000000100111100001000",
			2478 => "0000001111000000001010011100000100",
			2479 => "00000000000000000010011011010001",
			2480 => "00000000011111100010011011010001",
			2481 => "00000000000000000010011011010001",
			2482 => "00000000000000000010011011010001",
			2483 => "00000000000000000010011011010001",
			2484 => "0000000101000000000101001000010000",
			2485 => "0000000110000000000001000100000100",
			2486 => "00000000000000000010011100100101",
			2487 => "0000000001000000001001011000001000",
			2488 => "0000001100000000001001110100000100",
			2489 => "11111111110111110010011100100101",
			2490 => "00000000000000000010011100100101",
			2491 => "00000000000000000010011100100101",
			2492 => "0000000111000000001000011000000100",
			2493 => "00000000000000000010011100100101",
			2494 => "0000000110000000000101010000010100",
			2495 => "0000001100000000001011000000000100",
			2496 => "00000000000000000010011100100101",
			2497 => "0000001011000000000010001000000100",
			2498 => "00000000000000000010011100100101",
			2499 => "0000000001000000001101111100001000",
			2500 => "0000000001000000001101011100000100",
			2501 => "00000000000000000010011100100101",
			2502 => "00000000010100010010011100100101",
			2503 => "00000000000000000010011100100101",
			2504 => "00000000000000000010011100100101",
			2505 => "0000001101000000000111111100011100",
			2506 => "0000000011000000001001001000000100",
			2507 => "00000000000000000010011101100001",
			2508 => "0000001001000000000100111100010100",
			2509 => "0000001100000000000011011100000100",
			2510 => "00000000000000000010011101100001",
			2511 => "0000001100000000001011000000001100",
			2512 => "0000000110000000000000111100000100",
			2513 => "00000000000000000010011101100001",
			2514 => "0000001111000000001010011100000100",
			2515 => "00000000000000000010011101100001",
			2516 => "00000000101000000010011101100001",
			2517 => "00000000000000000010011101100001",
			2518 => "00000000000000000010011101100001",
			2519 => "00000000000000000010011101100001",
			2520 => "0000000011000000001000001100101100",
			2521 => "0000001010000000000000001000100000",
			2522 => "0000001111000000001001001000001100",
			2523 => "0000000001000000000110101000001000",
			2524 => "0000001110000000000100001000000100",
			2525 => "00000000000000000010011111001101",
			2526 => "00000000000011000010011111001101",
			2527 => "11111111010010100010011111001101",
			2528 => "0000000010000000001110110100010000",
			2529 => "0000000001000000000000111100001100",
			2530 => "0000001110000000001011000000000100",
			2531 => "00000000000000000010011111001101",
			2532 => "0000001011000000000100001000000100",
			2533 => "00000000000000000010011111001101",
			2534 => "00000000011100100010011111001101",
			2535 => "00000000000000000010011111001101",
			2536 => "00000000000000000010011111001101",
			2537 => "0000001111000000000000010000001000",
			2538 => "0000001011000000000100010000000100",
			2539 => "11111111100100000010011111001101",
			2540 => "00000000000000000010011111001101",
			2541 => "00000000000000000010011111001101",
			2542 => "0000000001000000000101011100001000",
			2543 => "0000000111000000000111010000000100",
			2544 => "00000000100011010010011111001101",
			2545 => "00000000000000000010011111001101",
			2546 => "00000000000000000010011111001101",
			2547 => "0000000101000000000110100100001100",
			2548 => "0000001100000000000110000100001000",
			2549 => "0000000110000000001101011100000100",
			2550 => "00000000000000000010100001000001",
			2551 => "11111110110011010010100001000001",
			2552 => "00000000000000000010100001000001",
			2553 => "0000000011000000001111010100011100",
			2554 => "0000000001000000001001011000010000",
			2555 => "0000000011000000000000110100000100",
			2556 => "00000000000000000010100001000001",
			2557 => "0000001100000000001000000000001000",
			2558 => "0000001100000000000011011100000100",
			2559 => "00000000000000000010100001000001",
			2560 => "00000000001010000010100001000001",
			2561 => "00000000000000000010100001000001",
			2562 => "0000001100000000000100011000000100",
			2563 => "00000000000000000010100001000001",
			2564 => "0000001100000000001001110100000100",
			2565 => "11111111101101010010100001000001",
			2566 => "00000000000000000010100001000001",
			2567 => "0000001001000000000100111100010000",
			2568 => "0000000011000000000010010100001100",
			2569 => "0000001100000000001001110100001000",
			2570 => "0000000011000000001010000100000100",
			2571 => "00000000000000000010100001000001",
			2572 => "00000000010011100010100001000001",
			2573 => "00000000000000000010100001000001",
			2574 => "00000000000000000010100001000001",
			2575 => "00000000000000000010100001000001",
			2576 => "0000000000000000000001010100110100",
			2577 => "0000000010000000001110010000100000",
			2578 => "0000000001000000001101011100011000",
			2579 => "0000001100000000000011011100001000",
			2580 => "0000001011000000000101101100000100",
			2581 => "00000000000000000010100011001101",
			2582 => "11111111111011100010100011001101",
			2583 => "0000000110000000001001011000000100",
			2584 => "00000000000000000010100011001101",
			2585 => "0000000111000000000110000100000100",
			2586 => "00000000000000000010100011001101",
			2587 => "0000000111000000000000001100000100",
			2588 => "00000000100010100010100011001101",
			2589 => "00000000000000000010100011001101",
			2590 => "0000000011000000001001100000000100",
			2591 => "11111111100100100010100011001101",
			2592 => "00000000000000000010100011001101",
			2593 => "0000001111000000001100000000001100",
			2594 => "0000000110000000000100110100001000",
			2595 => "0000000001000000000000111100000100",
			2596 => "00000000100111010010100011001101",
			2597 => "00000000000000000010100011001101",
			2598 => "00000000000000000010100011001101",
			2599 => "0000000111000000001000011000000100",
			2600 => "00000000000000000010100011001101",
			2601 => "00000000000010100010100011001101",
			2602 => "0000001111000000001111010100001000",
			2603 => "0000000011000000001000001100000100",
			2604 => "11111111011100110010100011001101",
			2605 => "00000000000000000010100011001101",
			2606 => "0000000001000000000000111100001000",
			2607 => "0000000001000000001111001100000100",
			2608 => "00000000000000000010100011001101",
			2609 => "00000000010001000010100011001101",
			2610 => "11111111100111000010100011001101",
			2611 => "0000000110000000000100110100100100",
			2612 => "0000000100000000000010010100100000",
			2613 => "0000001100000000001001110100011100",
			2614 => "0000000010000000000110010000010100",
			2615 => "0000000111000000001100101000001100",
			2616 => "0000001000000000000010101100001000",
			2617 => "0000000010000000000100001000000100",
			2618 => "00000000000000000010100100101001",
			2619 => "00000000001010100010100100101001",
			2620 => "00000000000000000010100100101001",
			2621 => "0000001100000000001000000000000100",
			2622 => "11111111110111110010100100101001",
			2623 => "00000000000000000010100100101001",
			2624 => "0000000001000000000000111100000100",
			2625 => "00000000010011010010100100101001",
			2626 => "00000000000000000010100100101001",
			2627 => "00000000000000000010100100101001",
			2628 => "00000000000000000010100100101001",
			2629 => "0000001111000000000110001100001000",
			2630 => "0000001000000000001000100100000100",
			2631 => "00000000000000000010100100101001",
			2632 => "11111111101011000010100100101001",
			2633 => "00000000000000000010100100101001",
			2634 => "0000001011000000000010001000101100",
			2635 => "0000001010000000000111101100100000",
			2636 => "0000000000000000001010100100010000",
			2637 => "0000000001000000000110101000001100",
			2638 => "0000000010000000000100001000000100",
			2639 => "00000000000000000010100110101101",
			2640 => "0000001001000000000000111100000100",
			2641 => "00000000010001000010100110101101",
			2642 => "00000000000000000010100110101101",
			2643 => "00000000000000000010100110101101",
			2644 => "0000001010000000000100111100000100",
			2645 => "11111111110111110010100110101101",
			2646 => "0000001111000000000010001000000100",
			2647 => "00000000000000000010100110101101",
			2648 => "0000000110000000001101111100000100",
			2649 => "00000000000101110010100110101101",
			2650 => "00000000000000000010100110101101",
			2651 => "0000000011000000001100000000001000",
			2652 => "0000000000000000000110011100000100",
			2653 => "00000000000000000010100110101101",
			2654 => "11111111011110010010100110101101",
			2655 => "00000000000000000010100110101101",
			2656 => "0000001001000000000100111100010100",
			2657 => "0000001011000000001011110100010000",
			2658 => "0000001100000000001011000000000100",
			2659 => "00000000000000000010100110101101",
			2660 => "0000001110000000000110010000000100",
			2661 => "00000000000000000010100110101101",
			2662 => "0000001100000000001001110100000100",
			2663 => "00000000011110010010100110101101",
			2664 => "00000000000000000010100110101101",
			2665 => "00000000000000000010100110101101",
			2666 => "00000000000000000010100110101101",
			2667 => "0000001000000000001001000100101100",
			2668 => "0000001110000000001000011000001100",
			2669 => "0000001110000000001011000000000100",
			2670 => "11111110011100010010101001001001",
			2671 => "0000001101000000001111011100000100",
			2672 => "00000100011001110010101001001001",
			2673 => "11111110100100110010101001001001",
			2674 => "0000000001000000000000111100011000",
			2675 => "0000000111000000001111011100010100",
			2676 => "0000001011000000000101110100010000",
			2677 => "0000001110000000001100010000001000",
			2678 => "0000000110000000000100110100000100",
			2679 => "00000010001010000010101001001001",
			2680 => "00000000110001100010101001001001",
			2681 => "0000001100000000001000000000000100",
			2682 => "00000100111001110010101001001001",
			2683 => "00000010110101000010101001001001",
			2684 => "11111110101101110010101001001001",
			2685 => "11111101101100100010101001001001",
			2686 => "0000001101000000000011001000000100",
			2687 => "11111110011011010010101001001001",
			2688 => "00000000011100110010101001001001",
			2689 => "0000001000000000000001010000010000",
			2690 => "0000000100000000001101101100001100",
			2691 => "0000000001000000000000111100001000",
			2692 => "0000000100000000001000001100000100",
			2693 => "11111110111100110010101001001001",
			2694 => "00000001000110110010101001001001",
			2695 => "11111110011101010010101001001001",
			2696 => "00000011010100000010101001001001",
			2697 => "0000001101000000000011000000001100",
			2698 => "0000001000000000001100011100001000",
			2699 => "0000001000000000001010110000000100",
			2700 => "11111110011100010010101001001001",
			2701 => "00000000000000000010101001001001",
			2702 => "11111110011000010010101001001001",
			2703 => "0000001000000000001110111100000100",
			2704 => "00000100111000000010101001001001",
			2705 => "11111110011010010010101001001001",
			2706 => "0000001100000000000011011100001100",
			2707 => "0000001101000000001010001100001000",
			2708 => "0000001010000000001100011000000100",
			2709 => "00000000000000000010101011010101",
			2710 => "11111110111101110010101011010101",
			2711 => "00000000000000000010101011010101",
			2712 => "0000000011000000001111010100100100",
			2713 => "0000001100000000001011000000011000",
			2714 => "0000001101000000001110101000010000",
			2715 => "0000000111000000001101111000001100",
			2716 => "0000000111000000000110000100000100",
			2717 => "00000000000000000010101011010101",
			2718 => "0000001100000000000110000100000100",
			2719 => "00000000001111110010101011010101",
			2720 => "00000000000000000010101011010101",
			2721 => "11111111110100010010101011010101",
			2722 => "0000001001000000000100111100000100",
			2723 => "00000000101101100010101011010101",
			2724 => "00000000000000000010101011010101",
			2725 => "0000000001000000001001011000001000",
			2726 => "0000001000000000000111110100000100",
			2727 => "00000000000000000010101011010101",
			2728 => "11111111001000000010101011010101",
			2729 => "00000000000000000010101011010101",
			2730 => "0000000001000000000000111100001000",
			2731 => "0000000111000000001111011100000100",
			2732 => "00000000101100100010101011010101",
			2733 => "00000000000000000010101011010101",
			2734 => "0000001101000000000110010000000100",
			2735 => "11111111110100010010101011010101",
			2736 => "0000001100000000001011011100001000",
			2737 => "0000001110000000000000010100000100",
			2738 => "00000000000101000010101011010101",
			2739 => "00000000000000000010101011010101",
			2740 => "00000000000000000010101011010101",
			2741 => "0000001010000000001010100000110000",
			2742 => "0000001110000000000101110100011000",
			2743 => "0000000110000000001101011100001000",
			2744 => "0000001110000000000100001000000100",
			2745 => "11111110100101010010101110001001",
			2746 => "00000100110110100010101110001001",
			2747 => "0000001011000000000100001000000100",
			2748 => "11111110001111110010101110001001",
			2749 => "0000001001000000000001000100001000",
			2750 => "0000000101000000000001101000000100",
			2751 => "11111111001010010010101110001001",
			2752 => "00000011100101010010101110001001",
			2753 => "11111110011110010010101110001001",
			2754 => "0000001001000000000100111100010100",
			2755 => "0000000111000000001111011100010000",
			2756 => "0000000011000000001010000100001100",
			2757 => "0000000101000000001111010000001000",
			2758 => "0000001110000000001110101000000100",
			2759 => "00000001011110110010101110001001",
			2760 => "00000010100001000010101110001001",
			2761 => "00000000011000000010101110001001",
			2762 => "00000100000000110010101110001001",
			2763 => "00000000100101100010101110001001",
			2764 => "11111110100000010010101110001001",
			2765 => "0000001010000000000010101100011000",
			2766 => "0000000010000000001010000100001100",
			2767 => "0000000011000000001000001100000100",
			2768 => "11111110011000100010101110001001",
			2769 => "0000000111000000001000011000000100",
			2770 => "00000010011000000010101110001001",
			2771 => "11111110011111100010101110001001",
			2772 => "0000001001000000000101010000001000",
			2773 => "0000000100000000001000100000000100",
			2774 => "00000010011110100010101110001001",
			2775 => "00000100110111000010101110001001",
			2776 => "11111110101111100010101110001001",
			2777 => "0000001010000000000010101100001000",
			2778 => "0000001101000000000100101000000100",
			2779 => "11111110100000000010101110001001",
			2780 => "00000001001100110010101110001001",
			2781 => "0000001101000000000011000000000100",
			2782 => "11111110010111100010101110001001",
			2783 => "0000001011000000000111111100000100",
			2784 => "00000010010011110010101110001001",
			2785 => "11111110011001010010101110001001",
			2786 => "0000000101000000000110100100001100",
			2787 => "0000000100000000000001101000000100",
			2788 => "00000000000000000010110000001101",
			2789 => "0000001110000000001000011000000100",
			2790 => "11111111011001000010110000001101",
			2791 => "00000000000000000010110000001101",
			2792 => "0000001010000000000000001000010000",
			2793 => "0000001110000000001011000000000100",
			2794 => "00000000000000000010110000001101",
			2795 => "0000001011000000000100001000000100",
			2796 => "00000000000000000010110000001101",
			2797 => "0000001001000000000100111100000100",
			2798 => "00000000010110000010110000001101",
			2799 => "00000000000000000010110000001101",
			2800 => "0000000011000000001000001100010100",
			2801 => "0000000101000000000111100000000100",
			2802 => "00000000000000000010110000001101",
			2803 => "0000001010000000001010100100001100",
			2804 => "0000001101000000000101110000000100",
			2805 => "00000000000000000010110000001101",
			2806 => "0000001011000000000101110100000100",
			2807 => "11111111101100000010110000001101",
			2808 => "00000000000000000010110000001101",
			2809 => "00000000000000000010110000001101",
			2810 => "0000001110000000001000101000010000",
			2811 => "0000000101000000000111100000000100",
			2812 => "00000000000000000010110000001101",
			2813 => "0000001011000000000001001000001000",
			2814 => "0000001010000000000001010000000100",
			2815 => "00000000010000010010110000001101",
			2816 => "00000000000000000010110000001101",
			2817 => "00000000000000000010110000001101",
			2818 => "00000000000000000010110000001101",
			2819 => "0000000011000000001100010000101000",
			2820 => "0000001010000000000111101100011100",
			2821 => "0000001100000000000110000100010100",
			2822 => "0000001111000000001010011100001000",
			2823 => "0000001011000000000101101100000100",
			2824 => "00000000000000000010110010110001",
			2825 => "11111111111100100010110010110001",
			2826 => "0000001100000000001000111100000100",
			2827 => "00000000000000000010110010110001",
			2828 => "0000000111000000001100101000000100",
			2829 => "00000000100011010010110010110001",
			2830 => "00000000000000000010110010110001",
			2831 => "0000000010000000001100100100000100",
			2832 => "11111111110001110010110010110001",
			2833 => "00000000000000000010110010110001",
			2834 => "0000001000000000000111110100000100",
			2835 => "00000000000000000010110010110001",
			2836 => "0000000111000000000001101000000100",
			2837 => "11111111000011000010110010110001",
			2838 => "00000000000000000010110010110001",
			2839 => "0000001001000000001100011000000100",
			2840 => "00000000000000000010110010110001",
			2841 => "0000001001000000000100111100011100",
			2842 => "0000001100000000001000000000001100",
			2843 => "0000000110000000000100110100001000",
			2844 => "0000000100000000000010000100000100",
			2845 => "00000000000000000010110010110001",
			2846 => "00000000101101010010110010110001",
			2847 => "00000000000000000010110010110001",
			2848 => "0000001101000000001010001000001000",
			2849 => "0000001101000000000111111100000100",
			2850 => "00000000000000000010110010110001",
			2851 => "11111111110101000010110010110001",
			2852 => "0000001101000000001100000000000100",
			2853 => "00000000000001110010110010110001",
			2854 => "00000000000000000010110010110001",
			2855 => "0000000011000000001000100000000100",
			2856 => "11111111111110110010110010110001",
			2857 => "0000001101000000001010001000000100",
			2858 => "00000000000000000010110010110001",
			2859 => "00000000000010000010110010110001",
			2860 => "0000001010000000001010100000110000",
			2861 => "0000001110000000001000011000001100",
			2862 => "0000001110000000001011000000000100",
			2863 => "11111110011011000010110101010101",
			2864 => "0000001101000000001111011100000100",
			2865 => "00000101101110100010110101010101",
			2866 => "11111110100010100010110101010101",
			2867 => "0000001001000000000100111100100000",
			2868 => "0000001011000000000101110100011100",
			2869 => "0000001110000000001100010000010000",
			2870 => "0000001010000000000000001000001000",
			2871 => "0000001001000000001110010100000100",
			2872 => "00000100110000010010110101010101",
			2873 => "00000010010011000010110101010101",
			2874 => "0000001001000000001111000000000100",
			2875 => "00000010010011100010110101010101",
			2876 => "11111111110110010010110101010101",
			2877 => "0000001100000000001001110100001000",
			2878 => "0000001100000000001000000000000100",
			2879 => "00000101101101000010110101010101",
			2880 => "00000011100010100010110101010101",
			2881 => "11111111000010000010110101010101",
			2882 => "11111110011101100010110101010101",
			2883 => "11111110011011110010110101010101",
			2884 => "0000001010000000000010101100010000",
			2885 => "0000000010000000001010000100001000",
			2886 => "0000001011000000000101110100000100",
			2887 => "11111110011011110010110101010101",
			2888 => "00000000011100000010110101010101",
			2889 => "0000000001000000000101011100000100",
			2890 => "00000011011111110010110101010101",
			2891 => "11111110101111100010110101010101",
			2892 => "0000001101000000000011000000001100",
			2893 => "0000001010000000000011101000001000",
			2894 => "0000001010000000000011101000000100",
			2895 => "11111110011011110010110101010101",
			2896 => "11111111111001110010110101010101",
			2897 => "11111110011000000010110101010101",
			2898 => "0000000010000000000011111000000100",
			2899 => "00000110010100110010110101010101",
			2900 => "11111110011001100010110101010101",
			2901 => "0000001100000000000011011100001000",
			2902 => "0000000110000000001101011100000100",
			2903 => "00000000000000000010110111100001",
			2904 => "11111111000111000010110111100001",
			2905 => "0000001101000000000111111100100100",
			2906 => "0000000110000000000100110100011000",
			2907 => "0000001111000000001100100100010000",
			2908 => "0000001100000000000110000100001100",
			2909 => "0000000110000000001001011000000100",
			2910 => "00000000000000000010110111100001",
			2911 => "0000000111000000000110000100000100",
			2912 => "00000000000000000010110111100001",
			2913 => "00000000100001010010110111100001",
			2914 => "11111111101000000010110111100001",
			2915 => "0000001001000000000100111100000100",
			2916 => "00000000101111100010110111100001",
			2917 => "00000000000000000010110111100001",
			2918 => "0000000101000000001111010000001000",
			2919 => "0000001010000000000000001000000100",
			2920 => "00000000000000000010110111100001",
			2921 => "11111111110001100010110111100001",
			2922 => "00000000000000000010110111100001",
			2923 => "0000000011000000001000001100001000",
			2924 => "0000001101000000001010001000000100",
			2925 => "11111111010010100010110111100001",
			2926 => "00000000000000000010110111100001",
			2927 => "0000000110000000001000010000010000",
			2928 => "0000001100000000001011000000000100",
			2929 => "00000000000000000010110111100001",
			2930 => "0000000110000000001010011000000100",
			2931 => "00000000000000000010110111100001",
			2932 => "0000001001000000001010100000000100",
			2933 => "00000000101010110010110111100001",
			2934 => "00000000000000000010110111100001",
			2935 => "00000000000000000010110111100001",
			2936 => "0000000111000000000110000100010000",
			2937 => "0000001111000000001011000000000100",
			2938 => "00000000000000000010111001110101",
			2939 => "0000000101000000001010011100001000",
			2940 => "0000000110000000001001011000000100",
			2941 => "00000000000000000010111001110101",
			2942 => "11111111011010110010111001110101",
			2943 => "00000000000000000010111001110101",
			2944 => "0000000111000000000001101000010100",
			2945 => "0000000000000000001100000100010000",
			2946 => "0000000110000000000000111100000100",
			2947 => "00000000000000000010111001110101",
			2948 => "0000001001000000001111000000001000",
			2949 => "0000001111000000001010011100000100",
			2950 => "00000000000000000010111001110101",
			2951 => "00000000100110000010111001110101",
			2952 => "00000000000000000010111001110101",
			2953 => "00000000000000000010111001110101",
			2954 => "0000000111000000001000011000010100",
			2955 => "0000001100000000000100011000000100",
			2956 => "00000000000000000010111001110101",
			2957 => "0000000100000000001000110100001100",
			2958 => "0000000110000000001101111100000100",
			2959 => "00000000000000000010111001110101",
			2960 => "0000001101000000001001010000000100",
			2961 => "00000000000000000010111001110101",
			2962 => "11111111100110000010111001110101",
			2963 => "00000000000000000010111001110101",
			2964 => "0000001100000000001011000000000100",
			2965 => "00000000000000000010111001110101",
			2966 => "0000001101000000000100101000000100",
			2967 => "00000000000000000010111001110101",
			2968 => "0000000110000000001000010000001000",
			2969 => "0000000101000000000001000000000100",
			2970 => "00000000000000000010111001110101",
			2971 => "00000000011011100010111001110101",
			2972 => "00000000000000000010111001110101",
			2973 => "0000001010000000001010100100110100",
			2974 => "0000000111000000000110000100010000",
			2975 => "0000001011000000001100101000001100",
			2976 => "0000001011000000000000001100000100",
			2977 => "11111110101000100010111100100001",
			2978 => "0000000101000000001001110100000100",
			2979 => "00000000100010000010111100100001",
			2980 => "00000000000000000010111100100001",
			2981 => "11111100101101000010111100100001",
			2982 => "0000000001000000000110101000000100",
			2983 => "00001011100100110010111100100001",
			2984 => "0000001001000000000100111100011100",
			2985 => "0000001111000000001011011100001100",
			2986 => "0000000001000000000111100100001000",
			2987 => "0000000001000000000111100100000100",
			2988 => "11111111011110010010111100100001",
			2989 => "00000000111110110010111100100001",
			2990 => "11111110100100010010111100100001",
			2991 => "0000001100000000001001110100001000",
			2992 => "0000001111000000001111010100000100",
			2993 => "00000001100100010010111100100001",
			2994 => "00000011011110000010111100100001",
			2995 => "0000001000000000001000100100000100",
			2996 => "00000001010100000010111100100001",
			2997 => "11111110011101110010111100100001",
			2998 => "11111110100110100010111100100001",
			2999 => "0000001010000000000111110100010000",
			3000 => "0000000010000000001000100000001100",
			3001 => "0000001011000000000101100100000100",
			3002 => "11111110010001010010111100100001",
			3003 => "0000001011000000001011011100000100",
			3004 => "00000001001001100010111100100001",
			3005 => "11111110100010000010111100100001",
			3006 => "00000011000000010010111100100001",
			3007 => "0000000101000000001111100100001100",
			3008 => "0000000010000000000010110000000100",
			3009 => "11111110011001010010111100100001",
			3010 => "0000000010000000001000001000000100",
			3011 => "00000101001110000010111100100001",
			3012 => "11111110011100110010111100100001",
			3013 => "0000001100000000001011011100000100",
			3014 => "00000100001111000010111100100001",
			3015 => "11111110100010110010111100100001",
			3016 => "0000001000000000001001000100101100",
			3017 => "0000001110000000001011000000000100",
			3018 => "11111110011101010010111110111101",
			3019 => "0000000001000000000000111100100000",
			3020 => "0000000111000000001111011100011100",
			3021 => "0000001110000000001110101000010000",
			3022 => "0000001100000000001100110000001000",
			3023 => "0000001011000000000100001000000100",
			3024 => "00000000011101000010111110111101",
			3025 => "00000011111110100010111110111101",
			3026 => "0000000111000000001101111000000100",
			3027 => "00000000001000000010111110111101",
			3028 => "11111110001100110010111110111101",
			3029 => "0000001011000000000101110100001000",
			3030 => "0000001110000000001100010000000100",
			3031 => "00000010000001000010111110111101",
			3032 => "00000011011100110010111110111101",
			3033 => "11111110110000100010111110111101",
			3034 => "11111101101101000010111110111101",
			3035 => "0000001101000000000011001000000100",
			3036 => "11111110011100010010111110111101",
			3037 => "00000000011111010010111110111101",
			3038 => "0000001010000000000010101100001100",
			3039 => "0000001111000000001010000100000100",
			3040 => "11111110011110100010111110111101",
			3041 => "0000000001000000000101011100000100",
			3042 => "00000011000101100010111110111101",
			3043 => "11111110101101100010111110111101",
			3044 => "0000001101000000000011000000010000",
			3045 => "0000001010000000000011101000001100",
			3046 => "0000001010000000000011101000000100",
			3047 => "11111110011101110010111110111101",
			3048 => "0000001000000000001010110000000100",
			3049 => "11111110110000100010111110111101",
			3050 => "00000010001010110010111110111101",
			3051 => "11111110011000100010111110111101",
			3052 => "0000001110000000000011010100000100",
			3053 => "00000011110111110010111110111101",
			3054 => "11111110011011000010111110111101",
			3055 => "0000001000000000001000100100110100",
			3056 => "0000001111000000000010001000011100",
			3057 => "0000001110000000000110100100010100",
			3058 => "0000000110000000001101011100001000",
			3059 => "0000000101000000001110110000000100",
			3060 => "11111110101100000011000010010001",
			3061 => "00001000100100110011000010010001",
			3062 => "0000001110000000001011000000000100",
			3063 => "11111110011001000011000010010001",
			3064 => "0000001101000000001111011100000100",
			3065 => "00000011001011000011000010010001",
			3066 => "11111110100111110011000010010001",
			3067 => "0000000110000000000000111100000100",
			3068 => "00010100110000010011000010010001",
			3069 => "11111110011101110011000010010001",
			3070 => "0000001001000000000100111100010100",
			3071 => "0000001011000000001110110000000100",
			3072 => "00001011011000010011000010010001",
			3073 => "0000000010000000001100100100000100",
			3074 => "11111110100000110011000010010001",
			3075 => "0000000011000000001010000100001000",
			3076 => "0000000010000000000010000100000100",
			3077 => "00000101010010000011000010010001",
			3078 => "00000001011110010011000010010001",
			3079 => "00001000101010110011000010010001",
			3080 => "11111110011010110011000010010001",
			3081 => "0000000000000000001001101000011000",
			3082 => "0000000001000000000000111100001100",
			3083 => "0000000010000000000111011000001000",
			3084 => "0000001001000000001111000000000100",
			3085 => "00000100010111100011000010010001",
			3086 => "11111110101010110011000010010001",
			3087 => "00001110010101000011000010010001",
			3088 => "0000000011000000000000010000000100",
			3089 => "11111110011000000011000010010001",
			3090 => "0000001011000000000101110100000100",
			3091 => "00000111000011000011000010010001",
			3092 => "11111110100010110011000010010001",
			3093 => "0000001010000000000010101100001100",
			3094 => "0000001101000000001111010000000100",
			3095 => "11111110011000000011000010010001",
			3096 => "0000000000000000001001101000000100",
			3097 => "11111110100010010011000010010001",
			3098 => "00000110010010100011000010010001",
			3099 => "0000001101000000000011000000000100",
			3100 => "11111110010101110011000010010001",
			3101 => "0000001101000000000010010100001100",
			3102 => "0000000101000000001000100000001000",
			3103 => "0000000101000000001111100100000100",
			3104 => "11111111011001100011000010010001",
			3105 => "00000001100111100011000010010001",
			3106 => "11111110101100110011000010010001",
			3107 => "11111110010110110011000010010001",
			3108 => "0000001001000000000100111100111100",
			3109 => "0000001110000000001010001000011100",
			3110 => "0000000000000000001100011100011000",
			3111 => "0000000111000000000000001100010000",
			3112 => "0000001100000000000011011100000100",
			3113 => "00000000000000000011000100010101",
			3114 => "0000001101000000001000011000000100",
			3115 => "00000000000000000011000100010101",
			3116 => "0000001100000000000110000100000100",
			3117 => "00000000010011100011000100010101",
			3118 => "00000000000000000011000100010101",
			3119 => "0000001101000000000000110100000100",
			3120 => "11111111111110110011000100010101",
			3121 => "00000000000000000011000100010101",
			3122 => "11111111010000110011000100010101",
			3123 => "0000000111000000001111011100011100",
			3124 => "0000000111000000001000011000010100",
			3125 => "0000000111000000000001101000001100",
			3126 => "0000001101000000000111111100001000",
			3127 => "0000000000000000000010101000000100",
			3128 => "00000000011100010011000100010101",
			3129 => "00000000000000000011000100010101",
			3130 => "00000000000000000011000100010101",
			3131 => "0000000001000000001001011000000100",
			3132 => "00000000000000000011000100010101",
			3133 => "11111111101001000011000100010101",
			3134 => "0000000011000000001100000000000100",
			3135 => "00000000000000000011000100010101",
			3136 => "00000000101100000011000100010101",
			3137 => "00000000000000000011000100010101",
			3138 => "0000000001000000000000111100000100",
			3139 => "00000000000000000011000100010101",
			3140 => "11111111100001110011000100010101",
			3141 => "0000000000000000000001010100110000",
			3142 => "0000000001000000000000111100101100",
			3143 => "0000000111000000001000011000101000",
			3144 => "0000001010000000000100111100011000",
			3145 => "0000001001000000000101011100001100",
			3146 => "0000001110000000000100001000000100",
			3147 => "00000000000000000011000110101001",
			3148 => "0000000001000000000110101000000100",
			3149 => "00000000100101000011000110101001",
			3150 => "00000000000000000011000110101001",
			3151 => "0000000110000000001001011000000100",
			3152 => "00000000000000000011000110101001",
			3153 => "0000001010000000001001100100000100",
			3154 => "11111111100111010011000110101001",
			3155 => "00000000000000000011000110101001",
			3156 => "0000000001000000000111100100000100",
			3157 => "00000000000000000011000110101001",
			3158 => "0000001001000000000100111100001000",
			3159 => "0000001111000000000010001000000100",
			3160 => "00000000000000000011000110101001",
			3161 => "00000000110000110011000110101001",
			3162 => "00000000000000000011000110101001",
			3163 => "00000000000000000011000110101001",
			3164 => "00000000000000000011000110101001",
			3165 => "0000001011000000000101100100001000",
			3166 => "0000000000000000000001110000000100",
			3167 => "00000000000000000011000110101001",
			3168 => "11111110110101000011000110101001",
			3169 => "0000001011000000000110110100001000",
			3170 => "0000001001000000000100111100000100",
			3171 => "00000000001110100011000110101001",
			3172 => "00000000000000000011000110101001",
			3173 => "0000000101000000001110010000001000",
			3174 => "0000001100000000000100011000000100",
			3175 => "00000000000000000011000110101001",
			3176 => "11111111011111010011000110101001",
			3177 => "00000000000000000011000110101001",
			3178 => "0000000000000000001011010101001100",
			3179 => "0000000110000000000100110100101000",
			3180 => "0000001110000000001110101000010100",
			3181 => "0000000110000000000001000100010000",
			3182 => "0000001100000000000110000100001100",
			3183 => "0000001110000000000100001000000100",
			3184 => "11111111110110000011001001011101",
			3185 => "0000000001000000000110101000000100",
			3186 => "00000001100000000011001001011101",
			3187 => "00000000100101000011001001011101",
			3188 => "11111111101100000011001001011101",
			3189 => "11111110011001100011001001011101",
			3190 => "0000001010000000001010100000010000",
			3191 => "0000000001000000000000111100001100",
			3192 => "0000001100000000000100011000000100",
			3193 => "00000001100011010011001001011101",
			3194 => "0000001100000000000100011000000100",
			3195 => "11111111010011100011001001011101",
			3196 => "00000001001101000011001001011101",
			3197 => "11111111111010000011001001011101",
			3198 => "11111111111111000011001001011101",
			3199 => "0000000011000000001000001100011000",
			3200 => "0000000100000000000111011000010000",
			3201 => "0000000101000000000111100000001000",
			3202 => "0000001100000000001010111000000100",
			3203 => "00000000000000000011001001011101",
			3204 => "11111111000011010011001001011101",
			3205 => "0000000001000000000000111100000100",
			3206 => "00000001000111010011001001011101",
			3207 => "00000000000000000011001001011101",
			3208 => "0000000001000000001001011000000100",
			3209 => "00000000000000000011001001011101",
			3210 => "11111110101000000011001001011101",
			3211 => "0000000001000000000101011100001000",
			3212 => "0000001100000000001001110100000100",
			3213 => "00000001010110100011001001011101",
			3214 => "00000000000000000011001001011101",
			3215 => "00000000000000000011001001011101",
			3216 => "0000000010000000000010110000000100",
			3217 => "11111110011010100011001001011101",
			3218 => "0000000110000000000101010000001000",
			3219 => "0000000001000000001101011100000100",
			3220 => "00000000000000000011001001011101",
			3221 => "00000001100111110011001001011101",
			3222 => "11111110111010110011001001011101",
			3223 => "0000001101000000001000011000001000",
			3224 => "0000000110000000001101011100000100",
			3225 => "00000000000000000011001100000001",
			3226 => "11111110101101000011001100000001",
			3227 => "0000001010000000001010100000100000",
			3228 => "0000000110000000000100110100010100",
			3229 => "0000001100000000000011011100000100",
			3230 => "00000000000000000011001100000001",
			3231 => "0000000011000000000110100100000100",
			3232 => "00000000000000000011001100000001",
			3233 => "0000001100000000001001110100001000",
			3234 => "0000001001000000000100111100000100",
			3235 => "00000000111000100011001100000001",
			3236 => "00000000000000000011001100000001",
			3237 => "00000000000000000011001100000001",
			3238 => "0000000011000000001010000100001000",
			3239 => "0000000111000000000001101000000100",
			3240 => "00000000000000000011001100000001",
			3241 => "11111111010100010011001100000001",
			3242 => "00000000000000000011001100000001",
			3243 => "0000000011000000001000001100010000",
			3244 => "0000001001000000001111000000001100",
			3245 => "0000001001000000001010011000000100",
			3246 => "11111111011000010011001100000001",
			3247 => "0000000010000000001011101100000100",
			3248 => "00000000010010100011001100000001",
			3249 => "00000000000000000011001100000001",
			3250 => "11111111001000110011001100000001",
			3251 => "0000000110000000001010011000010000",
			3252 => "0000000111000000000111010000001100",
			3253 => "0000001001000000000101010000001000",
			3254 => "0000001000000000001000010100000100",
			3255 => "00000000000000000011001100000001",
			3256 => "00000000111001100011001100000001",
			3257 => "00000000000000000011001100000001",
			3258 => "00000000000000000011001100000001",
			3259 => "0000001101000000001111101000000100",
			3260 => "11111111100010000011001100000001",
			3261 => "0000001100000000000010001000000100",
			3262 => "00000000001010000011001100000001",
			3263 => "00000000000000000011001100000001",
			3264 => "0000000000000000001101010001001100",
			3265 => "0000001010000000001010100000101000",
			3266 => "0000000110000000000100110100011000",
			3267 => "0000000110000000001001011000001000",
			3268 => "0000000001000000000110101000000100",
			3269 => "00000000000000000011001110011101",
			3270 => "11111111111011000011001110011101",
			3271 => "0000001100000000000011011100000100",
			3272 => "00000000000000000011001110011101",
			3273 => "0000000111000000000110000100000100",
			3274 => "00000000000000000011001110011101",
			3275 => "0000000001000000000000111100000100",
			3276 => "00000000111010000011001110011101",
			3277 => "00000000000000000011001110011101",
			3278 => "0000000011000000001010000100001100",
			3279 => "0000000001000000001001011000000100",
			3280 => "00000000000000000011001110011101",
			3281 => "0000001000000000001000100100000100",
			3282 => "00000000000000000011001110011101",
			3283 => "11111111010000010011001110011101",
			3284 => "00000000000000000011001110011101",
			3285 => "0000000011000000001000001100010000",
			3286 => "0000000010000000000110101100001100",
			3287 => "0000001111000000001100000000001000",
			3288 => "0000001111000000001100010000000100",
			3289 => "11111111110001010011001110011101",
			3290 => "00000000000000000011001110011101",
			3291 => "11111111010000100011001110011101",
			3292 => "00000000000000000011001110011101",
			3293 => "0000000001000000000101011100001100",
			3294 => "0000000111000000000111010000001000",
			3295 => "0000001000000000001000010100000100",
			3296 => "00000000000000000011001110011101",
			3297 => "00000000110110010011001110011101",
			3298 => "00000000000000000011001110011101",
			3299 => "0000000111000000000111110000000100",
			3300 => "11111111101100100011001110011101",
			3301 => "00000000000111100011001110011101",
			3302 => "11111110101111110011001110011101",
			3303 => "0000000000000000001011010101001100",
			3304 => "0000001001000000001111000000011000",
			3305 => "0000000111000000001101100000000100",
			3306 => "00000000000000000011010001001001",
			3307 => "0000000101000000001111010000010000",
			3308 => "0000000111000000001111011100001100",
			3309 => "0000001110000000001110101000001000",
			3310 => "0000001111000000001001110100000100",
			3311 => "00000001000011110011010001001001",
			3312 => "11111111110101000011010001001001",
			3313 => "00000001000101000011010001001001",
			3314 => "00000000000000000011010001001001",
			3315 => "00000000000000000011010001001001",
			3316 => "0000000101000000000101001000010100",
			3317 => "0000000000000000000101000100001000",
			3318 => "0000001101000000000101110000000100",
			3319 => "11111111110111000011010001001001",
			3320 => "00000000010000100011010001001001",
			3321 => "0000000100000000000110111100001000",
			3322 => "0000000111000000000110100100000100",
			3323 => "00000000000000000011010001001001",
			3324 => "11111110110010110011010001001001",
			3325 => "00000000000000000011010001001001",
			3326 => "0000000111000000001000011000010100",
			3327 => "0000000100000000001010000100001000",
			3328 => "0000001101000000000111111100000100",
			3329 => "00000000000000000011010001001001",
			3330 => "11111111001101110011010001001001",
			3331 => "0000000111000000001000011000001000",
			3332 => "0000000111000000001000011000000100",
			3333 => "00000000000000000011010001001001",
			3334 => "00000000100001010011010001001001",
			3335 => "00000000000000000011010001001001",
			3336 => "0000000111000000000111010000001000",
			3337 => "0000000001000000000101011100000100",
			3338 => "00000000110111010011010001001001",
			3339 => "00000000000000000011010001001001",
			3340 => "11111111110111000011010001001001",
			3341 => "0000001111000000000110001100000100",
			3342 => "11111110100111010011010001001001",
			3343 => "0000000110000000001000010000000100",
			3344 => "00000000101001100011010001001001",
			3345 => "00000000000000000011010001001001",
			3346 => "0000000000000000001001101001000100",
			3347 => "0000001110000000001110101000011000",
			3348 => "0000000010000000000000110100010100",
			3349 => "0000000001000000001101101000010000",
			3350 => "0000001110000000000001101000001100",
			3351 => "0000000001000000000110101000001000",
			3352 => "0000001101000000000110100100000100",
			3353 => "11111111010001010011010100001101",
			3354 => "00000001101010010011010100001101",
			3355 => "11111110110000110011010100001101",
			3356 => "00000001100011000011010100001101",
			3357 => "11111110111000110011010100001101",
			3358 => "11111110100100010011010100001101",
			3359 => "0000001001000000001111000000001000",
			3360 => "0000001011000000000010001000000100",
			3361 => "00000001100101100011010100001101",
			3362 => "11111111100011000011010100001101",
			3363 => "0000000011000000001100000000001000",
			3364 => "0000001010000000000000001000000100",
			3365 => "11111111111101010011010100001101",
			3366 => "11111101110001010011010100001101",
			3367 => "0000001100000000001000000000010000",
			3368 => "0000000000000000000001110000001000",
			3369 => "0000000011000000000110111100000100",
			3370 => "00000000011010110011010100001101",
			3371 => "00000001110100000011010100001101",
			3372 => "0000001110000000001111010100000100",
			3373 => "11111111000011000011010100001101",
			3374 => "00000000000000000011010100001101",
			3375 => "0000001001000000001111000000000100",
			3376 => "11111110001010100011010100001101",
			3377 => "0000001101000000001010001000000100",
			3378 => "11111111111110110011010100001101",
			3379 => "00000001011001100011010100001101",
			3380 => "0000000010000000000010110000010100",
			3381 => "0000001000000000000110011100010000",
			3382 => "0000001101000000001111010000000100",
			3383 => "11111110101101010011010100001101",
			3384 => "0000001011000000001011011100001000",
			3385 => "0000001110000000000110111100000100",
			3386 => "00000001011011000011010100001101",
			3387 => "00000000000000000011010100001101",
			3388 => "11111111000100000011010100001101",
			3389 => "11111110011010000011010100001101",
			3390 => "0000001010000000000001010000001000",
			3391 => "0000000001000000001101011000000100",
			3392 => "00000011000011010011010100001101",
			3393 => "00000000000000000011010100001101",
			3394 => "11111110100110110011010100001101",
			3395 => "0000001000000000001001000101001000",
			3396 => "0000001001000000000100111101000000",
			3397 => "0000001110000000001110101000101000",
			3398 => "0000001100000000001100110000011000",
			3399 => "0000001011000000000100001000010000",
			3400 => "0000000110000000001101011100001000",
			3401 => "0000000011000000000100001000000100",
			3402 => "11111111001101100011010111010001",
			3403 => "00000100010101110011010111010001",
			3404 => "0000001101000000001111011100000100",
			3405 => "11111110011111000011010111010001",
			3406 => "00000000000000000011010111010001",
			3407 => "0000000110000000000101011100000100",
			3408 => "00000101000001010011010111010001",
			3409 => "00000001101111010011010111010001",
			3410 => "0000000110000000000101011100001100",
			3411 => "0000000111000000001110001100001000",
			3412 => "0000001011000000001010111100000100",
			3413 => "11111111000100100011010111010001",
			3414 => "00000001001110010011010111010001",
			3415 => "11111110011101100011010111010001",
			3416 => "11111101111010100011010111010001",
			3417 => "0000000011000000001000001100010100",
			3418 => "0000000000000000000001010100001100",
			3419 => "0000001001000000000100111100001000",
			3420 => "0000001110000000000010000100000100",
			3421 => "00000001111001010011010111010001",
			3422 => "00000010111110010011010111010001",
			3423 => "11111110111100010011010111010001",
			3424 => "0000001001000000001111000000000100",
			3425 => "00000001000111100011010111010001",
			3426 => "11111110010001100011010111010001",
			3427 => "00000100001010010011010111010001",
			3428 => "0000000000000000001100000100000100",
			3429 => "11111110011101100011010111010001",
			3430 => "00000001011010100011010111010001",
			3431 => "0000001010000000000011101000010000",
			3432 => "0000000010000000000110101100001100",
			3433 => "0000001011000000000101100100000100",
			3434 => "11111110011011100011010111010001",
			3435 => "0000001110000000001100000000000100",
			3436 => "00000001100010100011010111010001",
			3437 => "11111110100001000011010111010001",
			3438 => "00000011111110110011010111010001",
			3439 => "0000000101000000001111100100000100",
			3440 => "11111110011000010011010111010001",
			3441 => "0000000101000000001000100000000100",
			3442 => "00000000010101110011010111010001",
			3443 => "11111110011101000011010111010001",
			3444 => "0000000000000000001011010101000100",
			3445 => "0000001000000000000111110100100000",
			3446 => "0000000010000000001101000100011100",
			3447 => "0000000001000000000111100100010000",
			3448 => "0000001110000000000100001000000100",
			3449 => "11111111010100100011011010001101",
			3450 => "0000000111000000001110001100001000",
			3451 => "0000001001000000000000111100000100",
			3452 => "00000010000100100011011010001101",
			3453 => "00000000110010100011011010001101",
			3454 => "00000000000000000011011010001101",
			3455 => "0000001100000000001100110000001000",
			3456 => "0000000111000000001110001100000100",
			3457 => "11111111101000110011011010001101",
			3458 => "00000000001101010011011010001101",
			3459 => "11111110101010110011011010001101",
			3460 => "00000001100101000011011010001101",
			3461 => "0000001110000000001110010000000100",
			3462 => "11111101010100010011011010001101",
			3463 => "0000001010000000000000001000000100",
			3464 => "00000001100100110011011010001101",
			3465 => "0000000010000000001100000000010000",
			3466 => "0000001101000000000111111100001000",
			3467 => "0000000100000000001100010000000100",
			3468 => "11111110100100100011011010001101",
			3469 => "00000000110000100011011010001101",
			3470 => "0000001100000000001001110100000100",
			3471 => "11111101110111010011011010001101",
			3472 => "00000000110110010011011010001101",
			3473 => "0000001010000000001010100000000100",
			3474 => "00000010010011100011011010001101",
			3475 => "0000000001000000000101011100000100",
			3476 => "00000000101011110011011010001101",
			3477 => "11111110110110010011011010001101",
			3478 => "0000001101000000000011000000010100",
			3479 => "0000001010000000000111110100010000",
			3480 => "0000001100000000000100011000000100",
			3481 => "11111110010111010011011010001101",
			3482 => "0000000000000000001111001000001000",
			3483 => "0000001100000000001000000000000100",
			3484 => "00000000000000000011011010001101",
			3485 => "11111111011001000011011010001101",
			3486 => "00000001000111000011011010001101",
			3487 => "11111110011001110011011010001101",
			3488 => "0000001110000000000011110100000100",
			3489 => "00000001111110100011011010001101",
			3490 => "11111111000011000011011010001101",
			3491 => "0000000111000000001101100000000100",
			3492 => "11111110011100100011011100011001",
			3493 => "0000000000000000000110011100001100",
			3494 => "0000000001000000001001011000001000",
			3495 => "0000001110000000000100001000000100",
			3496 => "00000000000000000011011100011001",
			3497 => "00000001000100000011011100011001",
			3498 => "00000000000000000011011100011001",
			3499 => "0000001011000000000101100100001100",
			3500 => "0000001000000000000111110100000100",
			3501 => "00000000000000000011011100011001",
			3502 => "0000001111000000001111100100000100",
			3503 => "11111110100001110011011100011001",
			3504 => "00000000000000000011011100011001",
			3505 => "0000000011000000001111010100010000",
			3506 => "0000001000000000001000100100001000",
			3507 => "0000001101000000001001010000000100",
			3508 => "11111111110010100011011100011001",
			3509 => "00000001001111000011011100011001",
			3510 => "0000000001000000001001011000000100",
			3511 => "00000000000000010011011100011001",
			3512 => "11111110010111110011011100011001",
			3513 => "0000000111000000001111011100001100",
			3514 => "0000000001000000000000111100001000",
			3515 => "0000000011000000001000001100000100",
			3516 => "00000000110000100011011100011001",
			3517 => "00000010010001000011011100011001",
			3518 => "11111111000100000011011100011001",
			3519 => "0000001101000000000011000000001000",
			3520 => "0000001100000000001011000000000100",
			3521 => "00000000000000000011011100011001",
			3522 => "11111110110000110011011100011001",
			3523 => "0000000111000000000000110100000100",
			3524 => "00000001000100010011011100011001",
			3525 => "00000000000000000011011100011001",
			3526 => "0000000000000000001011010101010100",
			3527 => "0000001000000000000111110100100000",
			3528 => "0000001111000000001100100100011100",
			3529 => "0000000001000000000111100100010000",
			3530 => "0000000011000000000110100100001000",
			3531 => "0000000110000000001111001100000100",
			3532 => "00000001010101100011011111110101",
			3533 => "11111110111011010011011111110101",
			3534 => "0000000111000000001110001100000100",
			3535 => "00000001111010100011011111110101",
			3536 => "00000000000000000011011111110101",
			3537 => "0000001100000000001100110000001000",
			3538 => "0000000111000000001110001100000100",
			3539 => "11111111100001100011011111110101",
			3540 => "00000000010000110011011111110101",
			3541 => "11111110100111100011011111110101",
			3542 => "00000001100101110011011111110101",
			3543 => "0000000011000000001001100000001100",
			3544 => "0000000111000000000001101000001000",
			3545 => "0000001111000000000010000000000100",
			3546 => "11111110001000100011011111110101",
			3547 => "00000000000000000011011111110101",
			3548 => "11111011001001100011011111110101",
			3549 => "0000001010000000000000001000001100",
			3550 => "0000000011000000001100010000001000",
			3551 => "0000000110000000001101111100000100",
			3552 => "00000001001111100011011111110101",
			3553 => "11111101111111000011011111110101",
			3554 => "00000001101010000011011111110101",
			3555 => "0000000011000000000111010100010000",
			3556 => "0000001011000000000100010000001000",
			3557 => "0000001111000000001100000000000100",
			3558 => "00000000101110100011011111110101",
			3559 => "11111110110100110011011111110101",
			3560 => "0000001100000000001000000000000100",
			3561 => "11111111010110010011011111110101",
			3562 => "11111011000100000011011111110101",
			3563 => "0000001100000000001001110100001000",
			3564 => "0000001001000000000100111100000100",
			3565 => "00000010000110100011011111110101",
			3566 => "00000000000000000011011111110101",
			3567 => "11111110101100110011011111110101",
			3568 => "0000001101000000000011000000010100",
			3569 => "0000001010000000000111110100010000",
			3570 => "0000001100000000000100011000000100",
			3571 => "11111110010100100011011111110101",
			3572 => "0000001011000000001011011100001000",
			3573 => "0000001011000000000101100100000100",
			3574 => "00000000000000000011011111110101",
			3575 => "00000001101001110011011111110101",
			3576 => "11111111001111010011011111110101",
			3577 => "11111110011001110011011111110101",
			3578 => "0000000111000000000000110100000100",
			3579 => "00000010000111100011011111110101",
			3580 => "11111110111101110011011111110101",
			3581 => "0000001000000000001001000101010000",
			3582 => "0000001000000000000111110100100000",
			3583 => "0000000010000000001101000100011100",
			3584 => "0000000001000000000111100100010000",
			3585 => "0000001110000000000100001000000100",
			3586 => "11111111001101000011100011001001",
			3587 => "0000000111000000001110001100001000",
			3588 => "0000000111000000001101100000000100",
			3589 => "00000000000000000011100011001001",
			3590 => "00000001111011000011100011001001",
			3591 => "00000000000000000011100011001001",
			3592 => "0000001100000000001100110000001000",
			3593 => "0000000111000000001110001100000100",
			3594 => "11111111011110010011100011001001",
			3595 => "00000000010110110011100011001001",
			3596 => "11111110100011110011100011001001",
			3597 => "00000001100110100011100011001001",
			3598 => "0000000010000000001110010000001000",
			3599 => "0000001010000000000111101100000100",
			3600 => "11111010011001000011100011001001",
			3601 => "11111111000100000011100011001001",
			3602 => "0000001010000000000000001000001100",
			3603 => "0000000011000000001100010000001000",
			3604 => "0000001001000000001111000000000100",
			3605 => "00000001011000000011100011001001",
			3606 => "11111100110010110011100011001001",
			3607 => "00000001101011000011100011001001",
			3608 => "0000000010000000001100000000010000",
			3609 => "0000001101000000000111111100001000",
			3610 => "0000000011000000000110111100000100",
			3611 => "11111111100011000011100011001001",
			3612 => "00000001011001110011100011001001",
			3613 => "0000001100000000001001110100000100",
			3614 => "11111101010110000011100011001001",
			3615 => "00000000110001100011100011001001",
			3616 => "0000001011000000000100010000001000",
			3617 => "0000001010000000001010100000000100",
			3618 => "00000010100111010011100011001001",
			3619 => "00000000110111010011100011001001",
			3620 => "11111110110010100011100011001001",
			3621 => "0000001101000000000011000000010100",
			3622 => "0000001010000000000111110100010000",
			3623 => "0000000010000000001000100000001100",
			3624 => "0000001100000000001000000000000100",
			3625 => "11111110010011110011100011001001",
			3626 => "0000001100000000001001001000000100",
			3627 => "00000000000000000011100011001001",
			3628 => "11111110111010000011100011001001",
			3629 => "00000001101101010011100011001001",
			3630 => "11111110011001110011100011001001",
			3631 => "0000001001000000001010011000000100",
			3632 => "11111110111000110011100011001001",
			3633 => "00000010010010100011100011001001",
			3634 => "0000001010000000000111110100111100",
			3635 => "0000001001000000001000010000111000",
			3636 => "0000001111000000001111010100110000",
			3637 => "0000000000000000000001010100100000",
			3638 => "0000000101000000000111100000010000",
			3639 => "0000001100000000001011000000001000",
			3640 => "0000000011000000000000110100000100",
			3641 => "00000000000010000011100101010101",
			3642 => "00000000111100000011100101010101",
			3643 => "0000001000000000000111110100000100",
			3644 => "00000000000000000011100101010101",
			3645 => "11111110110100110011100101010101",
			3646 => "0000001000000000001000100100001000",
			3647 => "0000000011000000001100000000000100",
			3648 => "00000000000000000011100101010101",
			3649 => "00000001010101110011100101010101",
			3650 => "0000001100000000001011000000000100",
			3651 => "00000000000000000011100101010101",
			3652 => "00000000010001000011100101010101",
			3653 => "0000000011000000001000001100001100",
			3654 => "0000000101000000000111100000001000",
			3655 => "0000000101000000000010110100000100",
			3656 => "11111111101000000011100101010101",
			3657 => "00000000001001100011100101010101",
			3658 => "11111110111110100011100101010101",
			3659 => "00000000011110010011100101010101",
			3660 => "0000001011000000000101110100000100",
			3661 => "00000001100010000011100101010101",
			3662 => "00000000000000000011100101010101",
			3663 => "11111111000011100011100101010101",
			3664 => "0000001101000000000011000000000100",
			3665 => "11111110011111110011100101010101",
			3666 => "0000000111000000000000110100000100",
			3667 => "00000000010011110011100101010101",
			3668 => "00000000000000000011100101010101",
			3669 => "0000000111000000001101100000000100",
			3670 => "11111110110110110011100111101001",
			3671 => "0000001010000000000111101100001000",
			3672 => "0000001110000000000100001000000100",
			3673 => "00000000000000000011100111101001",
			3674 => "00000000101101100011100111101001",
			3675 => "0000000011000000001010000100100000",
			3676 => "0000000011000000001100010000001100",
			3677 => "0000001000000000000111110100000100",
			3678 => "00000000000000000011100111101001",
			3679 => "0000001010000000000111101100000100",
			3680 => "00000000000000000011100111101001",
			3681 => "11111110111110010011100111101001",
			3682 => "0000001101000000000111111100001100",
			3683 => "0000000001000000000000111100001000",
			3684 => "0000000111000000001111011100000100",
			3685 => "00000000101111000011100111101001",
			3686 => "00000000000000000011100111101001",
			3687 => "00000000000000000011100111101001",
			3688 => "0000000111000000001111011100000100",
			3689 => "11111111000110100011100111101001",
			3690 => "00000000000000000011100111101001",
			3691 => "0000001011000000000010001000001000",
			3692 => "0000001101000000000111111100000100",
			3693 => "00000000000000000011100111101001",
			3694 => "11111111101101110011100111101001",
			3695 => "0000000111000000000111010000001100",
			3696 => "0000000001000000000101011100001000",
			3697 => "0000000111000000001000011000000100",
			3698 => "00000000000000000011100111101001",
			3699 => "00000001000010010011100111101001",
			3700 => "00000000000000000011100111101001",
			3701 => "0000001101000000001111101000000100",
			3702 => "11111111110100000011100111101001",
			3703 => "0000000111000000001110101100000100",
			3704 => "00000000000000010011100111101001",
			3705 => "00000000000000000011100111101001",
			3706 => "0000000111000000001101100000000100",
			3707 => "11111110101010010011101010010101",
			3708 => "0000001010000000000111101100010100",
			3709 => "0000000001000000000111100100001000",
			3710 => "0000001111000000000001111100000100",
			3711 => "00000000000000000011101010010101",
			3712 => "00000000110101000011101010010101",
			3713 => "0000000010000000001101000100001000",
			3714 => "0000001100000000001100110000000100",
			3715 => "00000000000000000011101010010101",
			3716 => "11111111011011100011101010010101",
			3717 => "00000000110100110011101010010101",
			3718 => "0000000101000000000101001000100000",
			3719 => "0000001100000000001000000000010100",
			3720 => "0000000111000000001000000000000100",
			3721 => "11111110111101010011101010010101",
			3722 => "0000001100000000000100011000001000",
			3723 => "0000000000000000001100000100000100",
			3724 => "00000000011111000011101010010101",
			3725 => "00000000000000000011101010010101",
			3726 => "0000001000000000001000100100000100",
			3727 => "00000000000000000011101010010101",
			3728 => "11111111101100000011101010010101",
			3729 => "0000000111000000000001101000000100",
			3730 => "00000000000000000011101010010101",
			3731 => "0000001100000000001001110100000100",
			3732 => "11111110110000010011101010010101",
			3733 => "00000000000000000011101010010101",
			3734 => "0000000001000000000000111100010100",
			3735 => "0000000111000000001111011100010000",
			3736 => "0000000011000000001010000100001000",
			3737 => "0000001111000000001100000000000100",
			3738 => "00000000001000000011101010010101",
			3739 => "11111111110100110011101010010101",
			3740 => "0000001000000000001000100100000100",
			3741 => "00000000000000000011101010010101",
			3742 => "00000001001111100011101010010101",
			3743 => "00000000000000000011101010010101",
			3744 => "0000000011000000001111100000001000",
			3745 => "0000001011000000000100010000000100",
			3746 => "00000000000000000011101010010101",
			3747 => "11111111011100110011101010010101",
			3748 => "00000000000101000011101010010101",
			3749 => "0000000111000000001101100000000100",
			3750 => "11111110011110100011101101000001",
			3751 => "0000000000000000000001010100111000",
			3752 => "0000000011000000000110111100110000",
			3753 => "0000001100000000000100011000011000",
			3754 => "0000001111000000001100100100001100",
			3755 => "0000001100000000000110000100001000",
			3756 => "0000001011000000000100001000000100",
			3757 => "00000000000000000011101101000001",
			3758 => "00000000111110010011101101000001",
			3759 => "11111111000110100011101101000001",
			3760 => "0000000001000000000000111100001000",
			3761 => "0000001100000000000100011000000100",
			3762 => "00000001011000010011101101000001",
			3763 => "00000000000000000011101101000001",
			3764 => "00000000000000000011101101000001",
			3765 => "0000000111000000000001101000001000",
			3766 => "0000001001000000001111000000000100",
			3767 => "00000000110010110011101101000001",
			3768 => "00000000000000000011101101000001",
			3769 => "0000000001000000001001011000001000",
			3770 => "0000001001000000001001100100000100",
			3771 => "00000000000000000011101101000001",
			3772 => "11111110100001000011101101000001",
			3773 => "0000000001000000000000111100000100",
			3774 => "00000000110001000011101101000001",
			3775 => "11111111010110010011101101000001",
			3776 => "0000000101000000001110000100000100",
			3777 => "00000000000000000011101101000001",
			3778 => "00000001011000100011101101000001",
			3779 => "0000000011000000001000001100001000",
			3780 => "0000001111000000000000010000000100",
			3781 => "11111111000010010011101101000001",
			3782 => "00000000000000000011101101000001",
			3783 => "0000000001000000000101011100001100",
			3784 => "0000000111000000001111011100000100",
			3785 => "00000001101101010011101101000001",
			3786 => "0000001100000000001001110100000100",
			3787 => "00000000000110010011101101000001",
			3788 => "11111111101001010011101101000001",
			3789 => "0000000101000000000111010100000100",
			3790 => "11111110110101010011101101000001",
			3791 => "00000000100111000011101101000001",
			3792 => "0000000111000000001101100000000100",
			3793 => "11111110101101100011101111110101",
			3794 => "0000001010000000000111101100010000",
			3795 => "0000000001000000001101011100001100",
			3796 => "0000001111000000000001111100000100",
			3797 => "00000000000000000011101111110101",
			3798 => "0000000100000000001001100000000100",
			3799 => "00000000100010100011101111110101",
			3800 => "00000000000000000011101111110101",
			3801 => "00000000000000000011101111110101",
			3802 => "0000000011000000000110111100011100",
			3803 => "0000000111000000000001101000001100",
			3804 => "0000000011000000000110010000000100",
			3805 => "11111111010111110011101111110101",
			3806 => "0000000110000000000100110100000100",
			3807 => "00000000011010100011101111110101",
			3808 => "00000000000000000011101111110101",
			3809 => "0000000110000000001101111100000100",
			3810 => "00000000000000000011101111110101",
			3811 => "0000001100000000000100011000000100",
			3812 => "00000000000000000011101111110101",
			3813 => "0000001100000000001001110100000100",
			3814 => "11111110111010100011101111110101",
			3815 => "00000000000000000011101111110101",
			3816 => "0000000111000000001000011000011000",
			3817 => "0000001111000000000111011000001100",
			3818 => "0000000111000000000001101000001000",
			3819 => "0000001001000000000100111100000100",
			3820 => "00000000100011010011101111110101",
			3821 => "00000000000000000011101111110101",
			3822 => "00000000000000000011101111110101",
			3823 => "0000001101000000000111111100000100",
			3824 => "00000000000000000011101111110101",
			3825 => "0000001101000000001110010000000100",
			3826 => "11111110110111000011101111110101",
			3827 => "00000000000000000011101111110101",
			3828 => "0000000001000000000000111100001100",
			3829 => "0000000111000000001111011100001000",
			3830 => "0000001101000000000100101000000100",
			3831 => "00000000000000000011101111110101",
			3832 => "00000000110011010011101111110101",
			3833 => "00000000000000000011101111110101",
			3834 => "0000000011000000001111100000000100",
			3835 => "11111111100101100011101111110101",
			3836 => "00000000000011010011101111110101",
			3837 => "0000000111000000001101100000000100",
			3838 => "11111110100000100011110010011011",
			3839 => "0000001010000000000001010001001100",
			3840 => "0000000111000000001000011000110000",
			3841 => "0000001010000000000111101100010100",
			3842 => "0000000010000000001101000100010000",
			3843 => "0000000001000000000110101000001000",
			3844 => "0000001100000000001000111000000100",
			3845 => "00000001001010010011110010011011",
			3846 => "00000000000000000011110010011011",
			3847 => "0000001100000000001100110000000100",
			3848 => "00000000000000000011110010011011",
			3849 => "11111111001100000011110010011011",
			3850 => "00000001001011010011110010011011",
			3851 => "0000000011000000001100010000001100",
			3852 => "0000000000000000000110011100000100",
			3853 => "00000000000000000011110010011011",
			3854 => "0000000111000000000001101000000100",
			3855 => "11111110110100110011110010011011",
			3856 => "00000000000000000011110010011011",
			3857 => "0000001010000000000000001000001000",
			3858 => "0000001001000000000100111100000100",
			3859 => "00000001000110000011110010011011",
			3860 => "00000000000000000011110010011011",
			3861 => "0000000110000000001101111100000100",
			3862 => "11111111001100100011110010011011",
			3863 => "00000000000000000011110010011011",
			3864 => "0000000111000000001111011100001100",
			3865 => "0000000001000000000000111100001000",
			3866 => "0000000010000000000110010000000100",
			3867 => "00000000000000000011110010011011",
			3868 => "00000001010001000011110010011011",
			3869 => "00000000000000000011110010011011",
			3870 => "0000001110000000001011111000000100",
			3871 => "11111111010101010011110010011011",
			3872 => "0000000001000000001101111100001000",
			3873 => "0000001000000000001001101000000100",
			3874 => "00000000110010000011110010011011",
			3875 => "00000000000000000011110010011011",
			3876 => "00000000000000000011110010011011",
			3877 => "11111111000001010011110010011011",
			3878 => "00000000000000000011110010011101",
			3879 => "00000000000000000011110010100001",
			3880 => "00000000000000000011110010100101",
			3881 => "00000000000000000011110010101001",
			3882 => "00000000000000000011110010101101",
			3883 => "00000000000000000011110010110001",
			3884 => "00000000000000000011110010110101",
			3885 => "00000000000000000011110010111001",
			3886 => "0000001000000000001001111100001000",
			3887 => "0000001111000000000001111100000100",
			3888 => "00000000000000000011110011010101",
			3889 => "00000000000101000011110011010101",
			3890 => "0000001111000000001100010100000100",
			3891 => "11111111111010000011110011010101",
			3892 => "00000000000000000011110011010101",
			3893 => "0000000011000000000111010100001000",
			3894 => "0000000011000000001101010100000100",
			3895 => "00000000000000000011110011110001",
			3896 => "11111111111010110011110011110001",
			3897 => "0000000011000000000010100100000100",
			3898 => "00000000000001000011110011110001",
			3899 => "00000000000000000011110011110001",
			3900 => "0000000001000000000110101000000100",
			3901 => "00000000000000000011110100001101",
			3902 => "0000001101000000001010001000001000",
			3903 => "0000000101000000000101001000000100",
			3904 => "11111111110101010011110100001101",
			3905 => "00000000000000000011110100001101",
			3906 => "00000000000000000011110100001101",
			3907 => "0000000011000000000111010100001100",
			3908 => "0000001001000000000000111100000100",
			3909 => "00000000000000000011110100101001",
			3910 => "0000001101000000001010001000000100",
			3911 => "11111111110010000011110100101001",
			3912 => "00000000000000000011110100101001",
			3913 => "00000000000000000011110100101001",
			3914 => "0000000101000000001111010000001100",
			3915 => "0000000111000000000001101000000100",
			3916 => "00000000000000000011110101001101",
			3917 => "0000000101000000001101000100000100",
			3918 => "00000000000000000011110101001101",
			3919 => "11111111110110010011110101001101",
			3920 => "0000000111000000000001001000000100",
			3921 => "00000000001000110011110101001101",
			3922 => "00000000000000000011110101001101",
			3923 => "0000001001000000000101011100001100",
			3924 => "0000001110000000000100001000000100",
			3925 => "00000000000000000011110101110001",
			3926 => "0000000000000000001100011100000100",
			3927 => "00000000000011100011110101110001",
			3928 => "00000000000000000011110101110001",
			3929 => "0000000110000000001101111100000100",
			3930 => "11111111110000110011110101110001",
			3931 => "00000000000000000011110101110001",
			3932 => "0000001011000000000101100100001100",
			3933 => "0000001100000000001100110000000100",
			3934 => "00000000000000000011110110011101",
			3935 => "0000001100000000001000000000000100",
			3936 => "11111111111010000011110110011101",
			3937 => "00000000000000000011110110011101",
			3938 => "0000000001000000000000111100001000",
			3939 => "0000000111000000000111010000000100",
			3940 => "00000000001110010011110110011101",
			3941 => "00000000000000000011110110011101",
			3942 => "00000000000000000011110110011101",
			3943 => "0000001010000000000000001000001100",
			3944 => "0000000000000000000010101100000100",
			3945 => "00000000000000000011110111001001",
			3946 => "0000000000000000000001110000000100",
			3947 => "00000000001100100011110111001001",
			3948 => "00000000000000000011110111001001",
			3949 => "0000001010000000000110011000001000",
			3950 => "0000000000000000000001010100000100",
			3951 => "00000000000000000011110111001001",
			3952 => "11111111111100110011110111001001",
			3953 => "00000000000000000011110111001001",
			3954 => "0000001011000000000100010000010000",
			3955 => "0000001011000000001000011000000100",
			3956 => "00000000000000000011110111101101",
			3957 => "0000000110000000000100110100001000",
			3958 => "0000000001000000000000111100000100",
			3959 => "00000000001111010011110111101101",
			3960 => "00000000000000000011110111101101",
			3961 => "00000000000000000011110111101101",
			3962 => "00000000000000000011110111101101",
			3963 => "0000000100000000001111100100010000",
			3964 => "0000000010000000001100010000000100",
			3965 => "00000000000000000011111000010001",
			3966 => "0000000010000000001010000100001000",
			3967 => "0000001000000000001001000100000100",
			3968 => "00000000001111000011111000010001",
			3969 => "00000000000000000011111000010001",
			3970 => "00000000000000000011111000010001",
			3971 => "00000000000000000011111000010001",
			3972 => "0000000111000000001000011000010000",
			3973 => "0000000111000000000001101000000100",
			3974 => "00000000000000000011111000110101",
			3975 => "0000000110000000001101111100000100",
			3976 => "00000000000000000011111000110101",
			3977 => "0000001101000000001001010000000100",
			3978 => "00000000000000000011111000110101",
			3979 => "11111111110011110011111000110101",
			3980 => "00000000000000000011111000110101",
			3981 => "0000000110000000000100110100010000",
			3982 => "0000001010000000001010100000001100",
			3983 => "0000000110000000000111101000000100",
			3984 => "00000000000000000011111001100001",
			3985 => "0000001010000000000000001000000100",
			3986 => "00000000010000000011111001100001",
			3987 => "00000000000000000011111001100001",
			3988 => "00000000000000000011111001100001",
			3989 => "0000001010000000000000001000000100",
			3990 => "00000000000000000011111001100001",
			3991 => "11111111111001000011111001100001",
			3992 => "0000001000000000001001111100001100",
			3993 => "0000001001000000000000111100001000",
			3994 => "0000001111000000000001111100000100",
			3995 => "00000000000000000011111010010101",
			3996 => "00000000001010110011111010010101",
			3997 => "00000000000000000011111010010101",
			3998 => "0000001011000000000101100100000100",
			3999 => "11111111110110100011111010010101",
			4000 => "0000001011000000000100010000000100",
			4001 => "00000000000010110011111010010101",
			4002 => "0000001011000000000111111100000100",
			4003 => "11111111111110000011111010010101",
			4004 => "00000000000000000011111010010101",
			4005 => "0000001010000000000000001000010000",
			4006 => "0000001010000000000100110100000100",
			4007 => "00000000000000000011111011001001",
			4008 => "0000000000000000000001010100001000",
			4009 => "0000001010000000000111101100000100",
			4010 => "00000000000100010011111011001001",
			4011 => "00000000000000000011111011001001",
			4012 => "00000000000000000011111011001001",
			4013 => "0000000000000000000101000100000100",
			4014 => "00000000000000000011111011001001",
			4015 => "0000001010000000000110011000000100",
			4016 => "11111111111100010011111011001001",
			4017 => "00000000000000000011111011001001",
			4018 => "0000000011000000001110110100001100",
			4019 => "0000001001000000000000111100000100",
			4020 => "00000000000000000011111011111101",
			4021 => "0000000001000000000110101000000100",
			4022 => "00000000000000000011111011111101",
			4023 => "11111111111010000011111011111101",
			4024 => "0000000010000000000111010100001100",
			4025 => "0000000111000000001111011100001000",
			4026 => "0000000001000000000000111100000100",
			4027 => "00000000001111110011111011111101",
			4028 => "00000000000000000011111011111101",
			4029 => "00000000000000000011111011111101",
			4030 => "00000000000000000011111011111101",
			4031 => "0000001000000000001001111100001100",
			4032 => "0000000001000000000110101000001000",
			4033 => "0000001110000000000100001000000100",
			4034 => "00000000000000000011111100111001",
			4035 => "00000000001110010011111100111001",
			4036 => "00000000000000000011111100111001",
			4037 => "0000000001000000001001011000001100",
			4038 => "0000000101000000000101001000001000",
			4039 => "0000001111000000000000010000000100",
			4040 => "11111111110000010011111100111001",
			4041 => "00000000000000000011111100111001",
			4042 => "00000000000000000011111100111001",
			4043 => "0000000001000000000000111100000100",
			4044 => "00000000000001100011111100111001",
			4045 => "00000000000000000011111100111001",
			4046 => "0000001001000000001100011000001000",
			4047 => "0000001100000000001100110000000100",
			4048 => "00000000000000000011111101101101",
			4049 => "11111111110110110011111101101101",
			4050 => "0000001001000000001111000000010000",
			4051 => "0000001100000000001000011000001100",
			4052 => "0000000001000000001111001100000100",
			4053 => "00000000000000000011111101101101",
			4054 => "0000001100000000000110000100000100",
			4055 => "00000000000000000011111101101101",
			4056 => "00000000001100100011111101101101",
			4057 => "00000000000000000011111101101101",
			4058 => "00000000000000000011111101101101",
			4059 => "0000001110000000001110101000001000",
			4060 => "0000001000000000001001111100000100",
			4061 => "00000000000000000011111110100001",
			4062 => "11111111110110010011111110100001",
			4063 => "0000000001000000000101011100010000",
			4064 => "0000000111000000000111010000001100",
			4065 => "0000000110000000001010011000001000",
			4066 => "0000001100000000000110000100000100",
			4067 => "00000000000000000011111110100001",
			4068 => "00000000010101000011111110100001",
			4069 => "00000000000000000011111110100001",
			4070 => "00000000000000000011111110100001",
			4071 => "00000000000000000011111110100001",
			4072 => "0000000001000000000110101000000100",
			4073 => "00000000000000000011111111001101",
			4074 => "0000001101000000001010001000010000",
			4075 => "0000001100000000001100110000000100",
			4076 => "00000000000000000011111111001101",
			4077 => "0000001100000000001001001000001000",
			4078 => "0000000111000000001111011100000100",
			4079 => "11111111101110100011111111001101",
			4080 => "00000000000000000011111111001101",
			4081 => "00000000000000000011111111001101",
			4082 => "00000000000000000011111111001101",
			4083 => "0000000011000000001110110100001100",
			4084 => "0000001101000000001010011100000100",
			4085 => "00000000000000000100000000001001",
			4086 => "0000000001000000000110101000000100",
			4087 => "00000000000000000100000000001001",
			4088 => "11111111111010110100000000001001",
			4089 => "0000000001000000001111001100000100",
			4090 => "00000000000000000100000000001001",
			4091 => "0000001011000000000101110100001100",
			4092 => "0000000001000000000000111100001000",
			4093 => "0000000110000000001011001100000100",
			4094 => "00000000010100100100000000001001",
			4095 => "00000000000000000100000000001001",
			4096 => "00000000000000000100000000001001",
			4097 => "00000000000000000100000000001001",
			4098 => "0000001011000000000101100100010000",
			4099 => "0000000010000000000000110100000100",
			4100 => "00000000000000000100000001001101",
			4101 => "0000001100000000001000000000001000",
			4102 => "0000000111000000001000011000000100",
			4103 => "11111111110111100100000001001101",
			4104 => "00000000000000000100000001001101",
			4105 => "00000000000000000100000001001101",
			4106 => "0000000110000000001101111100000100",
			4107 => "00000000000000000100000001001101",
			4108 => "0000000001000000001101111100001100",
			4109 => "0000000101000000001100100100000100",
			4110 => "00000000000000000100000001001101",
			4111 => "0000000110000000000101010000000100",
			4112 => "00000000001101100100000001001101",
			4113 => "00000000000000000100000001001101",
			4114 => "00000000000000000100000001001101",
			4115 => "0000000011000000001100010000010100",
			4116 => "0000001001000000000000111100001100",
			4117 => "0000000000000000000011101000001000",
			4118 => "0000001110000000000100001000000100",
			4119 => "00000000000000000100000010011001",
			4120 => "00000000001011000100000010011001",
			4121 => "00000000000000000100000010011001",
			4122 => "0000000001000000000110101000000100",
			4123 => "00000000000000000100000010011001",
			4124 => "11111111110100010100000010011001",
			4125 => "0000000001000000001111001100000100",
			4126 => "00000000000000000100000010011001",
			4127 => "0000000001000000001101111100001100",
			4128 => "0000000101000000001110101000000100",
			4129 => "00000000000000000100000010011001",
			4130 => "0000001010000000000001010000000100",
			4131 => "00000000001101100100000010011001",
			4132 => "00000000000000000100000010011001",
			4133 => "00000000000000000100000010011001",
			4134 => "0000001110000000001010001000010100",
			4135 => "0000001010000000000111101100010000",
			4136 => "0000000001000000000110101000001000",
			4137 => "0000001110000000000100001000000100",
			4138 => "00000000000000000100000011100101",
			4139 => "00000000010010100100000011100101",
			4140 => "0000000110000000000000111100000100",
			4141 => "11111111111001100100000011100101",
			4142 => "00000000000000000100000011100101",
			4143 => "11111111100000000100000011100101",
			4144 => "0000001001000000000100111100010000",
			4145 => "0000000111000000001000011000001100",
			4146 => "0000000111000000001011000000000100",
			4147 => "00000000000000000100000011100101",
			4148 => "0000001011000000000100000100000100",
			4149 => "00000000000000000100000011100101",
			4150 => "00000000011101110100000011100101",
			4151 => "00000000000000000100000011100101",
			4152 => "00000000000000000100000011100101",
			4153 => "0000000011000000001010000100011100",
			4154 => "0000001100000000001100110000010000",
			4155 => "0000001110000000000100001000000100",
			4156 => "00000000000000000100000100111001",
			4157 => "0000001100000000000100000000000100",
			4158 => "00000000000000000100000100111001",
			4159 => "0000001110000000000101110000000100",
			4160 => "00000000010000000100000100111001",
			4161 => "00000000000000000100000100111001",
			4162 => "0000001100000000001001110100001000",
			4163 => "0000001110000000001100010000000100",
			4164 => "11111111101111100100000100111001",
			4165 => "00000000000000000100000100111001",
			4166 => "00000000000000000100000100111001",
			4167 => "0000001100000000001011011100001100",
			4168 => "0000001100000000000111001000000100",
			4169 => "00000000000000000100000100111001",
			4170 => "0000001110000000000000010100000100",
			4171 => "00000000000110110100000100111001",
			4172 => "00000000000000000100000100111001",
			4173 => "00000000000000000100000100111001",
			4174 => "0000000111000000000110000100001100",
			4175 => "0000001111000000001010111100000100",
			4176 => "00000000000000000100000101111101",
			4177 => "0000000101000000001010011100000100",
			4178 => "11111111101111110100000101111101",
			4179 => "00000000000000000100000101111101",
			4180 => "0000001001000000001111000000010100",
			4181 => "0000000111000000000111010000010000",
			4182 => "0000000000000000001100000100001100",
			4183 => "0000000101000000001111010000001000",
			4184 => "0000001111000000001001001000000100",
			4185 => "00000000000000000100000101111101",
			4186 => "00000000010100110100000101111101",
			4187 => "00000000000000000100000101111101",
			4188 => "00000000000000000100000101111101",
			4189 => "00000000000000000100000101111101",
			4190 => "00000000000000000100000101111101",
			4191 => "0000000001000000001111001100010100",
			4192 => "0000001100000000001100110000010000",
			4193 => "0000000111000000001101100000000100",
			4194 => "00000000000000000100000111001001",
			4195 => "0000001110000000000100001000000100",
			4196 => "00000000000000000100000111001001",
			4197 => "0000000000000000000101000100000100",
			4198 => "00000000001000100100000111001001",
			4199 => "00000000000000000100000111001001",
			4200 => "11111111011110100100000111001001",
			4201 => "0000000001000000000000111100010000",
			4202 => "0000000111000000001111011100001100",
			4203 => "0000001101000000000010110100000100",
			4204 => "00000000000000000100000111001001",
			4205 => "0000001100000000000000001100000100",
			4206 => "00000000000000000100000111001001",
			4207 => "00000000011000100100000111001001",
			4208 => "00000000000000000100000111001001",
			4209 => "00000000000000000100000111001001",
			4210 => "0000001011000000000010001000011100",
			4211 => "0000000000000000000110011100010000",
			4212 => "0000001001000000000000111100001000",
			4213 => "0000001110000000000100001000000100",
			4214 => "00000000000000000100001000100101",
			4215 => "00000000010000100100001000100101",
			4216 => "0000001110000000000101100100000100",
			4217 => "11111111111011110100001000100101",
			4218 => "00000000000000000100001000100101",
			4219 => "0000000011000000001100000000001000",
			4220 => "0000000101000000001100100100000100",
			4221 => "11111111011111010100001000100101",
			4222 => "00000000000000000100001000100101",
			4223 => "00000000000000000100001000100101",
			4224 => "0000000111000000000111010000010000",
			4225 => "0000000001000000000101011100001100",
			4226 => "0000001100000000001011000000000100",
			4227 => "00000000000000000100001000100101",
			4228 => "0000001100000000001001110100000100",
			4229 => "00000000011110100100001000100101",
			4230 => "00000000000000000100001000100101",
			4231 => "00000000000000000100001000100101",
			4232 => "00000000000000000100001000100101",
			4233 => "0000000001000000000000111100011100",
			4234 => "0000001110000000001110101000001000",
			4235 => "0000000110000000000001000100000100",
			4236 => "00000000000000000100001001100001",
			4237 => "11111111111111010100001001100001",
			4238 => "0000000111000000001000011000010000",
			4239 => "0000001001000000000100111100001100",
			4240 => "0000001101000000001001011100001000",
			4241 => "0000000110000000001100011000000100",
			4242 => "00000000101101000100001001100001",
			4243 => "00000000000000000100001001100001",
			4244 => "00000000000000000100001001100001",
			4245 => "00000000000000000100001001100001",
			4246 => "00000000000000000100001001100001",
			4247 => "00000000000000000100001001100001",
			4248 => "0000000101000000000101001000010000",
			4249 => "0000000010000000000000110100000100",
			4250 => "00000000000000000100001010101101",
			4251 => "0000000001000000001001011000001000",
			4252 => "0000001100000000001001110100000100",
			4253 => "11111111110110000100001010101101",
			4254 => "00000000000000000100001010101101",
			4255 => "00000000000000000100001010101101",
			4256 => "0000001011000000000100010000000100",
			4257 => "00000000000000000100001010101101",
			4258 => "0000000110000000000101010000010000",
			4259 => "0000001100000000001011000000000100",
			4260 => "00000000000000000100001010101101",
			4261 => "0000000001000000001101111100001000",
			4262 => "0000000001000000001101011100000100",
			4263 => "00000000000000000100001010101101",
			4264 => "00000000010110010100001010101101",
			4265 => "00000000000000000100001010101101",
			4266 => "00000000000000000100001010101101",
			4267 => "0000001100000000001100110000010100",
			4268 => "0000001110000000000100001000000100",
			4269 => "00000000000000000100001100001001",
			4270 => "0000001001000000001101111100001100",
			4271 => "0000001100000000000100000000000100",
			4272 => "00000000000000000100001100001001",
			4273 => "0000001001000000001011101000000100",
			4274 => "00000000000000000100001100001001",
			4275 => "00000000010011000100001100001001",
			4276 => "00000000000000000100001100001001",
			4277 => "0000000011000000001010000100001100",
			4278 => "0000001100000000001001110100001000",
			4279 => "0000001110000000001100010000000100",
			4280 => "11111111101100110100001100001001",
			4281 => "00000000000000000100001100001001",
			4282 => "00000000000000000100001100001001",
			4283 => "0000001001000000001000010000001100",
			4284 => "0000001001000000001100011000000100",
			4285 => "00000000000000000100001100001001",
			4286 => "0000001100000000001000011000000100",
			4287 => "00000000010000110100001100001001",
			4288 => "00000000000000000100001100001001",
			4289 => "00000000000000000100001100001001",
			4290 => "0000000011000000001010000100011100",
			4291 => "0000001010000000000000001000001100",
			4292 => "0000000010000000001110010000001000",
			4293 => "0000000101000000001110101000000100",
			4294 => "11111111111100100100001101110101",
			4295 => "00000000000000000100001101110101",
			4296 => "00000000000000000100001101110101",
			4297 => "0000001111000000001111010100001100",
			4298 => "0000000000000000000101000100000100",
			4299 => "00000000000000000100001101110101",
			4300 => "0000000110000000001101111100000100",
			4301 => "00000000000000000100001101110101",
			4302 => "11111111011100110100001101110101",
			4303 => "00000000000000000100001101110101",
			4304 => "0000001100000000001001001000010000",
			4305 => "0000000000000000001011010100001100",
			4306 => "0000000111000000001000011000000100",
			4307 => "00000000000000000100001101110101",
			4308 => "0000000001000000000101011100000100",
			4309 => "00000000011110000100001101110101",
			4310 => "00000000000000000100001101110101",
			4311 => "00000000000000000100001101110101",
			4312 => "0000001011000000000111111100001000",
			4313 => "0000000111000000000001101000000100",
			4314 => "00000000000000000100001101110101",
			4315 => "11111111110110110100001101110101",
			4316 => "00000000000000000100001101110101",
			4317 => "0000000101000000001111010000100100",
			4318 => "0000000000000000000101000100010100",
			4319 => "0000001111000000001001001000001000",
			4320 => "0000000001000000001001111000000100",
			4321 => "00000000000000000100001111100001",
			4322 => "11111111110010110100001111100001",
			4323 => "0000000001000000001101101000001000",
			4324 => "0000001011000000000100001000000100",
			4325 => "00000000000000000100001111100001",
			4326 => "00000000010101100100001111100001",
			4327 => "00000000000000000100001111100001",
			4328 => "0000001101000000001010001000001100",
			4329 => "0000000101000000001100100100000100",
			4330 => "00000000000000000100001111100001",
			4331 => "0000001101000000000010011100000100",
			4332 => "00000000000000000100001111100001",
			4333 => "11111111100101000100001111100001",
			4334 => "00000000000000000100001111100001",
			4335 => "0000001010000000000001010000010000",
			4336 => "0000001011000000000010001000000100",
			4337 => "00000000000000000100001111100001",
			4338 => "0000000111000000001000011000000100",
			4339 => "00000000000000000100001111100001",
			4340 => "0000001001000000001010100000000100",
			4341 => "00000000001111110100001111100001",
			4342 => "00000000000000000100001111100001",
			4343 => "00000000000000000100001111100001",
			4344 => "0000000101000000001100100100011100",
			4345 => "0000000000000000000110011100001100",
			4346 => "0000001111000000001010011100000100",
			4347 => "00000000000000000100010001000101",
			4348 => "0000001111000000001110101000000100",
			4349 => "00000000000011110100010001000101",
			4350 => "00000000000000000100010001000101",
			4351 => "0000001111000000001100010000001100",
			4352 => "0000001101000000000101110000001000",
			4353 => "0000001000000000000111110100000100",
			4354 => "00000000000000000100010001000101",
			4355 => "11111111001100010100010001000101",
			4356 => "00000000000000000100010001000101",
			4357 => "00000000000000000100010001000101",
			4358 => "0000001010000000000001010000010100",
			4359 => "0000000001000000001101111100010000",
			4360 => "0000001100000000000111001000000100",
			4361 => "00000000000000000100010001000101",
			4362 => "0000000011000000001100010000000100",
			4363 => "00000000000000000100010001000101",
			4364 => "0000000110000000001000010000000100",
			4365 => "00000000010110100100010001000101",
			4366 => "00000000000000000100010001000101",
			4367 => "00000000000000000100010001000101",
			4368 => "00000000000000000100010001000101",
			4369 => "0000000101000000001111010000011100",
			4370 => "0000001100000000001011000000010000",
			4371 => "0000000000000000001100000100001100",
			4372 => "0000001010000000001101011000000100",
			4373 => "00000000000000000100010010101001",
			4374 => "0000001100000000000011011100000100",
			4375 => "00000000000000000100010010101001",
			4376 => "00000000010100000100010010101001",
			4377 => "00000000000000000100010010101001",
			4378 => "0000001000000000000111110100000100",
			4379 => "00000000000000000100010010101001",
			4380 => "0000000000000000001011010100000100",
			4381 => "11111111111001100100010010101001",
			4382 => "00000000000000000100010010101001",
			4383 => "0000000110000000000101010000010100",
			4384 => "0000001100000000001011000000000100",
			4385 => "00000000000000000100010010101001",
			4386 => "0000001001000000001010100000001100",
			4387 => "0000001010000000000001010000001000",
			4388 => "0000001011000000000010001000000100",
			4389 => "00000000000000000100010010101001",
			4390 => "00000000001110110100010010101001",
			4391 => "00000000000000000100010010101001",
			4392 => "00000000000000000100010010101001",
			4393 => "00000000000000000100010010101001",
			4394 => "0000000111000000001000000000011100",
			4395 => "0000000010000000000000110100010100",
			4396 => "0000000001000000000110101000010000",
			4397 => "0000000010000000000100001000000100",
			4398 => "00000000000000000100010100011101",
			4399 => "0000001100000000000100000000000100",
			4400 => "00000000000000000100010100011101",
			4401 => "0000000100000000000111001000000100",
			4402 => "00000000000000000100010100011101",
			4403 => "00000000010111110100010100011101",
			4404 => "00000000000000000100010100011101",
			4405 => "0000001100000000000100011000000100",
			4406 => "11111111100011110100010100011101",
			4407 => "00000000000000000100010100011101",
			4408 => "0000000011000000001111010100010100",
			4409 => "0000001100000000001011000000001000",
			4410 => "0000000001000000001001011000000100",
			4411 => "00000000010011100100010100011101",
			4412 => "00000000000000000100010100011101",
			4413 => "0000001000000000000111110100000100",
			4414 => "00000000000000000100010100011101",
			4415 => "0000000111000000000110100100000100",
			4416 => "00000000000000000100010100011101",
			4417 => "11111111110001000100010100011101",
			4418 => "0000001001000000000100111100001000",
			4419 => "0000000111000000001111011100000100",
			4420 => "00000000100110100100010100011101",
			4421 => "00000000000000000100010100011101",
			4422 => "00000000000000000100010100011101",
			4423 => "0000000011000000001000011000001000",
			4424 => "0000000110000000001101011100000100",
			4425 => "00000000000000000100010101100001",
			4426 => "11111111110111110100010101100001",
			4427 => "0000001010000000000000001000011000",
			4428 => "0000000110000000000100110100010100",
			4429 => "0000000110000000000000111100000100",
			4430 => "00000000000000000100010101100001",
			4431 => "0000001011000000000100001000000100",
			4432 => "00000000000000000100010101100001",
			4433 => "0000001111000000001010011100000100",
			4434 => "00000000000000000100010101100001",
			4435 => "0000000001000000000000111100000100",
			4436 => "00000000011100010100010101100001",
			4437 => "00000000000000000100010101100001",
			4438 => "00000000000000000100010101100001",
			4439 => "00000000000000000100010101100001",
			4440 => "0000001010000000000000001000010100",
			4441 => "0000001001000000000101011100001100",
			4442 => "0000000001000000000110101000001000",
			4443 => "0000001110000000000100001000000100",
			4444 => "00000000000000000100010111001101",
			4445 => "00000000010101010100010111001101",
			4446 => "00000000000000000100010111001101",
			4447 => "0000000010000000001101000100000100",
			4448 => "11111111111101110100010111001101",
			4449 => "00000000000001100100010111001101",
			4450 => "0000000011000000001010000100001100",
			4451 => "0000000001000000000000111100001000",
			4452 => "0000000010000000001010000100000100",
			4453 => "11111111110001100100010111001101",
			4454 => "00000000000000000100010111001101",
			4455 => "00000000000000000100010111001101",
			4456 => "0000001100000000001011000000000100",
			4457 => "00000000000000000100010111001101",
			4458 => "0000000001000000001101111100010000",
			4459 => "0000000111000000000001101000000100",
			4460 => "00000000000000000100010111001101",
			4461 => "0000000001000000001111001100000100",
			4462 => "00000000000000000100010111001101",
			4463 => "0000000101000000000010011100000100",
			4464 => "00000000010011100100010111001101",
			4465 => "00000000000000000100010111001101",
			4466 => "00000000000000000100010111001101",
			4467 => "0000000101000000001111010000100000",
			4468 => "0000000000000000000101000100011000",
			4469 => "0000001100000000001000000000010100",
			4470 => "0000001010000000001101011000000100",
			4471 => "00000000000000000100011000110001",
			4472 => "0000001100000000000011011100000100",
			4473 => "00000000000000000100011000110001",
			4474 => "0000001010000000000000001000001000",
			4475 => "0000001100000000001011000000000100",
			4476 => "00000000001100010100011000110001",
			4477 => "00000000000000000100011000110001",
			4478 => "00000000000000000100011000110001",
			4479 => "00000000000000000100011000110001",
			4480 => "0000001010000000000000001000000100",
			4481 => "00000000000000000100011000110001",
			4482 => "11111111111010100100011000110001",
			4483 => "0000001010000000000001010000010000",
			4484 => "0000001100000000001011000000000100",
			4485 => "00000000000000000100011000110001",
			4486 => "0000000001000000001101111100001000",
			4487 => "0000000111000000001000011000000100",
			4488 => "00000000000000000100011000110001",
			4489 => "00000000010000000100011000110001",
			4490 => "00000000000000000100011000110001",
			4491 => "00000000000000000100011000110001",
			4492 => "0000000000000000000001010100101100",
			4493 => "0000001110000000001000011000001100",
			4494 => "0000000001000000000110101000001000",
			4495 => "0000001110000000000100001000000100",
			4496 => "00000000000000000100011010010101",
			4497 => "00000000010010010100011010010101",
			4498 => "11111110111001100100011010010101",
			4499 => "0000001100000000001000000000010100",
			4500 => "0000000110000000000100110100010000",
			4501 => "0000000110000000000000111100000100",
			4502 => "00000000000000000100011010010101",
			4503 => "0000001001000000000100111100001000",
			4504 => "0000001110000000000101100100000100",
			4505 => "00000000000000000100011010010101",
			4506 => "00000000011101100100011010010101",
			4507 => "00000000000000000100011010010101",
			4508 => "00000000000000000100011010010101",
			4509 => "0000000010000000001110110100000100",
			4510 => "00000000000000000100011010010101",
			4511 => "0000000010000000001100010000000100",
			4512 => "11111111110111100100011010010101",
			4513 => "00000000000000000100011010010101",
			4514 => "0000000110000000001101111100000100",
			4515 => "00000000000000000100011010010101",
			4516 => "11111111011001100100011010010101",
			4517 => "0000000011000000001000001100101100",
			4518 => "0000001000000000001000100100100100",
			4519 => "0000001100000000001100110000010000",
			4520 => "0000000001000000000111100100001100",
			4521 => "0000001111000000000001111100000100",
			4522 => "00000000000000000100011100001001",
			4523 => "0000000001000000000010001100000100",
			4524 => "00000000000000000100011100001001",
			4525 => "00000000010011110100011100001001",
			4526 => "00000000000000000100011100001001",
			4527 => "0000000011000000001100010000001100",
			4528 => "0000000001000000000110101000000100",
			4529 => "00000000000000000100011100001001",
			4530 => "0000001000000000000100101100000100",
			4531 => "11111111011011010100011100001001",
			4532 => "00000000000000000100011100001001",
			4533 => "0000000001000000001001011000000100",
			4534 => "00000000010111100100011100001001",
			4535 => "00000000000000000100011100001001",
			4536 => "0000001111000000001111100100000100",
			4537 => "11111111101111000100011100001001",
			4538 => "00000000000000000100011100001001",
			4539 => "0000000110000000001000010000001100",
			4540 => "0000001100000000001011000000000100",
			4541 => "00000000000000000100011100001001",
			4542 => "0000000001000000001101111100000100",
			4543 => "00000000011001110100011100001001",
			4544 => "00000000000000000100011100001001",
			4545 => "00000000000000000100011100001001",
			4546 => "0000000110000000001001011000010000",
			4547 => "0000000001000000000110101000001100",
			4548 => "0000001110000000000100001000000100",
			4549 => "00000000000000000100011110000101",
			4550 => "0000000111000000001101100000000100",
			4551 => "00000000000000000100011110000101",
			4552 => "00000000011000010100011110000101",
			4553 => "00000000000000000100011110000101",
			4554 => "0000000101000000000101001000011100",
			4555 => "0000001000000000000111110100000100",
			4556 => "00000000000000000100011110000101",
			4557 => "0000000011000000001100010000001000",
			4558 => "0000001010000000000111101100000100",
			4559 => "00000000000000000100011110000101",
			4560 => "11111111010000100100011110000101",
			4561 => "0000001010000000000000001000000100",
			4562 => "00000000000000000100011110000101",
			4563 => "0000001110000000001001100000000100",
			4564 => "00000000000000000100011110000101",
			4565 => "0000000010000000001000100000000100",
			4566 => "11111111110010010100011110000101",
			4567 => "00000000000000000100011110000101",
			4568 => "0000000111000000001000011000001100",
			4569 => "0000000001000000000000111100001000",
			4570 => "0000001000000000001000100100000100",
			4571 => "00000000000000000100011110000101",
			4572 => "00000000100011000100011110000101",
			4573 => "00000000000000000100011110000101",
			4574 => "0000001101000000000110010000000100",
			4575 => "11111111111110010100011110000101",
			4576 => "00000000000000000100011110000101",
			4577 => "0000001011000000000010001000110000",
			4578 => "0000001010000000000111101100100000",
			4579 => "0000000000000000001010100100010000",
			4580 => "0000000001000000000110101000001100",
			4581 => "0000000010000000000100001000000100",
			4582 => "00000000000000000100100000001001",
			4583 => "0000000111000000001101100000000100",
			4584 => "00000000000000000100100000001001",
			4585 => "00000000001111010100100000001001",
			4586 => "00000000000000000100100000001001",
			4587 => "0000001010000000000100111100000100",
			4588 => "11111111111000110100100000001001",
			4589 => "0000001111000000000010001000000100",
			4590 => "00000000000000000100100000001001",
			4591 => "0000000110000000001101111100000100",
			4592 => "00000000000110010100100000001001",
			4593 => "00000000000000000100100000001001",
			4594 => "0000000011000000001100000000001100",
			4595 => "0000000000000000000110011100000100",
			4596 => "00000000000000000100100000001001",
			4597 => "0000000101000000001100100100000100",
			4598 => "11111111100000010100100000001001",
			4599 => "00000000000000000100100000001001",
			4600 => "00000000000000000100100000001001",
			4601 => "0000000111000000000111010000010000",
			4602 => "0000000001000000000101011100001100",
			4603 => "0000001100000000001011000000000100",
			4604 => "00000000000000000100100000001001",
			4605 => "0000001100000000001001110100000100",
			4606 => "00000000011101100100100000001001",
			4607 => "00000000000000000100100000001001",
			4608 => "00000000000000000100100000001001",
			4609 => "00000000000000000100100000001001",
			4610 => "0000000000000000000001010100110100",
			4611 => "0000000101000000001100100100100100",
			4612 => "0000000001000000001101011100010000",
			4613 => "0000001100000000000100011000001100",
			4614 => "0000000010000000000100001000000100",
			4615 => "00000000000000000100100010000101",
			4616 => "0000001010000000000111101100000100",
			4617 => "00000000001100100100100010000101",
			4618 => "00000000000000000100100010000101",
			4619 => "00000000000000000100100010000101",
			4620 => "0000001001000000001101011000000100",
			4621 => "00000000000000000100100010000101",
			4622 => "0000000010000000001001100000001100",
			4623 => "0000001100000000000100001000000100",
			4624 => "00000000000000000100100010000101",
			4625 => "0000001100000000001000000000000100",
			4626 => "11111111110010010100100010000101",
			4627 => "00000000000000000100100010000101",
			4628 => "00000000000000000100100010000101",
			4629 => "0000000101000000001111010000001100",
			4630 => "0000001100000000000100011000000100",
			4631 => "00000000000000000100100010000101",
			4632 => "0000001001000000000100111100000100",
			4633 => "00000000011000110100100010000101",
			4634 => "00000000000000000100100010000101",
			4635 => "00000000000000000100100010000101",
			4636 => "0000001111000000000110001100001000",
			4637 => "0000001010000000000000001000000100",
			4638 => "00000000000000000100100010000101",
			4639 => "11111111101101110100100010000101",
			4640 => "00000000000000000100100010000101",
			4641 => "0000000101000000000111100000110100",
			4642 => "0000000110000000001101111100100000",
			4643 => "0000001110000000000110100100001000",
			4644 => "0000000110000000001111001100000100",
			4645 => "00000000000000000100100100101001",
			4646 => "11111111101100000100100100101001",
			4647 => "0000001100000000001110001100010000",
			4648 => "0000001011000000000100001000000100",
			4649 => "00000000000000000100100100101001",
			4650 => "0000001111000000001010011100000100",
			4651 => "00000000000000000100100100101001",
			4652 => "0000000111000000001100101000000100",
			4653 => "00000000011111100100100100101001",
			4654 => "00000000000000000100100100101001",
			4655 => "0000000101000000001001010100000100",
			4656 => "11111111101111000100100100101001",
			4657 => "00000000001101000100100100101001",
			4658 => "0000000011000000001100000000010000",
			4659 => "0000000000000000001100011100000100",
			4660 => "00000000000000000100100100101001",
			4661 => "0000000101000000001100100100001000",
			4662 => "0000001101000000000010011100000100",
			4663 => "11111111000000000100100100101001",
			4664 => "00000000000000000100100100101001",
			4665 => "00000000000000000100100100101001",
			4666 => "00000000000000000100100100101001",
			4667 => "0000000110000000001101111100001100",
			4668 => "0000000010000000001110110100000100",
			4669 => "00000000001101110100100100101001",
			4670 => "0000001001000000001111000000000100",
			4671 => "11111111101110000100100100101001",
			4672 => "00000000000000000100100100101001",
			4673 => "0000000111000000001000011000001000",
			4674 => "0000001001000000000100111100000100",
			4675 => "00000000111001100100100100101001",
			4676 => "00000000000000000100100100101001",
			4677 => "0000000011000000001000100000000100",
			4678 => "11111111111101110100100100101001",
			4679 => "0000000011000000000010100100000100",
			4680 => "00000000000110010100100100101001",
			4681 => "00000000000000000100100100101001",
			4682 => "0000001110000000001010001000011100",
			4683 => "0000000000000000001100011100011000",
			4684 => "0000001010000000000100111100010000",
			4685 => "0000000101000000000001101000001100",
			4686 => "0000000011000000000110100100000100",
			4687 => "00000000000000000100100111000101",
			4688 => "0000000110000000000000111100000100",
			4689 => "00000000001111010100100111000101",
			4690 => "00000000000000000100100111000101",
			4691 => "11111111011000110100100111000101",
			4692 => "0000001111000000000010001000000100",
			4693 => "00000000000000000100100111000101",
			4694 => "00000000010110110100100111000101",
			4695 => "11111110101101100100100111000101",
			4696 => "0000001001000000000100111100100100",
			4697 => "0000001100000000001000000000001100",
			4698 => "0000000110000000000100110100001000",
			4699 => "0000000011000000001110110100000100",
			4700 => "00000000000000000100100111000101",
			4701 => "00000000110010110100100111000101",
			4702 => "00000000000000000100100111000101",
			4703 => "0000001110000000001100010000001100",
			4704 => "0000000000000000000101000100000100",
			4705 => "00000000001011110100100111000101",
			4706 => "0000001011000000000101110100000100",
			4707 => "11111111001111010100100111000101",
			4708 => "00000000000000000100100111000101",
			4709 => "0000001001000000001101011000000100",
			4710 => "00000000000000000100100111000101",
			4711 => "0000001100000000001001110100000100",
			4712 => "00000000100110000100100111000101",
			4713 => "00000000000000000100100111000101",
			4714 => "0000001101000000001010001000000100",
			4715 => "11111111101101000100100111000101",
			4716 => "0000000011000000001000001100000100",
			4717 => "00000000000000000100100111000101",
			4718 => "0000000101000000001111010000000100",
			4719 => "00000000000000000100100111000101",
			4720 => "00000000001100000100100111000101",
			4721 => "0000001000000000000110011100110100",
			4722 => "0000000001000000000000111100101100",
			4723 => "0000000011000000000111010100100000",
			4724 => "0000000000000000000001010100010100",
			4725 => "0000001111000000001100000000010000",
			4726 => "0000000011000000001110110100001000",
			4727 => "0000001000000000000111110100000100",
			4728 => "00000000011011110100101001000001",
			4729 => "11111111010001010100101001000001",
			4730 => "0000001001000000000100111100000100",
			4731 => "00000001001010000100101001000001",
			4732 => "00000000000000000100101001000001",
			4733 => "00000000000000000100101001000001",
			4734 => "0000000001000000001001011000001000",
			4735 => "0000001011000000000100000100000100",
			4736 => "11111111101111010100101001000001",
			4737 => "00000000010000000100101001000001",
			4738 => "11111111000101000100101001000001",
			4739 => "0000000010000000001100000000000100",
			4740 => "00000000000000000100101001000001",
			4741 => "0000000111000000001111011100000100",
			4742 => "00000001011000110100101001000001",
			4743 => "00000000000000000100101001000001",
			4744 => "0000001001000000000100111100000100",
			4745 => "00000000000000000100101001000001",
			4746 => "11111111000001000100101001000001",
			4747 => "0000001101000000000011000000000100",
			4748 => "11111110100001000100101001000001",
			4749 => "0000000111000000000000110100000100",
			4750 => "00000000001001100100101001000001",
			4751 => "00000000000000000100101001000001",
			4752 => "0000000111000000001000011000111000",
			4753 => "0000001011000000000010001000101100",
			4754 => "0000001010000000000111101100011000",
			4755 => "0000001100000000000110000100010000",
			4756 => "0000000000000000001010110000001100",
			4757 => "0000001110000000000100001000000100",
			4758 => "00000000000000000100101011001101",
			4759 => "0000000111000000001101100000000100",
			4760 => "00000000000000000100101011001101",
			4761 => "00000000010000110100101011001101",
			4762 => "00000000000000000100101011001101",
			4763 => "0000000010000000001100100100000100",
			4764 => "11111111110010100100101011001101",
			4765 => "00000000000000000100101011001101",
			4766 => "0000000101000000000001000000010000",
			4767 => "0000001111000000001111100100001100",
			4768 => "0000000111000000001000011000001000",
			4769 => "0000000000000000000110011100000100",
			4770 => "00000000000000000100101011001101",
			4771 => "11111111011100000100101011001101",
			4772 => "00000000000000000100101011001101",
			4773 => "00000000000000000100101011001101",
			4774 => "00000000000000000100101011001101",
			4775 => "0000000111000000000001101000000100",
			4776 => "00000000000000000100101011001101",
			4777 => "0000000001000000000000111100000100",
			4778 => "00000000100010000100101011001101",
			4779 => "00000000000000000100101011001101",
			4780 => "0000001101000000000110010000001100",
			4781 => "0000000000000000000101000100000100",
			4782 => "00000000000000000100101011001101",
			4783 => "0000001011000000001010010100000100",
			4784 => "11111111100010010100101011001101",
			4785 => "00000000000000000100101011001101",
			4786 => "00000000000000000100101011001101",
			4787 => "0000001100000000000011011100001000",
			4788 => "0000000110000000001101011100000100",
			4789 => "00000000000000000100101101001001",
			4790 => "11111111000100010100101101001001",
			4791 => "0000000011000000001000100000101000",
			4792 => "0000001000000000001000100100100000",
			4793 => "0000001011000000000010001000011000",
			4794 => "0000001111000000001100100100001100",
			4795 => "0000001100000000000110000100001000",
			4796 => "0000000110000000001001011000000100",
			4797 => "00000000000000000100101101001001",
			4798 => "00000000011010010100101101001001",
			4799 => "11111111100100100100101101001001",
			4800 => "0000001001000000001111000000001000",
			4801 => "0000000111000000001000011000000100",
			4802 => "00000000110101110100101101001001",
			4803 => "00000000000000000100101101001001",
			4804 => "00000000000000000100101101001001",
			4805 => "0000000001000000000000111100000100",
			4806 => "11111111111011100100101101001001",
			4807 => "00000000000000000100101101001001",
			4808 => "0000001111000000001111100100000100",
			4809 => "11111111100110110100101101001001",
			4810 => "00000000000000000100101101001001",
			4811 => "0000000110000000001000010000001100",
			4812 => "0000001100000000001000000000000100",
			4813 => "00000000000000000100101101001001",
			4814 => "0000000001000000001101111100000100",
			4815 => "00000000100110010100101101001001",
			4816 => "00000000000000000100101101001001",
			4817 => "00000000000000000100101101001001",
			4818 => "0000001101000000001010011100001000",
			4819 => "0000000110000000001101011100000100",
			4820 => "00000000000000000100101110110101",
			4821 => "11111110100011100100101110110101",
			4822 => "0000000001000000000101011100101100",
			4823 => "0000000011000000000111010100100000",
			4824 => "0000001011000000000010001000011000",
			4825 => "0000000110000000000100110100010000",
			4826 => "0000000011000000001100010000001000",
			4827 => "0000000110000000001101111100000100",
			4828 => "00000000011100110100101110110101",
			4829 => "11111111001110110100101110110101",
			4830 => "0000000110000000000100110100000100",
			4831 => "00000001000110010100101110110101",
			4832 => "00000000000000000100101110110101",
			4833 => "0000000011000000000110111100000100",
			4834 => "11111111011101100100101110110101",
			4835 => "00000000000000000100101110110101",
			4836 => "0000000010000000001110110100000100",
			4837 => "00000000000101110100101110110101",
			4838 => "11111110100010110100101110110101",
			4839 => "0000000111000000000111010000001000",
			4840 => "0000001011000000000010001000000100",
			4841 => "00000000000000000100101110110101",
			4842 => "00000001000010100100101110110101",
			4843 => "11111111111011010100101110110101",
			4844 => "11111111000100000100101110110101",
			4845 => "0000001100000000001100110000001100",
			4846 => "0000000000000000001010110000001000",
			4847 => "0000001110000000000100001000000100",
			4848 => "00000000000000000100110001000001",
			4849 => "00000000011000100100110001000001",
			4850 => "00000000000000000100110001000001",
			4851 => "0000000111000000001000000000001100",
			4852 => "0000001100000000001100110000000100",
			4853 => "00000000000000000100110001000001",
			4854 => "0000001100000000000100011000000100",
			4855 => "11111111100111100100110001000001",
			4856 => "00000000000000000100110001000001",
			4857 => "0000000110000000000100110100010000",
			4858 => "0000001100000000001000000000001100",
			4859 => "0000001001000000000100111100001000",
			4860 => "0000001101000000001110101000000100",
			4861 => "00000000000000000100110001000001",
			4862 => "00000000010001000100110001000001",
			4863 => "00000000000000000100110001000001",
			4864 => "00000000000000000100110001000001",
			4865 => "0000001110000000001111010100010000",
			4866 => "0000001100000000001011000000000100",
			4867 => "00000000000000000100110001000001",
			4868 => "0000000010000000001110110100000100",
			4869 => "00000000000000000100110001000001",
			4870 => "0000000101000000000010011100000100",
			4871 => "11111111101101010100110001000001",
			4872 => "00000000000000000100110001000001",
			4873 => "0000001100000000001000000000000100",
			4874 => "00000000000000000100110001000001",
			4875 => "0000001000000000001001101000001000",
			4876 => "0000001000000000001000010100000100",
			4877 => "00000000000000000100110001000001",
			4878 => "00000000001010110100110001000001",
			4879 => "00000000000000000100110001000001",
			4880 => "0000001010000000001010100100101100",
			4881 => "0000000111000000000110000100001100",
			4882 => "0000000110000000001101011100001000",
			4883 => "0000000111000000001101100000000100",
			4884 => "11111111010101110100110011011101",
			4885 => "00000000011000000100110011011101",
			4886 => "11111101111100110100110011011101",
			4887 => "0000001001000000000100111100011100",
			4888 => "0000001100000000001001110100010100",
			4889 => "0000000001000000000110101000000100",
			4890 => "00000111000000010100110011011101",
			4891 => "0000001010000000000100111100001000",
			4892 => "0000000001000000000111100100000100",
			4893 => "00000000111110110100110011011101",
			4894 => "11111110011111010100110011011101",
			4895 => "0000000011000000000111010100000100",
			4896 => "00000001011110100100110011011101",
			4897 => "00000010101010010100110011011101",
			4898 => "0000001000000000001000100100000100",
			4899 => "00000001001101100100110011011101",
			4900 => "11111110100000100100110011011101",
			4901 => "11111110101000100100110011011101",
			4902 => "0000000001000000001111001100000100",
			4903 => "11111110011000100100110011011101",
			4904 => "0000001001000000001101011000010000",
			4905 => "0000000010000000001101101100001000",
			4906 => "0000001110000000000010011100000100",
			4907 => "00000000000000000100110011011101",
			4908 => "00000001101110010100110011011101",
			4909 => "0000000111000000000010110100000100",
			4910 => "00001010110101010100110011011101",
			4911 => "00000000000000000100110011011101",
			4912 => "0000001011000000001001010000001100",
			4913 => "0000000001000000000101011100001000",
			4914 => "0000001000000000001100011100000100",
			4915 => "00000001011011000100110011011101",
			4916 => "11111110110101000100110011011101",
			4917 => "11111110011010000100110011011101",
			4918 => "00000011011011010100110011011101",
			4919 => "0000001101000000001010011100001000",
			4920 => "0000001010000000001100011000000100",
			4921 => "00000000000000000100110101010001",
			4922 => "11111110100011110100110101010001",
			4923 => "0000001001000000000101010000110000",
			4924 => "0000000011000000000111010100100000",
			4925 => "0000001011000000000010001000011000",
			4926 => "0000000000000000000001010100001100",
			4927 => "0000000011000000000111011000001000",
			4928 => "0000000111000000000001101000000100",
			4929 => "00000000100010000100110101010001",
			4930 => "11111111010100000100110101010001",
			4931 => "00000001001011110100110101010001",
			4932 => "0000000011000000001111010100001000",
			4933 => "0000001101000000000100101000000100",
			4934 => "11111111100110010100110101010001",
			4935 => "00000000000000000100110101010001",
			4936 => "00000000000000000100110101010001",
			4937 => "0000000010000000001110110100000100",
			4938 => "00000000001101100100110101010001",
			4939 => "11111110010111110100110101010001",
			4940 => "0000000111000000001111011100001000",
			4941 => "0000001001000000001000010000000100",
			4942 => "00000001010001110100110101010001",
			4943 => "00000000000000000100110101010001",
			4944 => "0000001100000000001001110100000100",
			4945 => "00000000000000000100110101010001",
			4946 => "11111111100101100100110101010001",
			4947 => "11111111000001110100110101010001",
			4948 => "0000001010000000001010100100101100",
			4949 => "0000000111000000000110000100001100",
			4950 => "0000000110000000001101011100001000",
			4951 => "0000000110000000001111001100000100",
			4952 => "11111111011011110100110111101101",
			4953 => "00000000010100010100110111101101",
			4954 => "11111101111111110100110111101101",
			4955 => "0000001001000000000100111100011100",
			4956 => "0000000111000000001111011100010100",
			4957 => "0000001111000000001111010100010000",
			4958 => "0000000000000000000001010100001000",
			4959 => "0000001100000000000011011100000100",
			4960 => "11111111001101010100110111101101",
			4961 => "00000001100011000100110111101101",
			4962 => "0000000111000000001000011000000100",
			4963 => "11111111010001100100110111101101",
			4964 => "00000001000110100100110111101101",
			4965 => "00000011010001000100110111101101",
			4966 => "0000000010000000000010000100000100",
			4967 => "00000000111010100100110111101101",
			4968 => "11111110100011100100110111101101",
			4969 => "11111110101010100100110111101101",
			4970 => "0000000001000000001111001100000100",
			4971 => "11111110011000100100110111101101",
			4972 => "0000000001000000001101011100001100",
			4973 => "0000000101000000001101000100000100",
			4974 => "11111111011011110100110111101101",
			4975 => "0000001100000000000100010000000100",
			4976 => "00000100000010110100110111101101",
			4977 => "00000000000000000100110111101101",
			4978 => "0000001011000000001001010000010000",
			4979 => "0000000001000000000101011100001100",
			4980 => "0000001111000000001011101100000100",
			4981 => "11111110111110000100110111101101",
			4982 => "0000000100000000001000001000000100",
			4983 => "00000001011110000100110111101101",
			4984 => "11111111110100000100110111101101",
			4985 => "11111110011010010100110111101101",
			4986 => "00000010110111000100110111101101",
			4987 => "0000000111000000001101100000000100",
			4988 => "11111110011101000100111001110001",
			4989 => "0000000000000000000110011100011000",
			4990 => "0000000001000000001101011100010000",
			4991 => "0000001100000000000100011000001000",
			4992 => "0000001110000000000100001000000100",
			4993 => "00000000000000000100111001110001",
			4994 => "00000001001101000100111001110001",
			4995 => "0000000010000000000010011100000100",
			4996 => "00000000000000000100111001110001",
			4997 => "00000000010001100100111001110001",
			4998 => "0000000011000000000010000000000100",
			4999 => "11111111001010010100111001110001",
			5000 => "00000001000001100100111001110001",
			5001 => "0000000101000000001110101000001100",
			5002 => "0000001000000000000111110100000100",
			5003 => "00000000000000000100111001110001",
			5004 => "0000001011000000001011011100000100",
			5005 => "11111110100000110100111001110001",
			5006 => "00000000000000000100111001110001",
			5007 => "0000000001000000001111001100000100",
			5008 => "11111110101101110100111001110001",
			5009 => "0000000001000000000000111100001100",
			5010 => "0000000010000000001010000100001000",
			5011 => "0000000111000000001000011000000100",
			5012 => "00000000101100100100111001110001",
			5013 => "11111110110001100100111001110001",
			5014 => "00000001111101010100111001110001",
			5015 => "0000001100000000001011011100000100",
			5016 => "11111110101110010100111001110001",
			5017 => "0000000110000000001001111100000100",
			5018 => "00000000111111110100111001110001",
			5019 => "00000000000000000100111001110001",
			5020 => "0000001010000000001010100101001100",
			5021 => "0000001110000000001110101000100000",
			5022 => "0000000001000000000111100100010000",
			5023 => "0000001110000000001010111000001000",
			5024 => "0000000110000000001111001100000100",
			5025 => "00000001010110000100111100110101",
			5026 => "11111110100011100100111100110101",
			5027 => "0000001100000000000011011100000100",
			5028 => "00000010001110010100111100110101",
			5029 => "00000110011111010100111100110101",
			5030 => "0000001100000000000110000100001100",
			5031 => "0000001011000000000001111100000100",
			5032 => "11111110001111100100111100110101",
			5033 => "0000000100000000000111010000000100",
			5034 => "11111111001011000100111100110101",
			5035 => "00000001011100100100111100110101",
			5036 => "11111110010111100100111100110101",
			5037 => "0000000001000000000000111100100100",
			5038 => "0000000111000000001000011000010100",
			5039 => "0000000100000000001010000100010000",
			5040 => "0000000110000000001101111100001000",
			5041 => "0000001010000000000000001000000100",
			5042 => "00000001110010110100111100110101",
			5043 => "00000001001011100100111100110101",
			5044 => "0000000011000000001100010000000100",
			5045 => "11111100001110100100111100110101",
			5046 => "00000000111100010100111100110101",
			5047 => "00000011011011100100111100110101",
			5048 => "0000001011000000000100010000001000",
			5049 => "0000000000000000000001010100000100",
			5050 => "00000001100000100100111100110101",
			5051 => "11111110000001110100111100110101",
			5052 => "0000001110000000001100010000000100",
			5053 => "11111100001101010100111100110101",
			5054 => "11111110011111100100111100110101",
			5055 => "0000001101000000000011001000000100",
			5056 => "11111110011111100100111100110101",
			5057 => "00000001010011010100111100110101",
			5058 => "0000001010000000000111110100001100",
			5059 => "0000000010000000000110101100000100",
			5060 => "11111110011011100100111100110101",
			5061 => "0000000001000000001110010100000100",
			5062 => "00000100111111100100111100110101",
			5063 => "11111111111110000100111100110101",
			5064 => "0000000101000000001111100100000100",
			5065 => "11111110011001110100111100110101",
			5066 => "0000000010000000001101000000000100",
			5067 => "00000010000101100100111100110101",
			5068 => "11111110100000010100111100110101",
			5069 => "0000001010000000000111110100111100",
			5070 => "0000000001000000000000111100110100",
			5071 => "0000000011000000000111010100101000",
			5072 => "0000000000000000000001010100011100",
			5073 => "0000000101000000000111100000010000",
			5074 => "0000000111000000000001101000001000",
			5075 => "0000000011000000000000110100000100",
			5076 => "00000000000010010100111111000001",
			5077 => "00000000110111100100111111000001",
			5078 => "0000000110000000001101111100000100",
			5079 => "00000000000000000100111111000001",
			5080 => "11111110111110000100111111000001",
			5081 => "0000001000000000001000100100001000",
			5082 => "0000000011000000001100000000000100",
			5083 => "00000000000000000100111111000001",
			5084 => "00000001010010010100111111000001",
			5085 => "00000000000000000100111111000001",
			5086 => "0000000101000000000111100000001000",
			5087 => "0000001101000000001110101100000100",
			5088 => "11111111101101000100111111000001",
			5089 => "00000000010101000100111111000001",
			5090 => "11111111000010000100111111000001",
			5091 => "0000000010000000001100000000000100",
			5092 => "00000000000000000100111111000001",
			5093 => "0000000111000000001111011100000100",
			5094 => "00000001011101010100111111000001",
			5095 => "00000000000000000100111111000001",
			5096 => "0000001001000000000100111100000100",
			5097 => "00000000000000000100111111000001",
			5098 => "11111111000000010100111111000001",
			5099 => "0000001101000000000011000000000100",
			5100 => "11111110100000010100111111000001",
			5101 => "0000000111000000000000110100000100",
			5102 => "00000000001110110100111111000001",
			5103 => "00000000000000000100111111000001",
			5104 => "0000000111000000001101100000000100",
			5105 => "11111110101011110101000001000101",
			5106 => "0000001010000000000111101100010000",
			5107 => "0000000001000000001101011100001100",
			5108 => "0000001110000000000100001000000100",
			5109 => "00000000000000000101000001000101",
			5110 => "0000000100000000001001100000000100",
			5111 => "00000000100111110101000001000101",
			5112 => "00000000000000000101000001000101",
			5113 => "00000000000000000101000001000101",
			5114 => "0000000101000000000101001000011000",
			5115 => "0000000111000000000001101000010000",
			5116 => "0000000111000000001000000000000100",
			5117 => "11111111000010000101000001000101",
			5118 => "0000001000000000001100011100001000",
			5119 => "0000001000000000000111110100000100",
			5120 => "00000000000000000101000001000101",
			5121 => "00000000010010100101000001000101",
			5122 => "00000000000000000101000001000101",
			5123 => "0000000111000000001111011100000100",
			5124 => "11111111000101010101000001000101",
			5125 => "00000000000000000101000001000101",
			5126 => "0000000001000000000000111100010000",
			5127 => "0000001011000000000010001000000100",
			5128 => "00000000000000000101000001000101",
			5129 => "0000000111000000001111011100001000",
			5130 => "0000000011000000001010000100000100",
			5131 => "00000000000000000101000001000101",
			5132 => "00000000111100010101000001000101",
			5133 => "00000000000000000101000001000101",
			5134 => "0000000011000000001111100000000100",
			5135 => "11111111100000010101000001000101",
			5136 => "00000000000011010101000001000101",
			5137 => "0000000000000000001011010100111100",
			5138 => "0000001100000000000001101000111000",
			5139 => "0000001010000000000111101100011000",
			5140 => "0000000010000000001100100100010100",
			5141 => "0000000001000000000111100100001100",
			5142 => "0000001111000000001011000000000100",
			5143 => "11111111010100110101000011100001",
			5144 => "0000000001000000001001111000000100",
			5145 => "00000000000000000101000011100001",
			5146 => "00000001011001000101000011100001",
			5147 => "0000001100000000001100110000000100",
			5148 => "00000000000000000101000011100001",
			5149 => "11111110101011010101000011100001",
			5150 => "00000001011101100101000011100001",
			5151 => "0000000011000000001100010000010000",
			5152 => "0000000110000000001101111100001000",
			5153 => "0000000001000000001111001100000100",
			5154 => "11111111100100010101000011100001",
			5155 => "00000000011110010101000011100001",
			5156 => "0000001100000000000100011000000100",
			5157 => "00000000000000000101000011100001",
			5158 => "11111101011110100101000011100001",
			5159 => "0000001010000000000000001000000100",
			5160 => "00000001010111010101000011100001",
			5161 => "0000000110000000001101111100000100",
			5162 => "11111110110000000101000011100001",
			5163 => "0000000111000000001000011000000100",
			5164 => "11111111101000110101000011100001",
			5165 => "00000000110001000101000011100001",
			5166 => "00000111001001110101000011100001",
			5167 => "0000001011000000000101100100000100",
			5168 => "11111110011001000101000011100001",
			5169 => "0000001011000000001011011100001000",
			5170 => "0000001001000000000100101100000100",
			5171 => "00000001001000110101000011100001",
			5172 => "00000000000000000101000011100001",
			5173 => "0000000101000000001111100100000100",
			5174 => "11111110101000010101000011100001",
			5175 => "00000000000000000101000011100001",
			5176 => "0000001000000000001000100100110100",
			5177 => "0000001110000000001000011000010100",
			5178 => "0000000110000000001101011100001000",
			5179 => "0000001010000000000100110100000100",
			5180 => "11111110101001000101000110110101",
			5181 => "00001000111101010101000110110101",
			5182 => "0000001110000000001011000000000100",
			5183 => "11111110011001100101000110110101",
			5184 => "0000000001000000000111100100000100",
			5185 => "00000101110100000101000110110101",
			5186 => "11111110011101110101000110110101",
			5187 => "0000000001000000000000111100011000",
			5188 => "0000000111000000001101111000000100",
			5189 => "00001001100111010101000110110101",
			5190 => "0000001110000000000111110000000100",
			5191 => "11111110011111100101000110110101",
			5192 => "0000001101000000000111111100001000",
			5193 => "0000000111000000001111011100000100",
			5194 => "00000011111111000101000110110101",
			5195 => "00000010011100110101000110110101",
			5196 => "0000001100000000001000000000000100",
			5197 => "00000100001100100101000110110101",
			5198 => "00000001001100110101000110110101",
			5199 => "0000000110000000001101111100000100",
			5200 => "00000001010011010101000110110101",
			5201 => "11111110011011010101000110110101",
			5202 => "0000000000000000001001101000011000",
			5203 => "0000000001000000000000111100010100",
			5204 => "0000000011000000000000010000010000",
			5205 => "0000001100000000001011000000000100",
			5206 => "00000100010100000101000110110101",
			5207 => "0000001010000000001010100000000100",
			5208 => "11111110011101110101000110110101",
			5209 => "0000000111000000001000011000000100",
			5210 => "00000011011100010101000110110101",
			5211 => "11111110101011100101000110110101",
			5212 => "00001001001111100101000110110101",
			5213 => "11111110011000100101000110110101",
			5214 => "0000001010000000000010101100001100",
			5215 => "0000000100000000001101101100000100",
			5216 => "11111110011001000101000110110101",
			5217 => "0000000001000000001100110100000100",
			5218 => "11111110100100010101000110110101",
			5219 => "00000101001011100101000110110101",
			5220 => "0000001101000000000011000000000100",
			5221 => "11111110010110010101000110110101",
			5222 => "0000001101000000000010010100001100",
			5223 => "0000000101000000001000100000001000",
			5224 => "0000000101000000001111100100000100",
			5225 => "11111111011111010101000110110101",
			5226 => "00000001011101110101000110110101",
			5227 => "11111110110000000101000110110101",
			5228 => "11111110010111100101000110110101",
			5229 => "0000001000000000001001000101001100",
			5230 => "0000000110000000000100110100101000",
			5231 => "0000001110000000001110101000010100",
			5232 => "0000000110000000000001000100010000",
			5233 => "0000001100000000000110000100001100",
			5234 => "0000001110000000000100001000000100",
			5235 => "11111111110010000101001001111001",
			5236 => "0000001001000000000101011100000100",
			5237 => "00000001100000110101001001111001",
			5238 => "00000000011111000101001001111001",
			5239 => "11111111101000100101001001111001",
			5240 => "11111110010110000101001001111001",
			5241 => "0000001001000000000100111100010000",
			5242 => "0000000111000000001111011100001100",
			5243 => "0000000111000000001000011000001000",
			5244 => "0000000111000000000001101000000100",
			5245 => "00000001011100100101001001111001",
			5246 => "00000000000000000101001001111001",
			5247 => "00000001110100000101001001111001",
			5248 => "00000000000000000101001001111001",
			5249 => "11111111100011110101001001111001",
			5250 => "0000000011000000001000001100011100",
			5251 => "0000000100000000000111011000010100",
			5252 => "0000001011000000000110110100001100",
			5253 => "0000001110000000001001100000001000",
			5254 => "0000001000000000001000100100000100",
			5255 => "00000000000000000101001001111001",
			5256 => "11111111000100110101001001111001",
			5257 => "00000000000000000101001001111001",
			5258 => "0000001001000000001111000000000100",
			5259 => "00000001001011100101001001111001",
			5260 => "11111111111101010101001001111001",
			5261 => "0000001100000000000100011000000100",
			5262 => "00000000000000000101001001111001",
			5263 => "11111110101100110101001001111001",
			5264 => "0000001011000000000101110100000100",
			5265 => "00000001011011010101001001111001",
			5266 => "11111111111100100101001001111001",
			5267 => "0000001011000000000101110100000100",
			5268 => "11111110011010000101001001111001",
			5269 => "0000001100000000001001110100001000",
			5270 => "0000000001000000000101011100000100",
			5271 => "00000001111010100101001001111001",
			5272 => "11111111111011000101001001111001",
			5273 => "0000001101000000000011000000000100",
			5274 => "11111110101000100101001001111001",
			5275 => "0000001101000000001111101000000100",
			5276 => "00000000000000000101001001111001",
			5277 => "11111111111101100101001001111001",
			5278 => "0000000000000000000010111101001100",
			5279 => "0000000011000000001010000100110000",
			5280 => "0000000000000000000101000100011100",
			5281 => "0000000010000000001101000100010100",
			5282 => "0000001001000000000000111100001100",
			5283 => "0000001110000000000100001000000100",
			5284 => "00000000000000000101001100010101",
			5285 => "0000000111000000001101100000000100",
			5286 => "00000000000000000101001100010101",
			5287 => "00000000100000010101001100010101",
			5288 => "0000001001000000001110010100000100",
			5289 => "11111111010101000101001100010101",
			5290 => "00000000000000000101001100010101",
			5291 => "0000000110000000001101111100000100",
			5292 => "00000000101101000101001100010101",
			5293 => "00000000000000000101001100010101",
			5294 => "0000001000000000001000100100000100",
			5295 => "00000000000000000101001100010101",
			5296 => "0000001010000000000000001000000100",
			5297 => "00000000000000000101001100010101",
			5298 => "0000001111000000001111010100001000",
			5299 => "0000001100000000001001110100000100",
			5300 => "11111111001001000101001100010101",
			5301 => "00000000000000000101001100010101",
			5302 => "00000000000000000101001100010101",
			5303 => "0000000111000000001111011100001100",
			5304 => "0000001001000000001000010000001000",
			5305 => "0000000110000000000100110100000100",
			5306 => "00000000000000000101001100010101",
			5307 => "00000000111110100101001100010101",
			5308 => "00000000000000000101001100010101",
			5309 => "0000000101000000001110010000000100",
			5310 => "11111111101000110101001100010101",
			5311 => "0000001001000000001010100000001000",
			5312 => "0000000110000000001000010000000100",
			5313 => "00000000011001010101001100010101",
			5314 => "00000000000000000101001100010101",
			5315 => "00000000000000000101001100010101",
			5316 => "11111110111101110101001100010101",
			5317 => "0000001010000000000010101101001100",
			5318 => "0000000001000000000000111101000000",
			5319 => "0000001110000000001110101000100000",
			5320 => "0000000000000000000110011000011100",
			5321 => "0000001100000000001100110000010000",
			5322 => "0000001111000000001011000000001000",
			5323 => "0000000110000000001111001100000100",
			5324 => "00000010011000010101001111011001",
			5325 => "11111110100100100101001111011001",
			5326 => "0000001001000000000101011100000100",
			5327 => "00000100101010000101001111011001",
			5328 => "00000001011100110101001111011001",
			5329 => "0000000111000000001110001100001000",
			5330 => "0000001001000000001011111100000100",
			5331 => "11111111000101110101001111011001",
			5332 => "00000001000110000101001111011001",
			5333 => "11111110011001110101001111011001",
			5334 => "11111101111100000101001111011001",
			5335 => "0000000011000000001000001100011000",
			5336 => "0000000000000000000001010100001100",
			5337 => "0000001001000000000100111100001000",
			5338 => "0000001110000000000010000100000100",
			5339 => "00000001110100000101001111011001",
			5340 => "00000010110111000101001111011001",
			5341 => "11111110111100010101001111011001",
			5342 => "0000001100000000001011000000000100",
			5343 => "00000010100111100101001111011001",
			5344 => "0000000011000000000111010100000100",
			5345 => "11111110100010000101001111011001",
			5346 => "00000000100110110101001111011001",
			5347 => "0000000111000000001000011000000100",
			5348 => "00000100000011010101001111011001",
			5349 => "00000010001110000101001111011001",
			5350 => "0000001001000000000100111100001000",
			5351 => "0000000101000000001001010000000100",
			5352 => "11111110111001100101001111011001",
			5353 => "00000001111111000101001111011001",
			5354 => "11111110011011110101001111011001",
			5355 => "0000001010000000000011101000001100",
			5356 => "0000000100000000001111101000000100",
			5357 => "11111110011101110101001111011001",
			5358 => "0000000000000000001000101100000100",
			5359 => "00000101001010000101001111011001",
			5360 => "11111111011011110101001111011001",
			5361 => "0000000101000000001111100100000100",
			5362 => "11111110011000100101001111011001",
			5363 => "0000000101000000001000100000000100",
			5364 => "00000000011000100101001111011001",
			5365 => "11111110011110010101001111011001",
			5366 => "0000001010000000001010100101010000",
			5367 => "0000001110000000001110101000101100",
			5368 => "0000000110000000001001011000011000",
			5369 => "0000001100000000000110000100010100",
			5370 => "0000001110000000000100001000000100",
			5371 => "11111110101111100101010010100101",
			5372 => "0000000001000000000110101000001000",
			5373 => "0000001100000000001000111000000100",
			5374 => "00000011000010100101010010100101",
			5375 => "00000000000000000101010010100101",
			5376 => "0000001001000000000101011100000100",
			5377 => "11111111000000000101010010100101",
			5378 => "00000000000000000101010010100101",
			5379 => "00001001100100110101010010100101",
			5380 => "0000001011000000000100001000000100",
			5381 => "11111110010011000101010010100101",
			5382 => "0000001100000000000110000100001100",
			5383 => "0000000100000000000111010000000100",
			5384 => "11111111000010100101010010100101",
			5385 => "0000000001000000000111100100000100",
			5386 => "00000001101100000101010010100101",
			5387 => "00000000000000000101010010100101",
			5388 => "11111110011010010101010010100101",
			5389 => "0000001001000000000100111100100000",
			5390 => "0000000111000000001111011100010100",
			5391 => "0000000011000000000111010100010000",
			5392 => "0000000110000000001101111100001000",
			5393 => "0000001101000000000111111100000100",
			5394 => "00000001101111100101010010100101",
			5395 => "00000000011011100101010010100101",
			5396 => "0000000011000000001100010000000100",
			5397 => "11111100101100000101010010100101",
			5398 => "00000000101001110101010010100101",
			5399 => "00000011010010010101010010100101",
			5400 => "0000000111000000001111011100001000",
			5401 => "0000001110000000001100010000000100",
			5402 => "00000001001000100101010010100101",
			5403 => "11111110100001000101010010100101",
			5404 => "11111101100101000101010010100101",
			5405 => "11111110100010100101010010100101",
			5406 => "0000001010000000000111110100001100",
			5407 => "0000000010000000000110101100000100",
			5408 => "11111110011100000101010010100101",
			5409 => "0000000011000000001000100000000100",
			5410 => "00000101010110010101010010100101",
			5411 => "00000001011101100101010010100101",
			5412 => "0000000101000000001111100100000100",
			5413 => "11111110011010000101010010100101",
			5414 => "0000000010000000001101000000000100",
			5415 => "00000001110010100101010010100101",
			5416 => "11111110100001110101010010100101",
			5417 => "0000000111000000001101100000000100",
			5418 => "11111110111000110101010100110001",
			5419 => "0000001010000000000111101100001100",
			5420 => "0000001110000000000100001000000100",
			5421 => "00000000000000000101010100110001",
			5422 => "0000001100000000000100011000000100",
			5423 => "00000000101100010101010100110001",
			5424 => "00000000000000000101010100110001",
			5425 => "0000000101000000000101001000011000",
			5426 => "0000001101000000001010001000010100",
			5427 => "0000001101000000000111111100010000",
			5428 => "0000000011000000001100010000001000",
			5429 => "0000001000000000000111110100000100",
			5430 => "00000000000000000101010100110001",
			5431 => "11111111000101110101010100110001",
			5432 => "0000000001000000001001011000000100",
			5433 => "00000000110100110101010100110001",
			5434 => "11111111111011100101010100110001",
			5435 => "11111110111101110101010100110001",
			5436 => "00000000000000000101010100110001",
			5437 => "0000001011000000000100010000001100",
			5438 => "0000001101000000000111111100000100",
			5439 => "00000000000111100101010100110001",
			5440 => "0000001101000000001010001000000100",
			5441 => "11111111100011010101010100110001",
			5442 => "00000000000000000101010100110001",
			5443 => "0000000111000000000111010000001100",
			5444 => "0000000001000000000000111100001000",
			5445 => "0000001101000000000111111100000100",
			5446 => "00000000000000000101010100110001",
			5447 => "00000000111100110101010100110001",
			5448 => "00000000000000000101010100110001",
			5449 => "0000001101000000001111101000000100",
			5450 => "11111111110101010101010100110001",
			5451 => "00000000000000000101010100110001",
			5452 => "0000001101000000001010011100001000",
			5453 => "0000001010000000001100011000000100",
			5454 => "00000000000000000101010110110101",
			5455 => "11111110100101010101010110110101",
			5456 => "0000000001000000000101011100111000",
			5457 => "0000000011000000000111010100101000",
			5458 => "0000001011000000000010001000100000",
			5459 => "0000000011000000001100010000010000",
			5460 => "0000001010000000000111101100001000",
			5461 => "0000001111000000001010011100000100",
			5462 => "00000000000000000101010110110101",
			5463 => "00000000100101000101010110110101",
			5464 => "0000001000000000000111110100000100",
			5465 => "00000000000000000101010110110101",
			5466 => "11111110111110100101010110110101",
			5467 => "0000000001000000001001011000001000",
			5468 => "0000000111000000001111011100000100",
			5469 => "00000001001011010101010110110101",
			5470 => "00000000000000000101010110110101",
			5471 => "0000000000000000000001010100000100",
			5472 => "00000000001010100101010110110101",
			5473 => "11111111100100010101010110110101",
			5474 => "0000000010000000001110110100000100",
			5475 => "00000000001010000101010110110101",
			5476 => "11111110011101100101010110110101",
			5477 => "0000000111000000000111010000001100",
			5478 => "0000001011000000000010001000000100",
			5479 => "00000000000000000101010110110101",
			5480 => "0000000111000000001111011100000100",
			5481 => "00000001001101110101010110110101",
			5482 => "00000000000000000101010110110101",
			5483 => "11111111110111110101010110110101",
			5484 => "11111111000001000101010110110101",
			5485 => "0000000000000000001100000101010100",
			5486 => "0000001100000000001000000000110100",
			5487 => "0000001110000000001110101000010100",
			5488 => "0000000110000000000001000100010000",
			5489 => "0000001100000000000110000100001100",
			5490 => "0000001110000000000100001000000100",
			5491 => "11111111110000110101011010001001",
			5492 => "0000001001000000000000111100000100",
			5493 => "00000001110101010101011010001001",
			5494 => "00000000011111110101011010001001",
			5495 => "11111111000111100101011010001001",
			5496 => "11111110001110000101011010001001",
			5497 => "0000001010000000000000001000001000",
			5498 => "0000000001000000000000111100000100",
			5499 => "00000001011110100101011010001001",
			5500 => "11111111111011000101011010001001",
			5501 => "0000000011000000001010000100001100",
			5502 => "0000001011000000000000011100000100",
			5503 => "00000000000000000101011010001001",
			5504 => "0000000000000000001100000100000100",
			5505 => "11111110100101010101011010001001",
			5506 => "00000000000000000101011010001001",
			5507 => "0000000000000000000001110000000100",
			5508 => "00000001110010000101011010001001",
			5509 => "0000000101000000000101001000000100",
			5510 => "11111111111010110101011010001001",
			5511 => "00000000000000000101011010001001",
			5512 => "0000000011000000001001100000000100",
			5513 => "11111101110000100101011010001001",
			5514 => "0000000100000000000111011000001000",
			5515 => "0000001010000000000000001000000100",
			5516 => "00000001100110010101011010001001",
			5517 => "00000000000000000101011010001001",
			5518 => "0000001100000000001000000000001000",
			5519 => "0000000000000000000001010100000100",
			5520 => "00000001001111000101011010001001",
			5521 => "00000000000000000101011010001001",
			5522 => "0000001000000000001000010100000100",
			5523 => "11111110001010000101011010001001",
			5524 => "0000001011000000000100010000000100",
			5525 => "00000001001101010101011010001001",
			5526 => "00000000000000000101011010001001",
			5527 => "0000001101000000001111010000000100",
			5528 => "11111110011010100101011010001001",
			5529 => "0000000110000000001011001100001000",
			5530 => "0000001001000000001000010000000100",
			5531 => "00000010000100110101011010001001",
			5532 => "11111111000011100101011010001001",
			5533 => "0000001101000000000011000000000100",
			5534 => "11111110100001100101011010001001",
			5535 => "0000001100000000001011011100000100",
			5536 => "00000001001011000101011010001001",
			5537 => "11111111100111010101011010001001",
			5538 => "0000000000000000001100000101100000",
			5539 => "0000001000000000001000100100100000",
			5540 => "0000001110000000000100001000000100",
			5541 => "11111111000000100101011101110101",
			5542 => "0000000001000000000110101000001100",
			5543 => "0000001011000000001101111000001000",
			5544 => "0000001100000000001000111000000100",
			5545 => "00000010101101110101011101110101",
			5546 => "00000000000000000101011101110101",
			5547 => "00000110011011110101011101110101",
			5548 => "0000001011000000000100001000000100",
			5549 => "11111110101101100101011101110101",
			5550 => "0000000001000000000000111100001000",
			5551 => "0000000110000000001101111100000100",
			5552 => "00000001101000000101011101110101",
			5553 => "00000000100110010101011101110101",
			5554 => "11111111001110100101011101110101",
			5555 => "0000000111000000001000011000100000",
			5556 => "0000000111000000000001101000010000",
			5557 => "0000001101000000000101110000001000",
			5558 => "0000000010000000001001100000000100",
			5559 => "11111110011000110101011101110101",
			5560 => "11111111111111000101011101110101",
			5561 => "0000000001000000000000111100000100",
			5562 => "00000001100001110101011101110101",
			5563 => "00000000000000000101011101110101",
			5564 => "0000000010000000000010000100001000",
			5565 => "0000000101000000000111100000000100",
			5566 => "00000000000011010101011101110101",
			5567 => "11111110100101110101011101110101",
			5568 => "0000000101000000001001010000000100",
			5569 => "11111100000111000101011101110101",
			5570 => "00000000000000000101011101110101",
			5571 => "0000000111000000001000011000010000",
			5572 => "0000001110000000001100010000001000",
			5573 => "0000001001000000001111000000000100",
			5574 => "00000001101000010101011101110101",
			5575 => "11111111001101110101011101110101",
			5576 => "0000001101000000001001011100000100",
			5577 => "00000111010111000101011101110101",
			5578 => "00000010011010010101011101110101",
			5579 => "0000000110000000000100110100000100",
			5580 => "00000001011111000101011101110101",
			5581 => "0000000100000000000000010000001000",
			5582 => "0000000101000000000101001000000100",
			5583 => "11111111111110100101011101110101",
			5584 => "11111110000110100101011101110101",
			5585 => "00000000110011000101011101110101",
			5586 => "0000000001000000001111001100000100",
			5587 => "11111110011000100101011101110101",
			5588 => "0000001001000000001101011000001000",
			5589 => "0000000110000000001011001100000100",
			5590 => "00000011101100100101011101110101",
			5591 => "11111111000110100101011101110101",
			5592 => "0000000101000000000000010000001000",
			5593 => "0000000110000000001010011000000100",
			5594 => "00000000111111010101011101110101",
			5595 => "11111110011010110101011101110101",
			5596 => "00000010100101110101011101110101",
			5597 => "0000000000000000001011010101001100",
			5598 => "0000001100000000000001101001001000",
			5599 => "0000001000000000000111110100011100",
			5600 => "0000001110000000001110101000010100",
			5601 => "0000000001000000000111100100001100",
			5602 => "0000001110000000001011000000001000",
			5603 => "0000001100000000000110000100000100",
			5604 => "11111111010111110101100000110001",
			5605 => "00000000010010100101100000110001",
			5606 => "00000001100010010101100000110001",
			5607 => "0000001100000000001100110000000100",
			5608 => "00000000000000000101100000110001",
			5609 => "11111110101110010101100000110001",
			5610 => "0000001001000000001001100100000100",
			5611 => "00000001011100100101100000110001",
			5612 => "00000000000000000101100000110001",
			5613 => "0000000011000000001100010000010100",
			5614 => "0000001100000000000100011000001100",
			5615 => "0000001101000000001110000100001000",
			5616 => "0000000111000000000110100100000100",
			5617 => "11111111010110110101100000110001",
			5618 => "00000000000000000101100000110001",
			5619 => "00000000000000000101100000110001",
			5620 => "0000001011000000000101100100000100",
			5621 => "00000000000000000101100000110001",
			5622 => "11111101101111000101100000110001",
			5623 => "0000001000000000001000100100001000",
			5624 => "0000001011000000000101100100000100",
			5625 => "00000000000000000101100000110001",
			5626 => "00000001011101010101100000110001",
			5627 => "0000000011000000001010000100001000",
			5628 => "0000001011000000000010001000000100",
			5629 => "00000000000000000101100000110001",
			5630 => "11111110100111110101100000110001",
			5631 => "0000000000000000000001010100000100",
			5632 => "00000001100001000101100000110001",
			5633 => "00000000000000000101100000110001",
			5634 => "00000011111100110101100000110001",
			5635 => "0000001011000000000101100100000100",
			5636 => "11111110011001100101100000110001",
			5637 => "0000001011000000001011011100001000",
			5638 => "0000001110000000000110111100000100",
			5639 => "00000001000110110101100000110001",
			5640 => "00000000000000000101100000110001",
			5641 => "0000000101000000001111100100000100",
			5642 => "11111110101010100101100000110001",
			5643 => "00000000000000000101100000110001",
			5644 => "0000000000000000001001101001011000",
			5645 => "0000001110000000001110101000100000",
			5646 => "0000000010000000000000110100011100",
			5647 => "0000000111000000001100101000011000",
			5648 => "0000001110000000000001101000010000",
			5649 => "0000001100000000000110000100001000",
			5650 => "0000001100000000000100000000000100",
			5651 => "00000000000000000101100100100101",
			5652 => "11111110101011010101100100100101",
			5653 => "0000000101000000000110100100000100",
			5654 => "00000010000010100101100100100101",
			5655 => "00000000000000000101100100100101",
			5656 => "0000001100000000000110000100000100",
			5657 => "00000001100111110101100100100101",
			5658 => "00000000000000000101100100100101",
			5659 => "11111110110100010101100100100101",
			5660 => "11111110011101010101100100100101",
			5661 => "0000001100000000001000000000011000",
			5662 => "0000001001000000000100111100010100",
			5663 => "0000000111000000001111011100010000",
			5664 => "0000000111000000001000011000001000",
			5665 => "0000001001000000001111000000000100",
			5666 => "00000001100101110101100100100101",
			5667 => "00000000000000100101100100100101",
			5668 => "0000000010000000000110010000000100",
			5669 => "00000000000000000101100100100101",
			5670 => "00000010010110100101100100100101",
			5671 => "11111111111010010101100100100101",
			5672 => "11111110111010110101100100100101",
			5673 => "0000001101000000001010001000010100",
			5674 => "0000000000000000000101000100001000",
			5675 => "0000000011000000001100000000000100",
			5676 => "00000000000000000101100100100101",
			5677 => "00000001010100100101100100100101",
			5678 => "0000000010000000001111010100001000",
			5679 => "0000001011000000001011011100000100",
			5680 => "00000000000000000101100100100101",
			5681 => "11111101001010010101100100100101",
			5682 => "00000000000000000101100100100101",
			5683 => "0000001011000000000100010000000100",
			5684 => "00000001111000000101100100100101",
			5685 => "0000001110000000000111010100000100",
			5686 => "11111111011011110101100100100101",
			5687 => "00000000110001100101100100100101",
			5688 => "0000000010000000000010110000010100",
			5689 => "0000001000000000000110011100010000",
			5690 => "0000001101000000001111010000000100",
			5691 => "11111110101011010101100100100101",
			5692 => "0000001011000000001011011100001000",
			5693 => "0000001110000000000110111100000100",
			5694 => "00000001100001110101100100100101",
			5695 => "00000000000000000101100100100101",
			5696 => "11111110111111100101100100100101",
			5697 => "11111110011010000101100100100101",
			5698 => "0000001010000000000001010000001100",
			5699 => "0000000101000000000010000000000100",
			5700 => "00000101011100010101100100100101",
			5701 => "0000000011000000001101001000000100",
			5702 => "00000000000000000101100100100101",
			5703 => "00000001110110110101100100100101",
			5704 => "11111110100100110101100100100101",
			5705 => "0000001000000000001001000101100000",
			5706 => "0000001000000000001000100100100000",
			5707 => "0000001110000000000100001000000100",
			5708 => "11111111000101010101101000011001",
			5709 => "0000000001000000000110101000000100",
			5710 => "00000010111101000101101000011001",
			5711 => "0000001111000000000010001000001100",
			5712 => "0000000001000000000111100100001000",
			5713 => "0000000111000000000110000100000100",
			5714 => "11111111101010100101101000011001",
			5715 => "00000001100100000101101000011001",
			5716 => "11111110101001110101101000011001",
			5717 => "0000001001000000001111000000000100",
			5718 => "00000001100111110101101000011001",
			5719 => "0000000110000000001101111100000100",
			5720 => "00000001010000100101101000011001",
			5721 => "11111111100000110101101000011001",
			5722 => "0000000111000000001000011000100000",
			5723 => "0000000111000000000001101000010000",
			5724 => "0000001101000000000101110000001000",
			5725 => "0000000010000000001001100000000100",
			5726 => "11111110010111110101101000011001",
			5727 => "00000000000000000101101000011001",
			5728 => "0000001001000000000100111100000100",
			5729 => "00000001100010010101101000011001",
			5730 => "00000000000000000101101000011001",
			5731 => "0000000010000000000010000100001000",
			5732 => "0000000101000000000111100000000100",
			5733 => "00000000000101000101101000011001",
			5734 => "11111110101101000101101000011001",
			5735 => "0000001111000000000110111100000100",
			5736 => "11111100100011100101101000011001",
			5737 => "00000000000000000101101000011001",
			5738 => "0000000111000000001000011000010000",
			5739 => "0000000011000000001010000100001000",
			5740 => "0000001001000000001111000000000100",
			5741 => "00000001001100000101101000011001",
			5742 => "11111111001101000101101000011001",
			5743 => "0000000001000000000000111100000100",
			5744 => "00000010110111010101101000011001",
			5745 => "00000000000000000101101000011001",
			5746 => "0000000110000000000100110100000100",
			5747 => "00000001010101010101101000011001",
			5748 => "0000001101000000000011001000001000",
			5749 => "0000000101000000000101001000000100",
			5750 => "00000000000000000101101000011001",
			5751 => "11111110001011110101101000011001",
			5752 => "00000000101110000101101000011001",
			5753 => "0000000001000000001111001100000100",
			5754 => "11111110011000100101101000011001",
			5755 => "0000001001000000001101011000001000",
			5756 => "0000001000000000001001101000000100",
			5757 => "00000010110111110101101000011001",
			5758 => "11111111100000100101101000011001",
			5759 => "0000000101000000000000010000001100",
			5760 => "0000001000000000000001010000001000",
			5761 => "0000001001000000000101010000000100",
			5762 => "00000000100111000101101000011001",
			5763 => "11111111001010100101101000011001",
			5764 => "11111110011011000101101000011001",
			5765 => "00000010001011110101101000011001",
			5766 => "0000000111000000001101100000000100",
			5767 => "11111110011111010101101011011101",
			5768 => "0000000111000000001000011000111100",
			5769 => "0000001000000000000111110100011000",
			5770 => "0000000010000000001101000100010000",
			5771 => "0000000110000000001101011100000100",
			5772 => "00000001010011010101101011011101",
			5773 => "0000001100000000001100110000001000",
			5774 => "0000001111000000001010011100000100",
			5775 => "11111111100000100101101011011101",
			5776 => "00000000101100110101101011011101",
			5777 => "11111111001000010101101011011101",
			5778 => "0000001001000000001001100100000100",
			5779 => "00000001010000100101101011011101",
			5780 => "00000000000000000101101011011101",
			5781 => "0000001101000000000010011100010100",
			5782 => "0000000000000000000110011100000100",
			5783 => "00000000000000000101101011011101",
			5784 => "0000001111000000000111011000001000",
			5785 => "0000000111000000000001101000000100",
			5786 => "11111110101011100101101011011101",
			5787 => "00000000000000000101101011011101",
			5788 => "0000000101000000001100100100000100",
			5789 => "11111111111001000101101011011101",
			5790 => "00000000000000000101101011011101",
			5791 => "0000001010000000000000001000000100",
			5792 => "00000001001001010101101011011101",
			5793 => "0000000110000000001101111100000100",
			5794 => "11111110110111010101101011011101",
			5795 => "0000000110000000001100011000000100",
			5796 => "00000000100110110101101011011101",
			5797 => "00000000000000000101101011011101",
			5798 => "0000000111000000001111011100010000",
			5799 => "0000001001000000001000010000001100",
			5800 => "0000000010000000000110010000000100",
			5801 => "00000000000000000101101011011101",
			5802 => "0000001101000000000101110000000100",
			5803 => "00000000000000000101101011011101",
			5804 => "00000001011001000101101011011101",
			5805 => "11111111111101100101101011011101",
			5806 => "0000001110000000001011111000000100",
			5807 => "11111111001101010101101011011101",
			5808 => "0000001001000000001010100000001100",
			5809 => "0000001000000000001001101000001000",
			5810 => "0000000110000000000101010000000100",
			5811 => "00000000111110100101101011011101",
			5812 => "00000000000000000101101011011101",
			5813 => "00000000000000000101101011011101",
			5814 => "11111111101011100101101011011101",
			5815 => "0000000111000000001101100000000100",
			5816 => "11111110011110000101101110010011",
			5817 => "0000001010000000000001010001010100",
			5818 => "0000001101000000001010001000111100",
			5819 => "0000001010000000000000001000100000",
			5820 => "0000001100000000000100011000010000",
			5821 => "0000000010000000001101000100001000",
			5822 => "0000000111000000001100101000000100",
			5823 => "00000000100111000101101110010011",
			5824 => "11111111000000010101101110010011",
			5825 => "0000000001000000000000111100000100",
			5826 => "00000001011011010101101110010011",
			5827 => "00000000000000000101101110010011",
			5828 => "0000000101000000001100100100001000",
			5829 => "0000000110000000001101111100000100",
			5830 => "00000000010011110101101110010011",
			5831 => "11111110100111000101101110010011",
			5832 => "0000000010000000001110110100000100",
			5833 => "00000001001000100101101110010011",
			5834 => "11111111110010100101101110010011",
			5835 => "0000000011000000001010000100001100",
			5836 => "0000001111000000001111010100001000",
			5837 => "0000000110000000001101111100000100",
			5838 => "00000000000000000101101110010011",
			5839 => "11111110110111100101101110010011",
			5840 => "00000000000000000101101110010011",
			5841 => "0000000010000000000111011000001000",
			5842 => "0000000111000000001000011000000100",
			5843 => "00000000110110000101101110010011",
			5844 => "00000000000000000101101110010011",
			5845 => "0000000010000000000110101100000100",
			5846 => "11111110110101000101101110010011",
			5847 => "00000000000000000101101110010011",
			5848 => "0000000111000000001111011100001000",
			5849 => "0000000001000000000000111100000100",
			5850 => "00000001101111000101101110010011",
			5851 => "00000000000000000101101110010011",
			5852 => "0000000011000000001000101000000100",
			5853 => "11111111001000100101101110010011",
			5854 => "0000000001000000001101111100001000",
			5855 => "0000001101000000000110010000000100",
			5856 => "00000000000000000101101110010011",
			5857 => "00000001000011100101101110010011",
			5858 => "11111111111111000101101110010011",
			5859 => "11111110111000110101101110010011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1940, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(3878, initial_addr_3'length));
	end generate gen_rom_4;

	gen_rom_5: if SELECT_ROM = 5 generate
		bank <= (
			0 => "00000000000000000000000000000101",
			1 => "00000000000000000000000000001001",
			2 => "00000000000000000000000000001101",
			3 => "00000000000000000000000000010001",
			4 => "00000000000000000000000000010101",
			5 => "00000000000000000000000000011001",
			6 => "00000000000000000000000000011101",
			7 => "00000000000000000000000000100001",
			8 => "00000000000000000000000000100101",
			9 => "00000000000000000000000000101001",
			10 => "00000000000000000000000000101101",
			11 => "00000000000000000000000000110001",
			12 => "00000000000000000000000000110101",
			13 => "00000000000000000000000000111001",
			14 => "00000000000000000000000000111101",
			15 => "00000000000000000000000001000001",
			16 => "00000000000000000000000001000101",
			17 => "00000000000000000000000001001001",
			18 => "00000000000000000000000001001101",
			19 => "00000000000000000000000001010001",
			20 => "00000000000000000000000001010101",
			21 => "00000000000000000000000001011001",
			22 => "00000000000000000000000001011101",
			23 => "00000000000000000000000001100001",
			24 => "00000000000000000000000001100101",
			25 => "00000000000000000000000001101001",
			26 => "00000000000000000000000001101101",
			27 => "00000000000000000000000001110001",
			28 => "00000000000000000000000001110101",
			29 => "00000000000000000000000001111001",
			30 => "00000000000000000000000001111101",
			31 => "00000000000000000000000010000001",
			32 => "00000000000000000000000010000101",
			33 => "0000000100000000001011001000000100",
			34 => "11111111010101010000000010010001",
			35 => "00000000000000000000000010010001",
			36 => "0000000100000000001011001000000100",
			37 => "11111111100011100000000010011101",
			38 => "00000000000000000000000010011101",
			39 => "0000000100000000001011001000000100",
			40 => "11111111110101010000000010101001",
			41 => "00000000000000000000000010101001",
			42 => "0000000111000000000111010000000100",
			43 => "11111111111101000000000010110101",
			44 => "00000000000000000000000010110101",
			45 => "0000000010000000001110000000000100",
			46 => "11111111110010110000000011000001",
			47 => "00000000000000000000000011000001",
			48 => "0000000100000000001011100100000100",
			49 => "11111111110000010000000011001101",
			50 => "00000000000000000000000011001101",
			51 => "0000001100000000000100011000000100",
			52 => "00000000000000000000000011011001",
			53 => "00000000000001010000000011011001",
			54 => "0000000100000000001011100100000100",
			55 => "11111111111010100000000011100101",
			56 => "00000000000000000000000011100101",
			57 => "0000000100000000000001100100000100",
			58 => "11111111111100000000000011110001",
			59 => "00000000000000000000000011110001",
			60 => "0000000100000000001011100100000100",
			61 => "11111111111001100000000011111101",
			62 => "00000000000000000000000011111101",
			63 => "0000001100000000000100011000000100",
			64 => "00000000000000000000000100001001",
			65 => "00000000000001000000000100001001",
			66 => "0000001100000000001001110100000100",
			67 => "11111111100011100000000100011101",
			68 => "0000000001000000001101011100000100",
			69 => "00000000010100010000000100011101",
			70 => "00000000000000000000000100011101",
			71 => "0000000111000000001111011100000100",
			72 => "11111111101011110000000100110001",
			73 => "0000000001000000001101011100000100",
			74 => "00000000001100000000000100110001",
			75 => "00000000000000000000000100110001",
			76 => "0000001100000000000100011000000100",
			77 => "00000000000000000000000101000101",
			78 => "0000001111000000000100101000000100",
			79 => "00000000000000000000000101000101",
			80 => "00000000000011000000000101000101",
			81 => "0000000111000000000111010000001000",
			82 => "0000000100000000001111101100000100",
			83 => "11111111001001000000000101100001",
			84 => "00000000000000000000000101100001",
			85 => "0000001001000000000100111100000100",
			86 => "00000000011101110000000101100001",
			87 => "00000000000000000000000101100001",
			88 => "0000000111000000001111011100001000",
			89 => "0000000100000000001010101000000100",
			90 => "11111111011010010000000101111101",
			91 => "00000000000000000000000101111101",
			92 => "0000000001000000000000111100000100",
			93 => "00000000011101000000000101111101",
			94 => "00000000000000000000000101111101",
			95 => "0000000010000000000101010100000100",
			96 => "11111110010110010000000110011001",
			97 => "0000001001000000001000010000001000",
			98 => "0000000110000000000101010000000100",
			99 => "00000011100000010000000110011001",
			100 => "00000010101000110000000110011001",
			101 => "11111110011011110000000110011001",
			102 => "0000001100000000000100011000000100",
			103 => "11111110111001100000000110110101",
			104 => "0000000001000000001111001100001000",
			105 => "0000001111000000000100101000000100",
			106 => "00000000000000000000000110110101",
			107 => "00000000100110110000000110110101",
			108 => "00000000000000000000000110110101",
			109 => "0000001100000000001001110100000100",
			110 => "11111111100001100000000111010001",
			111 => "0000000001000000001101011100001000",
			112 => "0000001000000000001101100000000100",
			113 => "00000000010110100000000111010001",
			114 => "00000000000000000000000111010001",
			115 => "00000000000000000000000111010001",
			116 => "0000001100000000000100011000000100",
			117 => "11111111110101000000000111101101",
			118 => "0000000010000000001111010100000100",
			119 => "00000000000000000000000111101101",
			120 => "0000000011000000000100000100000100",
			121 => "00000000000000000000000111101101",
			122 => "00000000000011000000000111101101",
			123 => "0000001100000000000100011000000100",
			124 => "11111111111101010000001000001001",
			125 => "0000000010000000001111010100000100",
			126 => "00000000000000000000001000001001",
			127 => "0000001111000000000100101000000100",
			128 => "00000000000000000000001000001001",
			129 => "00000000000111110000001000001001",
			130 => "0000001100000000000100011000000100",
			131 => "00000000000000000000001000100101",
			132 => "0000001111000000000100101000000100",
			133 => "00000000000000000000001000100101",
			134 => "0000000010000000001111010100000100",
			135 => "00000000000000000000001000100101",
			136 => "00000000000100110000001000100101",
			137 => "0000001100000000000100011000000100",
			138 => "00000000000000000000001001000001",
			139 => "0000000010000000001111010100000100",
			140 => "00000000000000000000001001000001",
			141 => "0000000011000000000100000100000100",
			142 => "00000000000000000000001001000001",
			143 => "00000000000110010000001001000001",
			144 => "0000000010000000000101010100001100",
			145 => "0000000100000000000000000100000100",
			146 => "11111110011010110000001001100101",
			147 => "0000000011000000000100000100000100",
			148 => "11111110011011010000001001100101",
			149 => "00000010101110010000001001100101",
			150 => "0000000001000000000000111100000100",
			151 => "00000001101001010000001001100101",
			152 => "11111110110100000000001001100101",
			153 => "0000000010000000000101010100001100",
			154 => "0000000111000000001111011100000100",
			155 => "11111110011001100000001010001001",
			156 => "0000001011000000000010001000000100",
			157 => "00000010001101100000001010001001",
			158 => "11111110011110000000001010001001",
			159 => "0000000001000000000000111100000100",
			160 => "00000001100111010000001010001001",
			161 => "11111111001000000000001010001001",
			162 => "0000000111000000001111011100001100",
			163 => "0000000010000000001110000000000100",
			164 => "11111110011100010000001010101101",
			165 => "0000000000000000001100001000000100",
			166 => "11111111111111100000001010101101",
			167 => "00000000000000000000001010101101",
			168 => "0000000001000000001111001100000100",
			169 => "00000001100000110000001010101101",
			170 => "11111111000100100000001010101101",
			171 => "0000001100000000001001110100001000",
			172 => "0000000100000000000100110000000100",
			173 => "11111110100000100000001011010001",
			174 => "00000000000000000000001011010001",
			175 => "0000000001000000001101011100001000",
			176 => "0000000000000000000101100100000100",
			177 => "00000001010001100000001011010001",
			178 => "00000000000000000000001011010001",
			179 => "11111111100011010000001011010001",
			180 => "0000001100000000001001110100001000",
			181 => "0000000100000000000100110000000100",
			182 => "11111110101101110000001011110101",
			183 => "00000000000000000000001011110101",
			184 => "0000000001000000000000111100001000",
			185 => "0000000111000000001000011000000100",
			186 => "00000000000000000000001011110101",
			187 => "00000000111000110000001011110101",
			188 => "00000000000000000000001011110101",
			189 => "0000001100000000000100011000000100",
			190 => "11111110100010010000001100011001",
			191 => "0000000001000000001111001100001000",
			192 => "0000000111000000001111011100000100",
			193 => "00000000000000000000001100011001",
			194 => "00000001001011000000001100011001",
			195 => "0000001100000000001011011100000100",
			196 => "11111111010101000000001100011001",
			197 => "00000000000000000000001100011001",
			198 => "0000001100000000000100011000000100",
			199 => "11111110101010000000001100111101",
			200 => "0000000001000000001111001100001000",
			201 => "0000001111000000000100101000000100",
			202 => "00000000000000000000001100111101",
			203 => "00000000111000110000001100111101",
			204 => "0000000000000000001101111000000100",
			205 => "11111111101001110000001100111101",
			206 => "00000000000000000000001100111101",
			207 => "0000000010000000000011110100010000",
			208 => "0000000010000000001110111000001000",
			209 => "0000000010000000000101010100000100",
			210 => "11010100011011100000001101101001",
			211 => "11010110010000110000001101101001",
			212 => "0000000001000000000111101000000100",
			213 => "11101010110110110000001101101001",
			214 => "11010100100001010000001101101001",
			215 => "0000000001000000001101111100000100",
			216 => "11101100000001000000001101101001",
			217 => "11010100101100000000001101101001",
			218 => "0000000100000000001011001000000100",
			219 => "11111110101110010000001110001101",
			220 => "0000001100000000000100011000000100",
			221 => "00000000000000000000001110001101",
			222 => "0000000001000000000000111100001000",
			223 => "0000000001000000000010001100000100",
			224 => "00000000000000000000001110001101",
			225 => "00000000100100000000001110001101",
			226 => "00000000000000000000001110001101",
			227 => "0000001100000000000100011000000100",
			228 => "11111110111011100000001110110001",
			229 => "0000000001000000001111001100001100",
			230 => "0000000110000000001010011000000100",
			231 => "00000000000000000000001110110001",
			232 => "0000000000000000000101110100000100",
			233 => "00000000100101010000001110110001",
			234 => "00000000000000000000001110110001",
			235 => "00000000000000000000001110110001",
			236 => "0000000100000000001011001000000100",
			237 => "11111111000110100000001111010101",
			238 => "0000001100000000000100011000000100",
			239 => "00000000000000000000001111010101",
			240 => "0000000001000000000000111100001000",
			241 => "0000000001000000000010001100000100",
			242 => "00000000000000000000001111010101",
			243 => "00000000010101010000001111010101",
			244 => "00000000000000000000001111010101",
			245 => "0000001100000000000100011000000100",
			246 => "11111111010001000000001111111001",
			247 => "0000000001000000000000111100001100",
			248 => "0000000010000000001111010100000100",
			249 => "00000000000000000000001111111001",
			250 => "0000000000000000000101110100000100",
			251 => "00000000101110010000001111111001",
			252 => "00000000000000000000001111111001",
			253 => "00000000000000000000001111111001",
			254 => "0000001100000000000100011000000100",
			255 => "00000000000000000000010000011101",
			256 => "0000000001000000000000111100001100",
			257 => "0000001111000000000100101000000100",
			258 => "00000000000000000000010000011101",
			259 => "0000000010000000001111010100000100",
			260 => "00000000000000000000010000011101",
			261 => "00000000011111100000010000011101",
			262 => "00000000000000000000010000011101",
			263 => "0000000010000000000101010100010000",
			264 => "0000001100000000000100011000000100",
			265 => "11111110010111110000010001001001",
			266 => "0000000100000000000000000100000100",
			267 => "11111110011010010000010001001001",
			268 => "0000000100000000000111001100000100",
			269 => "00000110110001110000010001001001",
			270 => "11111111000001000000010001001001",
			271 => "0000000001000000000000111100000100",
			272 => "00000001111010010000010001001001",
			273 => "11111110100011000000010001001001",
			274 => "0000000010000000000101010100010000",
			275 => "0000001100000000000100011000000100",
			276 => "11111110011001110000010001110101",
			277 => "0000000001000000001111001100001000",
			278 => "0000001111000000001011110100000100",
			279 => "00000000000000000000010001110101",
			280 => "00000010001010100000010001110101",
			281 => "11111110011100100000010001110101",
			282 => "0000000001000000001110010100000100",
			283 => "00000001100110110000010001110101",
			284 => "11111111001100000000010001110101",
			285 => "0000000010000000000101010100010000",
			286 => "0000000100000000001111101100000100",
			287 => "11111110011010000000010010100001",
			288 => "0000000000000000001010111100001000",
			289 => "0000001100000000000011011100000100",
			290 => "00000000000000000000010010100001",
			291 => "00000001011000100000010010100001",
			292 => "11111110100100100000010010100001",
			293 => "0000000001000000001110010100000100",
			294 => "00000001100101000000010010100001",
			295 => "11111111010110110000010010100001",
			296 => "0000000010000000000101010100010000",
			297 => "0000001010000000001010100100001100",
			298 => "0000000111000000000111010000000100",
			299 => "11111110110001010000010011001101",
			300 => "0000000100000000001000001100000100",
			301 => "00000000000000000000010011001101",
			302 => "00000001010010110000010011001101",
			303 => "11111110011010100000010011001101",
			304 => "0000000001000000000000111100000100",
			305 => "00000001100010100000010011001101",
			306 => "11111111101001100000010011001101",
			307 => "0000000100000000000000101100001000",
			308 => "0000001100000000000100000100000100",
			309 => "11111110011100000000010011111001",
			310 => "00000000000000000000010011111001",
			311 => "0000001100000000000100011000000100",
			312 => "11111110111011100000010011111001",
			313 => "0000000001000000001111001100001000",
			314 => "0000000001000000000010001100000100",
			315 => "00000000000000000000010011111001",
			316 => "00000001011111100000010011111001",
			317 => "00000000000000000000010011111001",
			318 => "0000001100000000001001110100010000",
			319 => "0000000010000000001000101000000100",
			320 => "11111110011010110000010100101101",
			321 => "0000000000000000000000001100000100",
			322 => "11111110111101100000010100101101",
			323 => "0000001010000000001001101000000100",
			324 => "00000001000001110000010100101101",
			325 => "00000000000000000000010100101101",
			326 => "0000000001000000000000111100001000",
			327 => "0000000000000000001011010100000100",
			328 => "00000000000000000000010100101101",
			329 => "00000001100100010000010100101101",
			330 => "11111110101100010000010100101101",
			331 => "0000000010000000001110111000010100",
			332 => "0000000010000000000101010100000100",
			333 => "11111110010011110000010101100001",
			334 => "0000001100000000001111011100000100",
			335 => "00000101111011010000010101100001",
			336 => "0000001100000000000100000100000100",
			337 => "11111110101010100000010101100001",
			338 => "0000001100000000000001011000000100",
			339 => "00000001011111010000010101100001",
			340 => "11111111000010010000010101100001",
			341 => "0000000001000000000111101000000100",
			342 => "00000110001110100000010101100001",
			343 => "11111110011010010000010101100001",
			344 => "0000001100000000000100011000000100",
			345 => "00000000000000000000010110001101",
			346 => "0000000110000000000010101100010000",
			347 => "0000000110000000001010011000000100",
			348 => "00000000000000000000010110001101",
			349 => "0000000011000000000100000100000100",
			350 => "00000000000000000000010110001101",
			351 => "0000000010000000001111010100000100",
			352 => "00000000000000000000010110001101",
			353 => "00000000001110110000010110001101",
			354 => "00000000000000000000010110001101",
			355 => "0000001100000000000100011000000100",
			356 => "11111110011110000000010111000001",
			357 => "0000000001000000001111001100010000",
			358 => "0000000110000000001010011000000100",
			359 => "00000000000000000000010111000001",
			360 => "0000000001000000000010001100000100",
			361 => "00000000000000000000010111000001",
			362 => "0000000001000000001111001100000100",
			363 => "00000001010010010000010111000001",
			364 => "00000000000000000000010111000001",
			365 => "0000001100000000001011011100000100",
			366 => "11111111000000010000010111000001",
			367 => "00000000000000000000010111000001",
			368 => "0000000010000000000101010100011000",
			369 => "0000001100000000000100011000000100",
			370 => "11111110011010000000010111111101",
			371 => "0000001110000000001001100000010000",
			372 => "0000000110000000001010011000000100",
			373 => "11111110111110000000010111111101",
			374 => "0000000110000000001011001100001000",
			375 => "0000000010000000001111010100000100",
			376 => "00000000000000000000010111111101",
			377 => "00000001110101000000010111111101",
			378 => "00000000000000000000010111111101",
			379 => "11111110011110010000010111111101",
			380 => "0000001001000000000100101100000100",
			381 => "00000001100110000000010111111101",
			382 => "11111111010100000000010111111101",
			383 => "0000000010000000000101010100011100",
			384 => "0000001100000000000100011000000100",
			385 => "11111110010111010000011001001011",
			386 => "0000001100000000000100011000000100",
			387 => "11111111010110100000011001001011",
			388 => "0000001100000000001001110100010000",
			389 => "0000001100000000001001110100000100",
			390 => "11111110011100100000011001001011",
			391 => "0000001100000000001001110100000100",
			392 => "00000000111110110000011001001011",
			393 => "0000001100000000001001110100000100",
			394 => "11111110101011110000011001001011",
			395 => "00000000000000000000011001001011",
			396 => "11111110010111110000011001001011",
			397 => "0000000001000000000000111100001000",
			398 => "0000001111000000001001001100000100",
			399 => "00000010111010110000011001001011",
			400 => "00000010000101010000011001001011",
			401 => "11111110011111010000011001001011",
			402 => "00000000000000000000011001001101",
			403 => "00000000000000000000011001010001",
			404 => "00000000000000000000011001010101",
			405 => "00000000000000000000011001011001",
			406 => "00000000000000000000011001011101",
			407 => "00000000000000000000011001100001",
			408 => "00000000000000000000011001100101",
			409 => "00000000000000000000011001101001",
			410 => "00000000000000000000011001101101",
			411 => "00000000000000000000011001110001",
			412 => "00000000000000000000011001110101",
			413 => "00000000000000000000011001111001",
			414 => "00000000000000000000011001111101",
			415 => "00000000000000000000011010000001",
			416 => "00000000000000000000011010000101",
			417 => "00000000000000000000011010001001",
			418 => "00000000000000000000011010001101",
			419 => "00000000000000000000011010010001",
			420 => "00000000000000000000011010010101",
			421 => "00000000000000000000011010011001",
			422 => "00000000000000000000011010011101",
			423 => "00000000000000000000011010100001",
			424 => "00000000000000000000011010100101",
			425 => "00000000000000000000011010101001",
			426 => "00000000000000000000011010101101",
			427 => "00000000000000000000011010110001",
			428 => "00000000000000000000011010110101",
			429 => "00000000000000000000011010111001",
			430 => "00000000000000000000011010111101",
			431 => "00000000000000000000011011000001",
			432 => "00000000000000000000011011000101",
			433 => "00000000000000000000011011001001",
			434 => "00000000000000000000011011001101",
			435 => "0000000100000000001011001000000100",
			436 => "11111111011110110000011011011001",
			437 => "00000000000000000000011011011001",
			438 => "0000000100000000001011001000000100",
			439 => "11111111110011000000011011100101",
			440 => "00000000000000000000011011100101",
			441 => "0000000111000000000111010000000100",
			442 => "11111111111011100000011011110001",
			443 => "00000000000000000000011011110001",
			444 => "0000000010000000001110000000000100",
			445 => "11111111110000100000011011111101",
			446 => "00000000000000000000011011111101",
			447 => "0000000111000000001111011100000100",
			448 => "00000000000000000000011100001001",
			449 => "00000000000000010000011100001001",
			450 => "0000000100000000001011100100000100",
			451 => "11111111110001110000011100010101",
			452 => "00000000000000000000011100010101",
			453 => "0000000111000000000011100000000100",
			454 => "00000000000000000000011100100001",
			455 => "00000000000000010000011100100001",
			456 => "0000000100000000001011100100000100",
			457 => "11111111111011010000011100101101",
			458 => "00000000000000000000011100101101",
			459 => "0000000100000000000001100100000100",
			460 => "11111111111100110000011100111001",
			461 => "00000000000000000000011100111001",
			462 => "0000000100000000001011100100000100",
			463 => "11111111111010110000011101000101",
			464 => "00000000000000000000011101000101",
			465 => "0000000010000000000101010100000100",
			466 => "11111110011001110000011101011001",
			467 => "0000000001000000000000111100000100",
			468 => "00000001110011100000011101011001",
			469 => "11111110100101100000011101011001",
			470 => "0000001100000000001001110100000100",
			471 => "11111111100101010000011101101101",
			472 => "0000000001000000001101011100000100",
			473 => "00000000010010000000011101101101",
			474 => "00000000000000000000011101101101",
			475 => "0000000111000000001111011100000100",
			476 => "11111111101101100000011110000001",
			477 => "0000000001000000001101011100000100",
			478 => "00000000001011010000011110000001",
			479 => "00000000000000000000011110000001",
			480 => "0000001100000000000100011000000100",
			481 => "00000000000000000000011110010101",
			482 => "0000000010000000001111010100000100",
			483 => "00000000000000000000011110010101",
			484 => "00000000000101000000011110010101",
			485 => "0000000111000000000111010000001000",
			486 => "0000000100000000001111101100000100",
			487 => "11111111001011110000011110110001",
			488 => "00000000000000000000011110110001",
			489 => "0000000001000000000000111100000100",
			490 => "00000000011011110000011110110001",
			491 => "00000000000000000000011110110001",
			492 => "0000000010000000000101010100000100",
			493 => "11111110010100110000011111001101",
			494 => "0000000001000000001110010100001000",
			495 => "0000001111000000001010110100000100",
			496 => "00000110100001100000011111001101",
			497 => "00000100011010100000011111001101",
			498 => "11111110011000000000011111001101",
			499 => "0000000010000000000101010100000100",
			500 => "11111110010111110000011111101001",
			501 => "0000000001000000000000111100001000",
			502 => "0000001111000000001001001100000100",
			503 => "00000011110101100000011111101001",
			504 => "00000010011001000000011111101001",
			505 => "11111110011100100000011111101001",
			506 => "0000001011000000001010001100000100",
			507 => "11111110111110000000100000000101",
			508 => "0000000001000000001111001100001000",
			509 => "0000000101000000000111100000000100",
			510 => "00000000000000000000100000000101",
			511 => "00000000100101100000100000000101",
			512 => "00000000000000000000100000000101",
			513 => "0000001100000000000100011000000100",
			514 => "11111111110010110000100000100001",
			515 => "0000000010000000001111010100000100",
			516 => "00000000000000000000100000100001",
			517 => "0000000011000000000100000100000100",
			518 => "00000000000000000000100000100001",
			519 => "00000000000011110000100000100001",
			520 => "0000000111000000000011100000000100",
			521 => "11111111111101010000100000111101",
			522 => "0000000010000000001111010100000100",
			523 => "00000000000000000000100000111101",
			524 => "0000000011000000000100000100000100",
			525 => "00000000000000000000100000111101",
			526 => "00000000000111010000100000111101",
			527 => "0000001100000000000100011000000100",
			528 => "00000000000000000000100001011001",
			529 => "0000000010000000001111010100000100",
			530 => "00000000000000000000100001011001",
			531 => "0000001101000000000010001000000100",
			532 => "00000000000000000000100001011001",
			533 => "00000000000110000000100001011001",
			534 => "0000001011000000001001110100000100",
			535 => "00000000000000000000100001110101",
			536 => "0000000010000000001111010100000100",
			537 => "00000000000000000000100001110101",
			538 => "0000001111000000000100101000000100",
			539 => "00000000000000000000100001110101",
			540 => "00000000000011010000100001110101",
			541 => "0000001011000000001001110100000100",
			542 => "00000000000000000000100010010001",
			543 => "0000000010000000001111010100000100",
			544 => "00000000000000000000100010010001",
			545 => "0000000011000000000100000100000100",
			546 => "00000000000000000000100010010001",
			547 => "00000000000011110000100010010001",
			548 => "0000000010000000000101010100001100",
			549 => "0000000111000000001111011100000100",
			550 => "11111110011001100000100010110101",
			551 => "0000001011000000000010001000000100",
			552 => "00000010111110100000100010110101",
			553 => "11111110011100100000100010110101",
			554 => "0000000001000000000000111100000100",
			555 => "00000001101000000000100010110101",
			556 => "11111111000000100000100010110101",
			557 => "0000000010000000000101010100001100",
			558 => "0000001010000000001010100100001000",
			559 => "0000001000000000000001010000000100",
			560 => "11111110101011110000100011011001",
			561 => "00000001100100110000100011011001",
			562 => "11111110011010010000100011011001",
			563 => "0000000001000000000000111100000100",
			564 => "00000001100100000000100011011001",
			565 => "11111111100011000000100011011001",
			566 => "0000001100000000001001110100001100",
			567 => "0000000010000000001110000000000100",
			568 => "11111110011100110000100011111101",
			569 => "0000000010000000001110000000000100",
			570 => "00000000000000000000100011111101",
			571 => "11111111110100100000100011111101",
			572 => "0000000001000000001101011100000100",
			573 => "00000001011010000000100011111101",
			574 => "11111111000101100000100011111101",
			575 => "0000001100000000001001110100001000",
			576 => "0000000100000000000100110000000100",
			577 => "11111110100001010000100100100001",
			578 => "00000000000000000000100100100001",
			579 => "0000000001000000001101011100001000",
			580 => "0000000000000000000101100100000100",
			581 => "00000001001111010000100100100001",
			582 => "00000000000000000000100100100001",
			583 => "11111111100110010000100100100001",
			584 => "0000000100000000001011100100001000",
			585 => "0000001111000000001101001000000100",
			586 => "11111110110001100000100101000101",
			587 => "00000000000000000000100101000101",
			588 => "0000001011000000001001110100000100",
			589 => "00000000000000000000100101000101",
			590 => "0000000001000000000010001100000100",
			591 => "00000000000000000000100101000101",
			592 => "00000000011101110000100101000101",
			593 => "0000001100000000000100011000000100",
			594 => "11111110100011000000100101101001",
			595 => "0000000001000000001111001100001000",
			596 => "0000000111000000001111011100000100",
			597 => "00000000000000000000100101101001",
			598 => "00000001001000000000100101101001",
			599 => "0000001100000000001011011100000100",
			600 => "11111111011000100000100101101001",
			601 => "00000000000000000000100101101001",
			602 => "0000001100000000000100011000000100",
			603 => "11111110101011010000100110001101",
			604 => "0000000001000000001111001100001000",
			605 => "0000001111000000000100101000000100",
			606 => "00000000000000000000100110001101",
			607 => "00000000110101100000100110001101",
			608 => "0000000000000000001101111000000100",
			609 => "11111111101100000000100110001101",
			610 => "00000000000000000000100110001101",
			611 => "0000000100000000001011001000000100",
			612 => "11111110011110000000100110110001",
			613 => "0000001100000000000100011000000100",
			614 => "11111111010011110000100110110001",
			615 => "0000000001000000000000111100001000",
			616 => "0000000001000000000010001100000100",
			617 => "00000000000000000000100110110001",
			618 => "00000001010010010000100110110001",
			619 => "00000000000000000000100110110001",
			620 => "0000000100000000001011001000000100",
			621 => "11111110110000000000100111010101",
			622 => "0000001011000000001001110100000100",
			623 => "00000000000000000000100111010101",
			624 => "0000000001000000000000111100001000",
			625 => "0000000001000000000010001100000100",
			626 => "00000000000000000000100111010101",
			627 => "00000000100001110000100111010101",
			628 => "00000000000000000000100111010101",
			629 => "0000000100000000001011001000000100",
			630 => "11111111000001100000100111111001",
			631 => "0000001100000000000100011000000100",
			632 => "00000000000000000000100111111001",
			633 => "0000001001000000001000010000001000",
			634 => "0000000011000000000100000100000100",
			635 => "00000000000000000000100111111001",
			636 => "00000000011000100000100111111001",
			637 => "00000000000000000000100111111001",
			638 => "0000000111000000000011100000000100",
			639 => "11111111001101000000101000011101",
			640 => "0000000001000000000000111100001100",
			641 => "0000000010000000001111010100000100",
			642 => "00000000000000000000101000011101",
			643 => "0000000001000000000010001100000100",
			644 => "00000000000000000000101000011101",
			645 => "00000000110011000000101000011101",
			646 => "00000000000000000000101000011101",
			647 => "0000001100000000000100011000000100",
			648 => "11111111100001100000101001000001",
			649 => "0000000001000000000000111100001100",
			650 => "0000000110000000001010011000000100",
			651 => "00000000000000000000101001000001",
			652 => "0000000000000000000101100100000100",
			653 => "00000000011100100000101001000001",
			654 => "00000000000000000000101001000001",
			655 => "00000000000000000000101001000001",
			656 => "0000001100000000000100011000000100",
			657 => "00000000000000000000101001100101",
			658 => "0000000001000000000000111100001100",
			659 => "0000001111000000000100101000000100",
			660 => "00000000000000000000101001100101",
			661 => "0000000110000000001010011000000100",
			662 => "00000000000000000000101001100101",
			663 => "00000000011100010000101001100101",
			664 => "00000000000000000000101001100101",
			665 => "0000000010000000000101010100010000",
			666 => "0000001100000000000100011000000100",
			667 => "11111110011001000000101010010001",
			668 => "0000000001000000001111001100001000",
			669 => "0000000011000000001100101100000100",
			670 => "11111111100011000000101010010001",
			671 => "00000011011001000000101010010001",
			672 => "11111110011010010000101010010001",
			673 => "0000000001000000000000111100000100",
			674 => "00000001101010000000101010010001",
			675 => "11111110110001000000101010010001",
			676 => "0000001111000000000010111000010000",
			677 => "0000001100000000000100011000000100",
			678 => "11111110011001110000101010111101",
			679 => "0000000001000000001111001100001000",
			680 => "0000000001000000000010001100000100",
			681 => "00000000000000000000101010111101",
			682 => "00000001111110100000101010111101",
			683 => "11111110011101000000101010111101",
			684 => "0000000001000000001011111100000100",
			685 => "00000001100110010000101010111101",
			686 => "11111111000001010000101010111101",
			687 => "0000000010000000000101010100010000",
			688 => "0000000000000000000000001100000100",
			689 => "11111110011010010000101011101001",
			690 => "0000001000000000000010011000001000",
			691 => "0000001100000000001010000000000100",
			692 => "00000000000000000000101011101001",
			693 => "00000001010000010000101011101001",
			694 => "11111110100110000000101011101001",
			695 => "0000000001000000001110010100000100",
			696 => "00000001100100100000101011101001",
			697 => "11111111011010000000101011101001",
			698 => "0000000100000000000000101100001000",
			699 => "0000000010000000000101010100000100",
			700 => "11111110011011010000101100010101",
			701 => "00000000000000000000101100010101",
			702 => "0000001100000000000100011000000100",
			703 => "11111110110100010000101100010101",
			704 => "0000000001000000001111001100001000",
			705 => "0000000001000000000010001100000100",
			706 => "00000000000000000000101100010101",
			707 => "00000001100001010000101100010101",
			708 => "00000000000000000000101100010101",
			709 => "0000000010000000000101010100010000",
			710 => "0000000100000000000000000100000100",
			711 => "11111110011110010000101101000001",
			712 => "0000001000000000000010011000001000",
			713 => "0000000010000000001100111000000100",
			714 => "00000000000000000000101101000001",
			715 => "00000000001101000000101101000001",
			716 => "00000000000000000000101101000001",
			717 => "0000001001000000001000010000000100",
			718 => "00000001001100110000101101000001",
			719 => "00000000000000000000101101000001",
			720 => "0000001100000000001001110100010000",
			721 => "0000000010000000001000101000000100",
			722 => "11111110011011000000101101110101",
			723 => "0000000000000000000000001100000100",
			724 => "11111111000000010000101101110101",
			725 => "0000001010000000001001101000000100",
			726 => "00000000111011010000101101110101",
			727 => "00000000000000000000101101110101",
			728 => "0000000001000000000000111100001000",
			729 => "0000000000000000001011010100000100",
			730 => "00000000000000000000101101110101",
			731 => "00000001100010100000101101110101",
			732 => "11111110101110110000101101110101",
			733 => "0000000100000000001011001000000100",
			734 => "11111110100100000000101110100001",
			735 => "0000001100000000000100011000000100",
			736 => "00000000000000000000101110100001",
			737 => "0000000001000000000000111100001100",
			738 => "0000000010000000001000101000000100",
			739 => "00000000000000000000101110100001",
			740 => "0000000100000000001111110100000100",
			741 => "00000000111110000000101110100001",
			742 => "00000000000000000000101110100001",
			743 => "00000000000000000000101110100001",
			744 => "0000001100000000000100011000000100",
			745 => "11111110011101000000101111010101",
			746 => "0000000001000000001111001100010000",
			747 => "0000000110000000001010011000000100",
			748 => "00000000000000000000101111010101",
			749 => "0000000001000000000010001100000100",
			750 => "00000000000000000000101111010101",
			751 => "0000000001000000001111001100000100",
			752 => "00000001011000110000101111010101",
			753 => "00000000000000000000101111010101",
			754 => "0000001100000000001011011100000100",
			755 => "11111110111001100000101111010101",
			756 => "00000000000000000000101111010101",
			757 => "0000000010000000000101010100011000",
			758 => "0000001100000000000100011000000100",
			759 => "11111110011001000000110000010001",
			760 => "0000000000000000000000001100001100",
			761 => "0000001110000000001001100000001000",
			762 => "0000001111000000000110111100000100",
			763 => "11111110100010010000110000010001",
			764 => "00000011001001110000110000010001",
			765 => "11111110011010000000110000010001",
			766 => "0000001111000000001011011100000100",
			767 => "00000000000000000000110000010001",
			768 => "00000010101011100000110000010001",
			769 => "0000000001000000000000111100000100",
			770 => "00000001101011000000110000010001",
			771 => "11111110110010110000110000010001",
			772 => "0000000010000000000101010100011100",
			773 => "0000001100000000000100011000000100",
			774 => "11111110011000110000110001010101",
			775 => "0000000000000000000000001100010000",
			776 => "0000001110000000001001100000001100",
			777 => "0000000011000000000110111100000100",
			778 => "11111110011111100000110001010101",
			779 => "0000001110000000000110010000000100",
			780 => "00000000000000000000110001010101",
			781 => "00000111000010110000110001010101",
			782 => "11111110011001100000110001010101",
			783 => "0000001111000000001011011100000100",
			784 => "11111111110101110000110001010101",
			785 => "00000100000010100000110001010101",
			786 => "0000000001000000000000111100000100",
			787 => "00000001101101100000110001010101",
			788 => "11111110101101100000110001010101",
			789 => "0000000010000000000101010100100000",
			790 => "0000001100000000000100011000000100",
			791 => "11111110011001000000110010100011",
			792 => "0000000000000000000000001100010100",
			793 => "0000001011000000001011011100010000",
			794 => "0000001011000000001011011100000100",
			795 => "11111110011110100000110010100011",
			796 => "0000001010000000001010100100001000",
			797 => "0000000100000000001110110100000100",
			798 => "00000000000000000000110010100011",
			799 => "00000110100100000000110010100011",
			800 => "11111111100010100000110010100011",
			801 => "11111110011010000000110010100011",
			802 => "0000001111000000001011011100000100",
			803 => "11111111111100100000110010100011",
			804 => "00000011001101110000110010100011",
			805 => "0000000001000000000000111100000100",
			806 => "00000001101100010000110010100011",
			807 => "11111110110000000000110010100011",
			808 => "00000000000000000000110010100101",
			809 => "00000000000000000000110010101001",
			810 => "00000000000000000000110010101101",
			811 => "00000000000000000000110010110001",
			812 => "00000000000000000000110010110101",
			813 => "00000000000000000000110010111001",
			814 => "00000000000000000000110010111101",
			815 => "00000000000000000000110011000001",
			816 => "00000000000000000000110011000101",
			817 => "00000000000000000000110011001001",
			818 => "00000000000000000000110011001101",
			819 => "00000000000000000000110011010001",
			820 => "00000000000000000000110011010101",
			821 => "00000000000000000000110011011001",
			822 => "00000000000000000000110011011101",
			823 => "00000000000000000000110011100001",
			824 => "00000000000000000000110011100101",
			825 => "00000000000000000000110011101001",
			826 => "00000000000000000000110011101101",
			827 => "00000000000000000000110011110001",
			828 => "00000000000000000000110011110101",
			829 => "00000000000000000000110011111001",
			830 => "00000000000000000000110011111101",
			831 => "00000000000000000000110100000001",
			832 => "00000000000000000000110100000101",
			833 => "00000000000000000000110100001001",
			834 => "00000000000000000000110100001101",
			835 => "00000000000000000000110100010001",
			836 => "00000000000000000000110100010101",
			837 => "00000000000000000000110100011001",
			838 => "00000000000000000000110100011101",
			839 => "00000000000000000000110100100001",
			840 => "0000000100000000001011001000000100",
			841 => "11111111010000100000110100101101",
			842 => "00000000000000000000110100101101",
			843 => "0000000100000000001011001000000100",
			844 => "11111111100001100000110100111001",
			845 => "00000000000000000000110100111001",
			846 => "0000000100000000001011001000000100",
			847 => "11111111110100000000110101000101",
			848 => "00000000000000000000110101000101",
			849 => "0000000111000000000111010000000100",
			850 => "11111111111100010000110101010001",
			851 => "00000000000000000000110101010001",
			852 => "0000000100000000001011001000000100",
			853 => "11111111110001110000110101011101",
			854 => "00000000000000000000110101011101",
			855 => "0000000111000000001111011100000100",
			856 => "00000000000000000000110101101001",
			857 => "00000000000000000000110101101001",
			858 => "0000000100000000001011100100000100",
			859 => "11111111110011010000110101110101",
			860 => "00000000000000000000110101110101",
			861 => "0000000100000000001011100100000100",
			862 => "11111111111001010000110110000001",
			863 => "00000000000000000000110110000001",
			864 => "0000000100000000000001100100000100",
			865 => "11111111111010110000110110001101",
			866 => "00000000000000000000110110001101",
			867 => "0000000100000000001011100100000100",
			868 => "11111111111000100000110110011001",
			869 => "00000000000000000000110110011001",
			870 => "0000001100000000000100011000000100",
			871 => "00000000000000000000110110100101",
			872 => "00000000000001010000110110100101",
			873 => "0000000010000000000101010100000100",
			874 => "11111110011010010000110110111001",
			875 => "0000001001000000001000010000000100",
			876 => "00000001110001000000110110111001",
			877 => "11111110100111010000110110111001",
			878 => "0000000111000000001111011100000100",
			879 => "11111111101001110000110111001101",
			880 => "0000000001000000001101011100000100",
			881 => "00000000001101000000110111001101",
			882 => "00000000000000000000110111001101",
			883 => "0000001100000000000100011000000100",
			884 => "00000000000000000000110111100001",
			885 => "0000001111000000000100101000000100",
			886 => "00000000000000000000110111100001",
			887 => "00000000000100000000110111100001",
			888 => "0000000010000000000101010100001000",
			889 => "0000000000000000000001111100000100",
			890 => "11111110100101110000110111111101",
			891 => "00000000000000000000110111111101",
			892 => "0000000001000000001110010100000100",
			893 => "00000000101111010000110111111101",
			894 => "00000000000000000000110111111101",
			895 => "0000000111000000000111010000001000",
			896 => "0000000100000000001111101100000100",
			897 => "11111111001110100000111000011001",
			898 => "00000000000000000000111000011001",
			899 => "0000000001000000000000111100000100",
			900 => "00000000011010000000111000011001",
			901 => "00000000000000000000111000011001",
			902 => "0000000010000000000101010100000100",
			903 => "11111110010101110000111000110101",
			904 => "0000000001000000000000111100001000",
			905 => "0000000110000000000101010000000100",
			906 => "00000100000110100000111000110101",
			907 => "00000010111111000000111000110101",
			908 => "11111110011010100000111000110101",
			909 => "0000001100000000000100011000000100",
			910 => "11111110101111110000111001010001",
			911 => "0000000001000000001111001100001000",
			912 => "0000000100000000001111110100000100",
			913 => "00000000110101010000111001010001",
			914 => "00000000000000000000111001010001",
			915 => "00000000000000000000111001010001",
			916 => "0000000000000000001001110000001100",
			917 => "0000001100000000000111010000001000",
			918 => "0000000010000000000011110100000100",
			919 => "11111111010011000000111001101101",
			920 => "00000000000000000000111001101101",
			921 => "00000000000000000000111001101101",
			922 => "00000000000000000000111001101101",
			923 => "0000001100000000000100011000000100",
			924 => "11111111110100000000111010001001",
			925 => "0000000010000000001111010100000100",
			926 => "00000000000000000000111010001001",
			927 => "0000000011000000000100000100000100",
			928 => "00000000000000000000111010001001",
			929 => "00000000000011010000111010001001",
			930 => "0000001100000000000100011000000100",
			931 => "11111111111100110000111010100101",
			932 => "0000000010000000001111010100000100",
			933 => "00000000000000000000111010100101",
			934 => "0000000011000000000100000100000100",
			935 => "00000000000000000000111010100101",
			936 => "00000000001000000000111010100101",
			937 => "0000001100000000000100011000000100",
			938 => "00000000000000000000111011000001",
			939 => "0000001111000000000100101000000100",
			940 => "00000000000000000000111011000001",
			941 => "0000000010000000001111010100000100",
			942 => "00000000000000000000111011000001",
			943 => "00000000000101100000111011000001",
			944 => "0000001100000000000100011000000100",
			945 => "00000000000000000000111011011101",
			946 => "0000001111000000000100101000000100",
			947 => "00000000000000000000111011011101",
			948 => "0000000010000000001111010100000100",
			949 => "00000000000000000000111011011101",
			950 => "00000000000100010000111011011101",
			951 => "0000000010000000000101010100001100",
			952 => "0000001100000000000100011000000100",
			953 => "11111110011000100000111100000001",
			954 => "0000001100000000000100011000000100",
			955 => "00000000000000000000111100000001",
			956 => "11111110100000100000111100000001",
			957 => "0000000001000000000000111100000100",
			958 => "00000001101111000000111100000001",
			959 => "11111110101001000000111100000001",
			960 => "0000000010000000000101010100001100",
			961 => "0000000111000000001111011100000100",
			962 => "11111110011001100000111100100101",
			963 => "0000001011000000000010001000000100",
			964 => "00000010100010100000111100100101",
			965 => "11111110011101010000111100100101",
			966 => "0000000001000000000000111100000100",
			967 => "00000001100111100000111100100101",
			968 => "11111111000100010000111100100101",
			969 => "0000001100000000001001110100001100",
			970 => "0000000010000000001110000000000100",
			971 => "11111110011100000000111101001001",
			972 => "0000000010000000001110000000000100",
			973 => "00000000000000000000111101001001",
			974 => "11111111110010010000111101001001",
			975 => "0000000001000000001101011100000100",
			976 => "00000001011110110000111101001001",
			977 => "11111110111110100000111101001001",
			978 => "0000001100000000001001110100001000",
			979 => "0000000100000000000100110000000100",
			980 => "11111110011111110000111101101101",
			981 => "00000000000000000000111101101101",
			982 => "0000000001000000001101011100001000",
			983 => "0000000000000000000101100100000100",
			984 => "00000001010100100000111101101101",
			985 => "00000000000000000000111101101101",
			986 => "11111111011111000000111101101101",
			987 => "0000000111000000001111011100001000",
			988 => "0000000100000000001111101100000100",
			989 => "11111110100011010000111110010001",
			990 => "00000000000000000000111110010001",
			991 => "0000000001000000000000111100001000",
			992 => "0000000000000000001011010100000100",
			993 => "00000000000000000000111110010001",
			994 => "00000001000101100000111110010001",
			995 => "11111111111011000000111110010001",
			996 => "0000000111000000001111011100001000",
			997 => "0000000100000000001111101100000100",
			998 => "11111110111011000000111110110101",
			999 => "00000000000000000000111110110101",
			1000 => "0000001001000000000100111100001000",
			1001 => "0000000000000000001011010100000100",
			1002 => "00000000000000000000111110110101",
			1003 => "00000000101010010000111110110101",
			1004 => "00000000000000000000111110110101",
			1005 => "0000001100000000000100011000000100",
			1006 => "11111110101000100000111111011001",
			1007 => "0000000001000000001111001100001000",
			1008 => "0000001111000000000100101000000100",
			1009 => "00000000000000000000111111011001",
			1010 => "00000000111100110000111111011001",
			1011 => "0000000010000000000001001100000100",
			1012 => "11111111100110110000111111011001",
			1013 => "00000000000000000000111111011001",
			1014 => "0000001100000000000100011000000100",
			1015 => "11111110101100100000111111111101",
			1016 => "0000001001000000001010011000001000",
			1017 => "0000000100000000001111110100000100",
			1018 => "00000000111001100000111111111101",
			1019 => "00000000000000000000111111111101",
			1020 => "0000001001000000000100111100000100",
			1021 => "00000000000000000000111111111101",
			1022 => "11111111111110100000111111111101",
			1023 => "0000000100000000001011001000000100",
			1024 => "11111110011111000001000000100001",
			1025 => "0000001100000000000100011000000100",
			1026 => "11111111011011010001000000100001",
			1027 => "0000000001000000000000111100001000",
			1028 => "0000000001000000000010001100000100",
			1029 => "00000000000000000001000000100001",
			1030 => "00000001001101010001000000100001",
			1031 => "00000000000000000001000000100001",
			1032 => "0000001100000000000100011000000100",
			1033 => "11111110110111010001000001000101",
			1034 => "0000000001000000001111001100001100",
			1035 => "0000000110000000001010011000000100",
			1036 => "00000000000000000001000001000101",
			1037 => "0000000000000000000101110100000100",
			1038 => "00000000101011000001000001000101",
			1039 => "00000000000000000001000001000101",
			1040 => "00000000000000000001000001000101",
			1041 => "0000000100000000001011001000000100",
			1042 => "11111111000100000001000001101001",
			1043 => "0000000111000000000011100000000100",
			1044 => "00000000000000000001000001101001",
			1045 => "0000000001000000000000111100001000",
			1046 => "0000000001000000000010001100000100",
			1047 => "00000000000000000001000001101001",
			1048 => "00000000010110110001000001101001",
			1049 => "00000000000000000001000001101001",
			1050 => "0000001100000000000100011000000100",
			1051 => "11111111001110100001000010001101",
			1052 => "0000000001000000000000111100001100",
			1053 => "0000000010000000001111010100000100",
			1054 => "00000000000000000001000010001101",
			1055 => "0000000000000000000101110100000100",
			1056 => "00000000110000110001000010001101",
			1057 => "00000000000000000001000010001101",
			1058 => "00000000000000000001000010001101",
			1059 => "0000001100000000000100011000000100",
			1060 => "11111111100101110001000010110001",
			1061 => "0000000001000000000000111100001100",
			1062 => "0000000000000000001011010100000100",
			1063 => "00000000000000000001000010110001",
			1064 => "0000000001000000000010001100000100",
			1065 => "00000000000000000001000010110001",
			1066 => "00000000011010010001000010110001",
			1067 => "00000000000000000001000010110001",
			1068 => "0000000010000000000101010100010000",
			1069 => "0000001100000000000100011000000100",
			1070 => "11111110010111100001000011011101",
			1071 => "0000000000000000000110000100000100",
			1072 => "11111110011001110001000011011101",
			1073 => "0000001000000000001001110000000100",
			1074 => "00001101101010010001000011011101",
			1075 => "11111111000101000001000011011101",
			1076 => "0000000001000000000000111100000100",
			1077 => "00000001111111010001000011011101",
			1078 => "11111110100001100001000011011101",
			1079 => "0000000010000000000101010100010000",
			1080 => "0000001100000000000100011000000100",
			1081 => "11111110011001010001000100001001",
			1082 => "0000000001000000001111001100001000",
			1083 => "0000000110000000001010011000000100",
			1084 => "11111111110101000001000100001001",
			1085 => "00000010101010010001000100001001",
			1086 => "11111110011010110001000100001001",
			1087 => "0000000001000000000000111100000100",
			1088 => "00000001101000100001000100001001",
			1089 => "11111110110111010001000100001001",
			1090 => "0000000010000000000101010100010000",
			1091 => "0000000100000000001111101100000100",
			1092 => "11111110011010000001000100110101",
			1093 => "0000001000000000000010111100001000",
			1094 => "0000000010000000000110100000000100",
			1095 => "00000000000000000001000100110101",
			1096 => "00000001011110010001000100110101",
			1097 => "11111110100010110001000100110101",
			1098 => "0000000001000000001110010100000100",
			1099 => "00000001100101100001000100110101",
			1100 => "11111111010011110001000100110101",
			1101 => "0000000010000000000101010100010000",
			1102 => "0000001010000000001010100100001100",
			1103 => "0000000111000000000111010000000100",
			1104 => "11111110101110100001000101100001",
			1105 => "0000000100000000001000001100000100",
			1106 => "00000000000000000001000101100001",
			1107 => "00000001011110000001000101100001",
			1108 => "11111110011010100001000101100001",
			1109 => "0000000001000000000000111100000100",
			1110 => "00000001100011010001000101100001",
			1111 => "11111111100110100001000101100001",
			1112 => "0000000010000000000101010100010000",
			1113 => "0000001000000000001000110000000100",
			1114 => "11111110011011100001000110001101",
			1115 => "0000001100000000000100011000000100",
			1116 => "11111110110111010001000110001101",
			1117 => "0000000010000000000001011100000100",
			1118 => "00000000000000000001000110001101",
			1119 => "00000001001000000001000110001101",
			1120 => "0000000001000000000000111100000100",
			1121 => "00000001011101110001000110001101",
			1122 => "11111111110000100001000110001101",
			1123 => "0000000111000000001111011100001000",
			1124 => "0000000100000000001111101100000100",
			1125 => "11111110111101100001000110111001",
			1126 => "00000000000000000001000110111001",
			1127 => "0000001100000000001001110100000100",
			1128 => "00000000000000000001000110111001",
			1129 => "0000000110000000000010101100001000",
			1130 => "0000000000000000001011010100000100",
			1131 => "00000000000000000001000110111001",
			1132 => "00000000010000100001000110111001",
			1133 => "00000000000000000001000110111001",
			1134 => "0000001100000000001001110100010000",
			1135 => "0000000010000000001000101000000100",
			1136 => "11111110011011000001000111101101",
			1137 => "0000000100000000000100110000000100",
			1138 => "11111111000010110001000111101101",
			1139 => "0000001010000000001011010100000100",
			1140 => "00000000110101100001000111101101",
			1141 => "00000000000000000001000111101101",
			1142 => "0000000001000000001101011100000100",
			1143 => "00000001100001100001000111101101",
			1144 => "0000000001000000000000111100000100",
			1145 => "00000000000000000001000111101101",
			1146 => "11111110110001110001000111101101",
			1147 => "0000000100000000001011001000000100",
			1148 => "11111110100101000001001000011001",
			1149 => "0000001100000000000100011000000100",
			1150 => "00000000000000000001001000011001",
			1151 => "0000000001000000000000111100001100",
			1152 => "0000000010000000001000101000000100",
			1153 => "00000000000000000001001000011001",
			1154 => "0000000100000000001111110100000100",
			1155 => "00000000111010000001001000011001",
			1156 => "00000000000000000001001000011001",
			1157 => "00000000000000000001001000011001",
			1158 => "0000001100000000000100011000000100",
			1159 => "11111110011101100001001001001101",
			1160 => "0000000001000000001111001100010000",
			1161 => "0000000110000000001010011000000100",
			1162 => "00000000000000000001001001001101",
			1163 => "0000000001000000000010001100000100",
			1164 => "00000000000000000001001001001101",
			1165 => "0000000001000000001111001100000100",
			1166 => "00000001010101110001001001001101",
			1167 => "00000000000000000001001001001101",
			1168 => "0000001100000000001011011100000100",
			1169 => "11111110111101000001001001001101",
			1170 => "00000000000000000001001001001101",
			1171 => "0000001111000000000010111000011000",
			1172 => "0000000100000000001011100100000100",
			1173 => "11111110011000110001001010001001",
			1174 => "0000001111000000000100101000000100",
			1175 => "11111110011001000001001010001001",
			1176 => "0000000110000000001001100100000100",
			1177 => "00000101111111110001001010001001",
			1178 => "0000000001000000000111100100000100",
			1179 => "00000001110101110001001010001001",
			1180 => "0000000000000000000011011100000100",
			1181 => "00000000000000000001001010001001",
			1182 => "11111111011101010001001010001001",
			1183 => "0000000001000000000000111100000100",
			1184 => "00000001110110010001001010001001",
			1185 => "11111110011111010001001010001001",
			1186 => "0000000010000000000101010100011100",
			1187 => "0000001100000000000100011000000100",
			1188 => "11111110010111000001001011010101",
			1189 => "0000001100000000000100011000000100",
			1190 => "11111111010000000001001011010101",
			1191 => "0000001100000000001001110100010000",
			1192 => "0000001100000000001001110100000100",
			1193 => "11111110011011100001001011010101",
			1194 => "0000001100000000001001110100000100",
			1195 => "00000001000100010001001011010101",
			1196 => "0000001100000000001001110100000100",
			1197 => "11111110101001000001001011010101",
			1198 => "00000000000000000001001011010101",
			1199 => "11111110010111100001001011010101",
			1200 => "0000001001000000001000010000001000",
			1201 => "0000001111000000001001001100000100",
			1202 => "00000011010100010001001011010101",
			1203 => "00000010001101110001001011010101",
			1204 => "11111110011101110001001011010101",
			1205 => "0000000011000000000010111000101000",
			1206 => "0000000011000000000011110000100000",
			1207 => "0000000110000000001000010000010100",
			1208 => "0000001101000000001010000100010000",
			1209 => "0000000011000000000101000000000100",
			1210 => "11111110010101010001001100110011",
			1211 => "0000000011000000001100001100001000",
			1212 => "0000000011000000001100001100000100",
			1213 => "11111111001011000001001100110011",
			1214 => "11111111110001100001001100110011",
			1215 => "11111110010110100001001100110011",
			1216 => "00000000011011110001001100110011",
			1217 => "0000000001000000001111001100001000",
			1218 => "0000000011000000001101101100000100",
			1219 => "11111110101011000001001100110011",
			1220 => "00000011111010010001001100110011",
			1221 => "11111110010101010001001100110011",
			1222 => "0000000000000000000111111000000100",
			1223 => "11111110010111010001001100110011",
			1224 => "00000011100011000001001100110011",
			1225 => "0000000001000000001110010100000100",
			1226 => "00000011100001010001001100110011",
			1227 => "11111110010111110001001100110011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(402, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(808, initial_addr_3'length));
	end generate gen_rom_5;

	gen_rom_6: if SELECT_ROM = 6 generate
		bank <= (
			0 => "00000000000000000000000000000101",
			1 => "00000000000000000000000000001001",
			2 => "00000000000000000000000000001101",
			3 => "00000000000000000000000000010001",
			4 => "00000000000000000000000000010101",
			5 => "00000000000000000000000000011001",
			6 => "00000000000000000000000000011101",
			7 => "00000000000000000000000000100001",
			8 => "00000000000000000000000000100101",
			9 => "00000000000000000000000000101001",
			10 => "00000000000000000000000000101101",
			11 => "00000000000000000000000000110001",
			12 => "00000000000000000000000000110101",
			13 => "00000000000000000000000000111001",
			14 => "00000000000000000000000000111101",
			15 => "00000000000000000000000001000001",
			16 => "00000000000000000000000001000101",
			17 => "00000000000000000000000001001001",
			18 => "00000000000000000000000001001101",
			19 => "00000000000000000000000001010001",
			20 => "00000000000000000000000001010101",
			21 => "00000000000000000000000001011001",
			22 => "00000000000000000000000001011101",
			23 => "00000000000000000000000001100001",
			24 => "00000000000000000000000001100101",
			25 => "00000000000000000000000001101001",
			26 => "00000000000000000000000001101101",
			27 => "00000000000000000000000001110001",
			28 => "00000000000000000000000001110101",
			29 => "00000000000000000000000001111001",
			30 => "0000000010000000000111100000000100",
			31 => "00000000000000000000000010000101",
			32 => "11111111111110010000000010000101",
			33 => "0000000011000000001010101100000100",
			34 => "00000000000000000000000010010001",
			35 => "11111111110100100000000010010001",
			36 => "0000000010000000001100100100000100",
			37 => "00000000000000000000000010011101",
			38 => "11111111111010000000000010011101",
			39 => "0000000010000000001100100100000100",
			40 => "00000000000000000000000010101001",
			41 => "11111111111111000000000010101001",
			42 => "0000000110000000001101111100001000",
			43 => "0000000110000000001011111100000100",
			44 => "00000000000000000000000010111101",
			45 => "00000000001000010000000010111101",
			46 => "00000000000000000000000010111101",
			47 => "0000000110000000001101111100001000",
			48 => "0000000110000000001011111100000100",
			49 => "00000000000000000000000011010001",
			50 => "00000000000111100000000011010001",
			51 => "00000000000000000000000011010001",
			52 => "0000000100000000001011100100001000",
			53 => "0000001101000000001001110100000100",
			54 => "11111111101001000000000011100101",
			55 => "00000000000000000000000011100101",
			56 => "00000000000000000000000011100101",
			57 => "0000000110000000001101111100001000",
			58 => "0000000110000000001011111100000100",
			59 => "00000000000000000000000011111001",
			60 => "00000000000100110000000011111001",
			61 => "00000000000000000000000011111001",
			62 => "0000000110000000001101111100001000",
			63 => "0000000110000000001011111100000100",
			64 => "00000000000000000000000100001101",
			65 => "00000000000100000000000100001101",
			66 => "00000000000000000000000100001101",
			67 => "0000000010000000001100100100000100",
			68 => "00000000000000000000000100100001",
			69 => "0000000011000000000111000000000100",
			70 => "00000000000000000000000100100001",
			71 => "11111111111010000000000100100001",
			72 => "0000000110000000001101111100001000",
			73 => "0000000110000000001011111100000100",
			74 => "00000000000000000000000100110101",
			75 => "00000000000100000000000100110101",
			76 => "00000000000000000000000100110101",
			77 => "0000000110000000001101111100001000",
			78 => "0000000110000000001011111100000100",
			79 => "00000000000000000000000101001001",
			80 => "00000000000111110000000101001001",
			81 => "00000000000000000000000101001001",
			82 => "0000000110000000001101111100001000",
			83 => "0000000110000000001011111100000100",
			84 => "00000000000000000000000101011101",
			85 => "00000000000011010000000101011101",
			86 => "00000000000000000000000101011101",
			87 => "0000000110000000001101111100001000",
			88 => "0000000110000000001011111100000100",
			89 => "00000000000000000000000101110001",
			90 => "00000000000110110000000101110001",
			91 => "00000000000000000000000101110001",
			92 => "0000000110000000001101111100001000",
			93 => "0000000110000000001011111100000100",
			94 => "00000000000000000000000110001101",
			95 => "00000000000110000000000110001101",
			96 => "0000000010000000000111100000000100",
			97 => "00000000000000000000000110001101",
			98 => "11111111110000000000000110001101",
			99 => "0000000110000000001101111100001100",
			100 => "0000000010000000000111100000001000",
			101 => "0000000110000000001011111100000100",
			102 => "00000000000000000000000110101001",
			103 => "00000000001110100000000110101001",
			104 => "00000000000000000000000110101001",
			105 => "11111111110101000000000110101001",
			106 => "0000000010000000000111100000001100",
			107 => "0000000110000000001101111100001000",
			108 => "0000000110000000001011111100000100",
			109 => "00000000000000000000000111001101",
			110 => "00000000010001010000000111001101",
			111 => "00000000000000000000000111001101",
			112 => "0000000010000000001000001100000100",
			113 => "11111111100101000000000111001101",
			114 => "00000000000000000000000111001101",
			115 => "0000001101000000001001110100001000",
			116 => "0000000011000000000001110100000100",
			117 => "00000000000000000000000111110001",
			118 => "11111111110000110000000111110001",
			119 => "0000001110000000001100101100000100",
			120 => "00000000000000000000000111110001",
			121 => "0000001110000000000111011000000100",
			122 => "00000000001110110000000111110001",
			123 => "00000000000000000000000111110001",
			124 => "0000000100000000000011011000000100",
			125 => "11111111010110110000001000010101",
			126 => "0000001100000000000011011100001100",
			127 => "0000000110000000001101111100001000",
			128 => "0000000110000000000111101000000100",
			129 => "00000000000000000000001000010101",
			130 => "00000000011011100000001000010101",
			131 => "00000000000000000000001000010101",
			132 => "00000000000000000000001000010101",
			133 => "0000000110000000001101111100010000",
			134 => "0000000011000000000100011000000100",
			135 => "00000000000000000000001000111001",
			136 => "0000000110000000001011111100000100",
			137 => "00000000000000000000001000111001",
			138 => "0000001101000000001001110100000100",
			139 => "00000000000000000000001000111001",
			140 => "00000000011000000000001000111001",
			141 => "00000000000000000000001000111001",
			142 => "0000000110000000001101111100010000",
			143 => "0000000110000000001011111100000100",
			144 => "00000000000000000000001001100101",
			145 => "0000001000000000000100010100001000",
			146 => "0000001000000000001001000100000100",
			147 => "00000000000000000000001001100101",
			148 => "00000000001001110000001001100101",
			149 => "00000000000000000000001001100101",
			150 => "0000000011000000000111000100000100",
			151 => "00000000000000000000001001100101",
			152 => "11111111101110110000001001100101",
			153 => "0000000110000000001101111100010000",
			154 => "0000000011000000000100011000001000",
			155 => "0000000100000000000100111000000100",
			156 => "11111111111100100000001010011001",
			157 => "00000000000000000000001010011001",
			158 => "0000000100000000001111101000000100",
			159 => "00000000000000000000001010011001",
			160 => "00000000011111000000001010011001",
			161 => "0000000100000000001010010000001000",
			162 => "0000000101000000000001101000000100",
			163 => "11111111011010110000001010011001",
			164 => "00000000000000000000001010011001",
			165 => "00000000000000000000001010011001",
			166 => "0000001110000000000001010100010000",
			167 => "0000001000000000000100000000001100",
			168 => "0000001111000000000001111100001000",
			169 => "0000000100000000001110001000000100",
			170 => "00000010010100100000001011010101",
			171 => "00000011011111100000001011010101",
			172 => "11111110011001100000001011010101",
			173 => "11111110011000010000001011010101",
			174 => "0000001111000000000001111100001100",
			175 => "0000000111000000000000101000001000",
			176 => "0000000001000000001100100000000100",
			177 => "00000011100111110000001011010101",
			178 => "11111110100100100000001011010101",
			179 => "11111110010111000000001011010101",
			180 => "11111110010110100000001011010101",
			181 => "0000000010000000000111100000010100",
			182 => "0000000001000000001100110100010000",
			183 => "0000000110000000001101111100001100",
			184 => "0000000110000000001011111100000100",
			185 => "00000000000000000000001100001001",
			186 => "0000000000000000000001001000000100",
			187 => "00000000001010000000001100001001",
			188 => "00000000000000000000001100001001",
			189 => "00000000000000000000001100001001",
			190 => "00000000000000000000001100001001",
			191 => "0000000011000000000111000000000100",
			192 => "00000000000000000000001100001001",
			193 => "11111111101101000000001100001001",
			194 => "0000000100000000000011011000000100",
			195 => "11111110011111000000001100110101",
			196 => "0000000110000000001101111100010000",
			197 => "0000000111000000001110001100001100",
			198 => "0000000110000000001110010100000100",
			199 => "00000000000000000000001100110101",
			200 => "0000000010000000001110110100000100",
			201 => "00000001000101100000001100110101",
			202 => "00000000000000000000001100110101",
			203 => "11111111111101110000001100110101",
			204 => "11111111000100000000001100110101",
			205 => "0000000110000000001101111100010100",
			206 => "0000001101000000001010111100000100",
			207 => "00000000000000000000001101100001",
			208 => "0000000010000000001110101000000100",
			209 => "00000000000000000000001101100001",
			210 => "0000000011000000001100001000000100",
			211 => "00000000000000000000001101100001",
			212 => "0000001011000000000101100100000100",
			213 => "00000000011110100000001101100001",
			214 => "00000000000000000000001101100001",
			215 => "00000000000000000000001101100001",
			216 => "0000000001000000000000011000010100",
			217 => "0000000101000000001010111000010000",
			218 => "0000000110000000001101111100001100",
			219 => "0000000110000000000111101000000100",
			220 => "00000000000000000000001110100101",
			221 => "0000000010000000001100010100000100",
			222 => "00000001010001010000001110100101",
			223 => "00000000000000000000001110100101",
			224 => "00000000000000000000001110100101",
			225 => "11111111101111010000001110100101",
			226 => "0000001101000000001010011100000100",
			227 => "11111110100000010000001110100101",
			228 => "0000001100000000001000111000001000",
			229 => "0000001110000000000010001000000100",
			230 => "00000001001111010000001110100101",
			231 => "00000000000000000000001110100101",
			232 => "11111110111110000000001110100101",
			233 => "0000000100000000000011011000000100",
			234 => "11111110110111100000001111011001",
			235 => "0000001100000000000011011100010100",
			236 => "0000001011000000001100001000001100",
			237 => "0000001001000000000000011000001000",
			238 => "0000001111000000001010111000000100",
			239 => "00000000001110100000001111011001",
			240 => "00000000000000000000001111011001",
			241 => "11111111111001100000001111011001",
			242 => "0000000110000000001100011000000100",
			243 => "00000000110000110000001111011001",
			244 => "00000000000000000000001111011001",
			245 => "00000000000000000000001111011001",
			246 => "0000000100000000001011100100011000",
			247 => "0000001000000000000110011000001000",
			248 => "0000000010000000000111010100000100",
			249 => "11111110111000110000010000100101",
			250 => "00000001110110110000010000100101",
			251 => "0000000100000000001101110100000100",
			252 => "11111110011011100000010000100101",
			253 => "0000001101000000001001110100000100",
			254 => "11111110110100000000010000100101",
			255 => "0000001101000000000001011000000100",
			256 => "00000000111110000000010000100101",
			257 => "00000000000000000000010000100101",
			258 => "0000001011000000001001110000001100",
			259 => "0000000010000000000011001000001000",
			260 => "0000000110000000001110010100000100",
			261 => "00000000000000000000010000100101",
			262 => "00000001011110000000010000100101",
			263 => "00000000000000000000010000100101",
			264 => "11111110110010100000010000100101",
			265 => "0000001101000000001001110100011000",
			266 => "0000000100000000001011100100001000",
			267 => "0000001111000000000011011100000100",
			268 => "00000000000000000000010001110001",
			269 => "11111111000100110000010001110001",
			270 => "0000000010000000000011001000001100",
			271 => "0000001010000000000010101000001000",
			272 => "0000001010000000000101000100000100",
			273 => "00000000000000000000010001110001",
			274 => "00000000001101110000010001110001",
			275 => "00000000000000000000010001110001",
			276 => "00000000000000000000010001110001",
			277 => "0000001010000000000110011000001100",
			278 => "0000000100000000001111101000000100",
			279 => "00000000000000000000010001110001",
			280 => "0000000001000000001101101000000100",
			281 => "00000000101010110000010001110001",
			282 => "00000000000000000000010001110001",
			283 => "00000000000000000000010001110001",
			284 => "0000000110000000001101111100011100",
			285 => "0000001101000000001010111100010000",
			286 => "0000001111000000001010111000001100",
			287 => "0000000100000000000000101100000100",
			288 => "00000000000000000000010010101101",
			289 => "0000000110000000001110010100000100",
			290 => "00000000000000000000010010101101",
			291 => "00000000010101100000010010101101",
			292 => "11111111010001010000010010101101",
			293 => "0000001001000000001110100000000100",
			294 => "00000000000000000000010010101101",
			295 => "0000000100000000001111101000000100",
			296 => "00000000000000000000010010101101",
			297 => "00000001001110110000010010101101",
			298 => "11111111000101100000010010101101",
			299 => "0000000110000000001101111100011100",
			300 => "0000001101000000001010111100001100",
			301 => "0000001111000000001010111000001000",
			302 => "0000001010000000000110011100000100",
			303 => "00000000000000000000010011101001",
			304 => "00000000001011010000010011101001",
			305 => "11111111011111010000010011101001",
			306 => "0000000100000000001011110000000100",
			307 => "00000000000000000000010011101001",
			308 => "0000001001000000001110100000000100",
			309 => "00000000000000000000010011101001",
			310 => "0000000110000000000001111000000100",
			311 => "00000000000000000000010011101001",
			312 => "00000000101100000000010011101001",
			313 => "11111111010101000000010011101001",
			314 => "0000000110000000000001111000011100",
			315 => "0000000011000000000111000000001000",
			316 => "0000000110000000000111101000000100",
			317 => "00000000000000000000010100111101",
			318 => "00000000100001110000010100111101",
			319 => "0000000011000000000100011000001100",
			320 => "0000001111000000000101101100000100",
			321 => "00000000000000000000010100111101",
			322 => "0000000001000000001110011100000100",
			323 => "00000000000000000000010100111101",
			324 => "11111111010011000000010100111101",
			325 => "0000001010000000001010100100000100",
			326 => "00000000000000000000010100111101",
			327 => "00000000100110000000010100111101",
			328 => "0000000101000000000100000100001000",
			329 => "0000000011000000000111000100000100",
			330 => "00000000000000000000010100111101",
			331 => "11111110101101000000010100111101",
			332 => "0000001011000000000111001000000100",
			333 => "00000000000000000000010100111101",
			334 => "11111111101011000000010100111101",
			335 => "0000000100000000000011011000001100",
			336 => "0000001000000000000110011000001000",
			337 => "0000000000000000001001101000000100",
			338 => "11111111010000010000010110000001",
			339 => "00000001000101000000010110000001",
			340 => "11111110011110000000010110000001",
			341 => "0000000110000000001101111100010100",
			342 => "0000000111000000001110001100010000",
			343 => "0000000110000000000111101000000100",
			344 => "00000000000000000000010110000001",
			345 => "0000000001000000000000011000000100",
			346 => "00000001010111010000010110000001",
			347 => "0000000100000000000000100000000100",
			348 => "00000000110001100000010110000001",
			349 => "11111111011110110000010110000001",
			350 => "11111111110000000000010110000001",
			351 => "11111110111111100000010110000001",
			352 => "0000000100000000000011011000000100",
			353 => "11111111011011010000010110110101",
			354 => "0000001100000000000011011100010100",
			355 => "0000000110000000001101111100010000",
			356 => "0000000110000000001110010100000100",
			357 => "00000000000000000000010110110101",
			358 => "0000000010000000001100000000001000",
			359 => "0000001000000000000100010100000100",
			360 => "00000000011010010000010110110101",
			361 => "00000000000000000000010110110101",
			362 => "00000000000000000000010110110101",
			363 => "00000000000000000000010110110101",
			364 => "00000000000000000000010110110101",
			365 => "0000000110000000001101111100011100",
			366 => "0000000011000000000100011000010100",
			367 => "0000000001000000000000011000010000",
			368 => "0000000101000000000011100000001100",
			369 => "0000000110000000001110010100000100",
			370 => "00000000000000000000010111110001",
			371 => "0000000010000000000011001000000100",
			372 => "00000000111100100000010111110001",
			373 => "00000000000000000000010111110001",
			374 => "00000000000000000000010111110001",
			375 => "11111110110110110000010111110001",
			376 => "0000000100000000001111101000000100",
			377 => "00000000000000000000010111110001",
			378 => "00000001010010000000010111110001",
			379 => "11111110101000100000010111110001",
			380 => "0000001011000000000110000100010100",
			381 => "0000000100000000000101100000001000",
			382 => "0000000001000000001100100000000100",
			383 => "00000000000000000000011001000101",
			384 => "11111110100001110000011001000101",
			385 => "0000000010000000000011001000001000",
			386 => "0000001000000000001011000100000100",
			387 => "00000001000000010000011001000101",
			388 => "00000000000000000000011001000101",
			389 => "00000000000000000000011001000101",
			390 => "0000001100000000000100001000010100",
			391 => "0000001010000000000001010000010000",
			392 => "0000000100000000001111101000000100",
			393 => "00000000000000000000011001000101",
			394 => "0000000001000000001101101000001000",
			395 => "0000001100000000000100000000000100",
			396 => "00000000000000000000011001000101",
			397 => "00000001011110110000011001000101",
			398 => "00000000000000000000011001000101",
			399 => "11111111100110010000011001000101",
			400 => "11111111001100000000011001000101",
			401 => "0000000110000000001101111100100000",
			402 => "0000000011000000000100011000010100",
			403 => "0000001010000000000110011100000100",
			404 => "11111111010100100000011010001001",
			405 => "0000000001000000000000011000001100",
			406 => "0000000101000000000100011000001000",
			407 => "0000001111000000001010011100000100",
			408 => "00000000100101110000011010001001",
			409 => "00000000000000000000011010001001",
			410 => "00000000000000000000011010001001",
			411 => "00000000000000000000011010001001",
			412 => "0000000100000000001111101000000100",
			413 => "00000000000000000000011010001001",
			414 => "0000000101000000000111001000000100",
			415 => "00000000000000000000011010001001",
			416 => "00000000111111100000011010001001",
			417 => "11111111001011100000011010001001",
			418 => "0000000110000000001101111100100000",
			419 => "0000000011000000000100011000010100",
			420 => "0000000001000000000000011000010000",
			421 => "0000000101000000000100011000001100",
			422 => "0000000010000000000011001000001000",
			423 => "0000001010000000000110011100000100",
			424 => "00000000000000000000011011001101",
			425 => "00000000011010010000011011001101",
			426 => "00000000000000000000011011001101",
			427 => "00000000000000000000011011001101",
			428 => "11111111100010000000011011001101",
			429 => "0000000100000000001111101000000100",
			430 => "00000000000000000000011011001101",
			431 => "0000000101000000000111001000000100",
			432 => "00000000000000000000011011001101",
			433 => "00000000101001000000011011001101",
			434 => "11111111011101010000011011001101",
			435 => "0000001110000000000001010100011000",
			436 => "0000000110000000001101111100010000",
			437 => "0000000010000000000011001000001100",
			438 => "0000000110000000001110010100000100",
			439 => "00000000000000000000011100101001",
			440 => "0000001000000000001011000100000100",
			441 => "00000001100111010000011100101001",
			442 => "00000000000000000000011100101001",
			443 => "00000000000000000000011100101001",
			444 => "0000000110000000001101111100000100",
			445 => "00000000000000000000011100101001",
			446 => "11111111010000100000011100101001",
			447 => "0000000100000000000011011000000100",
			448 => "11111110011010000000011100101001",
			449 => "0000000110000000001101111100010000",
			450 => "0000001110000000001100001000001100",
			451 => "0000000010000000001100100100001000",
			452 => "0000000100000000001011100100000100",
			453 => "11111111010010000000011100101001",
			454 => "00000001000100100000011100101001",
			455 => "11111110110010010000011100101001",
			456 => "00000001111010010000011100101001",
			457 => "11111110100000110000011100101001",
			458 => "0000000001000000000000011000010100",
			459 => "0000000101000000001010111000010000",
			460 => "0000000110000000001101111100001100",
			461 => "0000000110000000001110010100000100",
			462 => "11111111110010000000011110000101",
			463 => "0000000010000000000011001000000100",
			464 => "00000001100111100000011110000101",
			465 => "00000000000000000000011110000101",
			466 => "11111111010111000000011110000101",
			467 => "11111110110010010000011110000101",
			468 => "0000001000000000000110011000001000",
			469 => "0000000100000000001000100000000100",
			470 => "11111110110001110000011110000101",
			471 => "00000010110100000000011110000101",
			472 => "0000000100000000000011011000000100",
			473 => "11111110011010110000011110000101",
			474 => "0000000100000000000001101100001100",
			475 => "0000001101000000001011011100000100",
			476 => "11111111111100100000011110000101",
			477 => "0000000101000000000001011000000100",
			478 => "00000000111110010000011110000101",
			479 => "00000000000000000000011110000101",
			480 => "11111110111110010000011110000101",
			481 => "0000000100000000000011011000001100",
			482 => "0000001000000000000110011000001000",
			483 => "0000000000000000001011010100000100",
			484 => "11111110111001110000011111010001",
			485 => "00000010000010000000011111010001",
			486 => "11111110011011010000011111010001",
			487 => "0000000110000000001101111100011000",
			488 => "0000000111000000001110001100010100",
			489 => "0000000110000000001110010100000100",
			490 => "00000000000000000000011111010001",
			491 => "0000000001000000000000011000001000",
			492 => "0000000010000000000011001000000100",
			493 => "00000001100101010000011111010001",
			494 => "00000000000000000000011111010001",
			495 => "0000000001000000000110000000000100",
			496 => "11111111101110110000011111010001",
			497 => "00000000111010010000011111010001",
			498 => "11111111010101110000011111010001",
			499 => "11111110101011110000011111010001",
			500 => "0000000011000000000111000000010000",
			501 => "0000000110000000001101111100001100",
			502 => "0000001111000000000001111100001000",
			503 => "0000001000000000000000101000000100",
			504 => "00000010011000100000100000110101",
			505 => "00000001000111100000100000110101",
			506 => "00000000000010010000100000110101",
			507 => "11111110011110000000100000110101",
			508 => "0000001111000000001101010100010000",
			509 => "0000000101000000001010111100001100",
			510 => "0000000001000000001100100000001000",
			511 => "0000000101000000000011011100000100",
			512 => "00000010010000110000100000110101",
			513 => "00000011101010100000100000110101",
			514 => "11111110100100110000100000110101",
			515 => "11111110011000010000100000110101",
			516 => "0000000100000000000011011000000100",
			517 => "11111110010110110000100000110101",
			518 => "0000000110000000001101111100001100",
			519 => "0000000110000000000001111000000100",
			520 => "11111110011001100000100000110101",
			521 => "0000000100000000001111011000000100",
			522 => "00001010000001010000100000110101",
			523 => "11111110011110000000100000110101",
			524 => "11111110010111010000100000110101",
			525 => "0000000100000000000011011000001100",
			526 => "0000001000000000000110011000001000",
			527 => "0000000100000000001111100100000100",
			528 => "11111111010100100000100010001001",
			529 => "00000001000000000000100010001001",
			530 => "11111110011110100000100010001001",
			531 => "0000000110000000001101111100011100",
			532 => "0000000111000000001110001100011000",
			533 => "0000000001000000000000011000001100",
			534 => "0000000110000000000111101000000100",
			535 => "00000000000000000000100010001001",
			536 => "0000000010000000000011001000000100",
			537 => "00000001011000100000100010001001",
			538 => "00000000000000000000100010001001",
			539 => "0000001000000000001111001000001000",
			540 => "0000000110000000000101011100000100",
			541 => "00000000000000000000100010001001",
			542 => "00000001001010010000100010001001",
			543 => "11111111001110110000100010001001",
			544 => "11111111110101000000100010001001",
			545 => "11111111000010110000100010001001",
			546 => "0000000011000000000111000000001100",
			547 => "0000000110000000001101111100001000",
			548 => "0000001111000000001010111000000100",
			549 => "00000001110010100000100011111101",
			550 => "11111111100110010000100011111101",
			551 => "11111110100110110000100011111101",
			552 => "0000001111000000001010111000010100",
			553 => "0000000101000000001010111100010000",
			554 => "0000000100000000001011100100000100",
			555 => "11111110101010000000100011111101",
			556 => "0000000111000000000100010100001000",
			557 => "0000000101000000001000111000000100",
			558 => "11111111100110100000100011111101",
			559 => "00000001100111110000100011111101",
			560 => "00000011110110100000100011111101",
			561 => "11111110011010110000100011111101",
			562 => "0000000100000000000011011000001100",
			563 => "0000000110000000001110010100001000",
			564 => "0000000110000000001011111100000100",
			565 => "11111110011110010000100011111101",
			566 => "00000001110110000000100011111101",
			567 => "11111110011001010000100011111101",
			568 => "0000000110000000001101111100001100",
			569 => "0000000101000000001100101000000100",
			570 => "11111110011001110000100011111101",
			571 => "0000001011000000000111001000000100",
			572 => "00000110010100110000100011111101",
			573 => "11111110100111010000100011111101",
			574 => "11111110011001010000100011111101",
			575 => "0000000011000000001000101100010100",
			576 => "0000000110000000001101111100010000",
			577 => "0000000110000000001110010100000100",
			578 => "11111110100010000000100110000001",
			579 => "0000000010000000001110010000001000",
			580 => "0000000000000000000101001000000100",
			581 => "00000001101101000000100110000001",
			582 => "11111111100011000000100110000001",
			583 => "00000110001001010000100110000001",
			584 => "11111110101101010000100110000001",
			585 => "0000000001000000000000011000100000",
			586 => "0000000010000000000111100000001100",
			587 => "0000000011000000000011111100001000",
			588 => "0000000110000000001101111100000100",
			589 => "00000001010001000000100110000001",
			590 => "11111111010001000000100110000001",
			591 => "00000011001110000000100110000001",
			592 => "0000001001000000001110100000001100",
			593 => "0000000010000000000101001000001000",
			594 => "0000000010000000000101001000000100",
			595 => "11111111000011010000100110000001",
			596 => "00000000110001000000100110000001",
			597 => "11111110011001100000100110000001",
			598 => "0000001100000000001010000000000100",
			599 => "00000000000000000000100110000001",
			600 => "00000010000011100000100110000001",
			601 => "0000000100000000001101110100000100",
			602 => "11111110011010000000100110000001",
			603 => "0000000110000000001101111100001000",
			604 => "0000000110000000000111101000000100",
			605 => "00000000000000000000100110000001",
			606 => "00000001100000010000100110000001",
			607 => "11111110011010100000100110000001",
			608 => "0000000100000000000011011000010000",
			609 => "0000000110000000001110010100001100",
			610 => "0000000010000000001110101000000100",
			611 => "00000000000000000000100111100101",
			612 => "0000000011000000000001111100000100",
			613 => "00000000000000000000100111100101",
			614 => "00000000010001100000100111100101",
			615 => "11111110100010000000100111100101",
			616 => "0000000110000000001101111100100000",
			617 => "0000000111000000001110001100011100",
			618 => "0000000100000000000000101100001100",
			619 => "0000001000000000001001101000001000",
			620 => "0000001010000000001000100100000100",
			621 => "00000000000000000000100111100101",
			622 => "00000000011111110000100111100101",
			623 => "11111111101010010000100111100101",
			624 => "0000000110000000001110010100000100",
			625 => "00000000000000000000100111100101",
			626 => "0000000010000000001110110100001000",
			627 => "0000001000000000001011000100000100",
			628 => "00000001000101010000100111100101",
			629 => "00000000000000000000100111100101",
			630 => "00000000000000000000100111100101",
			631 => "00000000000000000000100111100101",
			632 => "11111111010000000000100111100101",
			633 => "0000000011000000000111000000001100",
			634 => "0000000110000000001101111100001000",
			635 => "0000000110000000000111101000000100",
			636 => "00000000000000000000101001100001",
			637 => "00000001101001100000101001100001",
			638 => "11111111000010010000101001100001",
			639 => "0000000100000000000011011000001100",
			640 => "0000001000000000000110011000001000",
			641 => "0000000000000000001001101000000100",
			642 => "11111110011110000000101001100001",
			643 => "00000101101110010000101001100001",
			644 => "11111110011001010000101001100001",
			645 => "0000000010000000001110000100011000",
			646 => "0000000110000000001101111100010100",
			647 => "0000001100000000000000101000001100",
			648 => "0000000001000000000000011000001000",
			649 => "0000000110000000000111101000000100",
			650 => "00000000000000000000101001100001",
			651 => "00000001101110100000101001100001",
			652 => "11111110111001110000101001100001",
			653 => "0000000001000000001110011100000100",
			654 => "00000000000000000000101001100001",
			655 => "00000010110011110000101001100001",
			656 => "11111111000110100000101001100001",
			657 => "0000000110000000001101111100001100",
			658 => "0000000110000000000001111000000100",
			659 => "11111110100100100000101001100001",
			660 => "0000000100000000001111110100000100",
			661 => "00000001100110100000101001100001",
			662 => "11111111011111010000101001100001",
			663 => "11111110011011010000101001100001",
			664 => "0000001110000000000001110000010100",
			665 => "0000000110000000001101111100010000",
			666 => "0000001111000000001010111000001100",
			667 => "0000000000000000000111100000001000",
			668 => "0000000100000000000000000100000100",
			669 => "00000000000000000000101011101101",
			670 => "00000001101000100000101011101101",
			671 => "00000000000000000000101011101101",
			672 => "11111111100000100000101011101101",
			673 => "11111110111111000000101011101101",
			674 => "0000000100000000000011011000001100",
			675 => "0000000110000000001110010100001000",
			676 => "0000000110000000001011111100000100",
			677 => "11111110101000000000101011101101",
			678 => "00000000011010000000101011101101",
			679 => "11111110011001110000101011101101",
			680 => "0000001000000000001111001000001100",
			681 => "0000000011000000000100011000000100",
			682 => "11111111111110100000101011101101",
			683 => "0000001100000000001100110000000100",
			684 => "00000010011101000000101011101101",
			685 => "00000000000000000000101011101101",
			686 => "0000000010000000001110101000001100",
			687 => "0000000001000000001100100000001000",
			688 => "0000000000000000000101001000000100",
			689 => "00000001100100000000101011101101",
			690 => "00000000000000000000101011101101",
			691 => "11111111000011010000101011101101",
			692 => "0000000110000000001101111100001100",
			693 => "0000000110000000001101111100000100",
			694 => "11111110111010100000101011101101",
			695 => "0000000101000000000001101000000100",
			696 => "00000000100101100000101011101101",
			697 => "00000000000000000000101011101101",
			698 => "11111110011101110000101011101101",
			699 => "0000000011000000001000101100010100",
			700 => "0000000110000000001101111100010000",
			701 => "0000000110000000001110010100000100",
			702 => "11111110011111100000101110000011",
			703 => "0000000000000000000101001000001000",
			704 => "0000000010000000001110010000000100",
			705 => "00000001110110000000101110000011",
			706 => "00000000000000110000101110000011",
			707 => "11111111001101000000101110000011",
			708 => "11111110011111110000101110000011",
			709 => "0000001111000000001010111000010000",
			710 => "0000001101000000001100101100001100",
			711 => "0000000001000000001100100000001000",
			712 => "0000000101000000001001110000000100",
			713 => "00000000000000000000101110000011",
			714 => "00000010111010100000101110000011",
			715 => "11111110101001000000101110000011",
			716 => "11111110011010010000101110000011",
			717 => "0000000100000000000011011000001100",
			718 => "0000000110000000001110010100001000",
			719 => "0000000110000000001011111100000100",
			720 => "11111110011101100000101110000011",
			721 => "00000001111010110000101110000011",
			722 => "11111110011000010000101110000011",
			723 => "0000000010000000000111100000001000",
			724 => "0000000110000000001101111100000100",
			725 => "00000001100111010000101110000011",
			726 => "11111111011111100000101110000011",
			727 => "0000000010000000001110110100010000",
			728 => "0000000010000000001110110100001000",
			729 => "0000000100000000001010010000000100",
			730 => "11111110011011010000101110000011",
			731 => "11111111011100010000101110000011",
			732 => "0000000100000000000001001100000100",
			733 => "00000100011000010000101110000011",
			734 => "11111110111001110000101110000011",
			735 => "11111110011001000000101110000011",
			736 => "00000000000000000000101110000101",
			737 => "00000000000000000000101110001001",
			738 => "00000000000000000000101110001101",
			739 => "00000000000000000000101110010001",
			740 => "00000000000000000000101110010101",
			741 => "00000000000000000000101110011001",
			742 => "00000000000000000000101110011101",
			743 => "00000000000000000000101110100001",
			744 => "00000000000000000000101110100101",
			745 => "00000000000000000000101110101001",
			746 => "00000000000000000000101110101101",
			747 => "00000000000000000000101110110001",
			748 => "00000000000000000000101110110101",
			749 => "00000000000000000000101110111001",
			750 => "00000000000000000000101110111101",
			751 => "00000000000000000000101111000001",
			752 => "00000000000000000000101111000101",
			753 => "00000000000000000000101111001001",
			754 => "00000000000000000000101111001101",
			755 => "00000000000000000000101111010001",
			756 => "00000000000000000000101111010101",
			757 => "00000000000000000000101111011001",
			758 => "00000000000000000000101111011101",
			759 => "00000000000000000000101111100001",
			760 => "00000000000000000000101111100101",
			761 => "00000000000000000000101111101001",
			762 => "00000000000000000000101111101101",
			763 => "00000000000000000000101111110001",
			764 => "00000000000000000000101111110101",
			765 => "0000000100000000000011011000000100",
			766 => "11111111101010110000110000000001",
			767 => "00000000000000000000110000000001",
			768 => "0000000010000000000111100000000100",
			769 => "00000000000000000000110000001101",
			770 => "11111111111110100000110000001101",
			771 => "0000000011000000001010101100000100",
			772 => "00000000000000000000110000011001",
			773 => "11111111110110000000110000011001",
			774 => "0000000010000000001100100100000100",
			775 => "00000000000000000000110000100101",
			776 => "11111111111010110000110000100101",
			777 => "0000000110000000001101111100001000",
			778 => "0000000110000000000111101000000100",
			779 => "00000000000000000000110000111001",
			780 => "00000000000101000000110000111001",
			781 => "11111111111000000000110000111001",
			782 => "0000000110000000001101111100001000",
			783 => "0000000110000000001011111100000100",
			784 => "00000000000000000000110001001101",
			785 => "00000000000111000000110001001101",
			786 => "00000000000000000000110001001101",
			787 => "0000000110000000001101111100001000",
			788 => "0000000110000000001011111100000100",
			789 => "00000000000000000000110001100001",
			790 => "00000000000101110000110001100001",
			791 => "00000000000000000000110001100001",
			792 => "0000000100000000001011100100001000",
			793 => "0000000011000000000100011000000100",
			794 => "11111111101111100000110001110101",
			795 => "00000000000000000000110001110101",
			796 => "00000000000000000000110001110101",
			797 => "0000000110000000001101111100001000",
			798 => "0000000110000000001011111100000100",
			799 => "00000000000000000000110010001001",
			800 => "00000000000011110000110010001001",
			801 => "00000000000000000000110010001001",
			802 => "0000000110000000001101111100001000",
			803 => "0000000110000000001011111100000100",
			804 => "00000000000000000000110010011101",
			805 => "00000000000100010000110010011101",
			806 => "00000000000000000000110010011101",
			807 => "0000000010000000001100100100000100",
			808 => "00000000000000000000110010110001",
			809 => "0000000011000000000111000000000100",
			810 => "00000000000000000000110010110001",
			811 => "11111111111010100000110010110001",
			812 => "0000000110000000001101111100001000",
			813 => "0000000110000000001011111100000100",
			814 => "00000000000000000000110011000101",
			815 => "00000000000011100000110011000101",
			816 => "00000000000000000000110011000101",
			817 => "0000000110000000001101111100001000",
			818 => "0000000110000000001011111100000100",
			819 => "00000000000000000000110011011001",
			820 => "00000000000111000000110011011001",
			821 => "00000000000000000000110011011001",
			822 => "0000000110000000001101111100001000",
			823 => "0000000110000000001011111100000100",
			824 => "00000000000000000000110011101101",
			825 => "00000000000011000000110011101101",
			826 => "00000000000000000000110011101101",
			827 => "0000000110000000001101111100001000",
			828 => "0000000110000000001011111100000100",
			829 => "00000000000000000000110100000001",
			830 => "00000000000110000000110100000001",
			831 => "00000000000000000000110100000001",
			832 => "0000000100000000000101100000001100",
			833 => "0000001111000000000011011100000100",
			834 => "00000000000000000000110100011101",
			835 => "0000000101000000000110100100000100",
			836 => "11111111001010010000110100011101",
			837 => "00000000000000000000110100011101",
			838 => "00000000000000000000110100011101",
			839 => "0000000110000000001101111100001100",
			840 => "0000000110000000001011111100000100",
			841 => "00000000000000000000110100111001",
			842 => "0000000110000000001101111100000100",
			843 => "00000000001010110000110100111001",
			844 => "00000000000000000000110100111001",
			845 => "11111111111000000000110100111001",
			846 => "0000000010000000000111100000001100",
			847 => "0000000110000000001101111100001000",
			848 => "0000000110000000001011111100000100",
			849 => "00000000000000000000110101011101",
			850 => "00000000010000010000110101011101",
			851 => "00000000000000000000110101011101",
			852 => "0000000010000000001000001100000100",
			853 => "11111111100111000000110101011101",
			854 => "00000000000000000000110101011101",
			855 => "0000000110000000001101111100010000",
			856 => "0000000011000000000100011000000100",
			857 => "00000000000000000000110110000001",
			858 => "0000000000000000001011010100000100",
			859 => "00000000000000000000110110000001",
			860 => "0000001101000000001011000000000100",
			861 => "00000000000000000000110110000001",
			862 => "00000000011000110000110110000001",
			863 => "11111111100111010000110110000001",
			864 => "0000000100000000000011011000000100",
			865 => "11111111011001000000110110100101",
			866 => "0000001100000000000011011100001100",
			867 => "0000000010000000001110110100001000",
			868 => "0000001000000000000100010100000100",
			869 => "00000000010010010000110110100101",
			870 => "00000000000000000000110110100101",
			871 => "00000000000000000000110110100101",
			872 => "00000000000000000000110110100101",
			873 => "0000000010000000000111100000010000",
			874 => "0000000001000000001100110100001100",
			875 => "0000000100000000001111101000000100",
			876 => "00000000000000000000110111010001",
			877 => "0000000100000000001101110000000100",
			878 => "00000000000011110000110111010001",
			879 => "00000000000000000000110111010001",
			880 => "00000000000000000000110111010001",
			881 => "0000000011000000000111000000000100",
			882 => "00000000000000000000110111010001",
			883 => "11111111110000010000110111010001",
			884 => "0000000110000000001101111100010000",
			885 => "0000000110000000001011111100000100",
			886 => "00000000000000000000110111111101",
			887 => "0000000000000000001011010100000100",
			888 => "00000000000000000000110111111101",
			889 => "0000001000000000000100010100000100",
			890 => "00000000001001000000110111111101",
			891 => "00000000000000000000110111111101",
			892 => "0000000011000000000111000100000100",
			893 => "00000000000000000000110111111101",
			894 => "11111111110000010000110111111101",
			895 => "0000000011000000000111000000001100",
			896 => "0000000110000000001101111100001000",
			897 => "0000001111000000000111001000000100",
			898 => "00000100010110100000111000110001",
			899 => "11111110100110010000111000110001",
			900 => "11111110011001110000111000110001",
			901 => "0000001111000000000001111100001100",
			902 => "0000000101000000001010111100001000",
			903 => "0000000001000000001100100000000100",
			904 => "00000100011001010000111000110001",
			905 => "11111110100001000000111000110001",
			906 => "11111110010110010000111000110001",
			907 => "11111110010101100000111000110001",
			908 => "0000000011000000000111000000010000",
			909 => "0000000110000000001101111100001100",
			910 => "0000001111000000000111001000001000",
			911 => "0000001010000000000001110100000100",
			912 => "00000010111110010000111001101101",
			913 => "00000000111011110000111001101101",
			914 => "11111110110001100000111001101101",
			915 => "11111110011001110000111001101101",
			916 => "0000001111000000000001111100001100",
			917 => "0000001011000000000000101000001000",
			918 => "0000000001000000001100100000000100",
			919 => "00000010111100100000111001101101",
			920 => "11111110100111010000111001101101",
			921 => "11111110010111100000111001101101",
			922 => "11111110010111010000111001101101",
			923 => "0000000010000000000111100000010100",
			924 => "0000000001000000001100110100010000",
			925 => "0000000110000000001101111100001100",
			926 => "0000000110000000001011111100000100",
			927 => "00000000000000000000111010100001",
			928 => "0000000100000000001101110000000100",
			929 => "00000000001001010000111010100001",
			930 => "00000000000000000000111010100001",
			931 => "00000000000000000000111010100001",
			932 => "00000000000000000000111010100001",
			933 => "0000000011000000000111000000000100",
			934 => "00000000000000000000111010100001",
			935 => "11111111101110110000111010100001",
			936 => "0000000100000000000011011000000100",
			937 => "11111110110101100000111011001101",
			938 => "0000000111000000000110000100010000",
			939 => "0000000110000000001101111100001100",
			940 => "0000000110000000000111101000000100",
			941 => "00000000000000000000111011001101",
			942 => "0000001000000000001011000100000100",
			943 => "00000000101000010000111011001101",
			944 => "00000000000000000000111011001101",
			945 => "00000000000000000000111011001101",
			946 => "00000000000000000000111011001101",
			947 => "0000000011000000000111000000010000",
			948 => "0000000110000000001101111100001100",
			949 => "0000001111000000000111001000001000",
			950 => "0000001101000000001101100000000100",
			951 => "00000010101000000000111100010001",
			952 => "00000000101110110000111100010001",
			953 => "11111110110110110000111100010001",
			954 => "11111110011011110000111100010001",
			955 => "0000001111000000000001111100001100",
			956 => "0000001011000000000000101000001000",
			957 => "0000000001000000001100100000000100",
			958 => "00000010100110000000111100010001",
			959 => "11111110101001100000111100010001",
			960 => "11111110011000000000111100010001",
			961 => "0000000110000000001101111100000100",
			962 => "11111110011100010000111100010001",
			963 => "11111110010110100000111100010001",
			964 => "0000000100000000000011011000001000",
			965 => "0000000110000000001110010100000100",
			966 => "00000000000000000000111101010101",
			967 => "11111110110000110000111101010101",
			968 => "0000000010000000000111100000010000",
			969 => "0000000110000000001101111100001100",
			970 => "0000000100000000001101110000001000",
			971 => "0000000110000000000111101000000100",
			972 => "00000000000000000000111101010101",
			973 => "00000000110110100000111101010101",
			974 => "00000000000000000000111101010101",
			975 => "00000000000000000000111101010101",
			976 => "0000001000000000000110001000000100",
			977 => "00000000000000000000111101010101",
			978 => "0000000011000000000111000000000100",
			979 => "00000000000000000000111101010101",
			980 => "11111111100110100000111101010101",
			981 => "0000000011000000001010101100001100",
			982 => "0000001010000000000010101000001000",
			983 => "0000001001000000000000011000000100",
			984 => "00000110000101010000111110100001",
			985 => "00000100001111010000111110100001",
			986 => "11111110101010010000111110100001",
			987 => "0000000011000000001000101100001100",
			988 => "0000000000000000001001001000001000",
			989 => "0000000101000000001000111000000100",
			990 => "11111110100001000000111110100001",
			991 => "00000111011000010000111110100001",
			992 => "11111110010111110000111110100001",
			993 => "0000001111000000000001111100001100",
			994 => "0000001011000000000000101000001000",
			995 => "0000001001000000000110000000000100",
			996 => "00000110001101100000111110100001",
			997 => "11111110100001000000111110100001",
			998 => "11111110010101100000111110100001",
			999 => "11111110010100100000111110100001",
			1000 => "0000000001000000000000011000010100",
			1001 => "0000000101000000001010111000010000",
			1002 => "0000000110000000001101111100001100",
			1003 => "0000000110000000000111101000000100",
			1004 => "00000000000000000000111111101101",
			1005 => "0000000010000000000011001000000100",
			1006 => "00000001100000100000111111101101",
			1007 => "00000000000000000000111111101101",
			1008 => "11111111101001000000111111101101",
			1009 => "11111111000101000000111111101101",
			1010 => "0000001000000000000110011000001000",
			1011 => "0000000010000000000111010100000100",
			1012 => "11111110111110110000111111101101",
			1013 => "00000001011101110000111111101101",
			1014 => "0000001101000000001001110100000100",
			1015 => "11111110011100010000111111101101",
			1016 => "0000001101000000001001110100000100",
			1017 => "00000000100101010000111111101101",
			1018 => "11111110110100100000111111101101",
			1019 => "0000000110000000001101111100011100",
			1020 => "0000000011000000000100011000010000",
			1021 => "0000000000000000001001110000000100",
			1022 => "11111110110010000001000000101001",
			1023 => "0000000010000000000111100000001000",
			1024 => "0000000000000000001100100100000100",
			1025 => "00000000111001110001000000101001",
			1026 => "00000000000000000001000000101001",
			1027 => "00000000000000000001000000101001",
			1028 => "0000000000000000001011010100000100",
			1029 => "00000000000000000001000000101001",
			1030 => "0000001101000000001001001000000100",
			1031 => "00000000000000000001000000101001",
			1032 => "00000001011011010001000000101001",
			1033 => "11111110100101110001000000101001",
			1034 => "0000000110000000001101111100011100",
			1035 => "0000001101000000001010111100010000",
			1036 => "0000001001000000000110000000001100",
			1037 => "0000001111000000001010111000001000",
			1038 => "0000000110000000001110010100000100",
			1039 => "00000000000000000001000001100101",
			1040 => "00000000010100000001000001100101",
			1041 => "00000000000000000001000001100101",
			1042 => "11111111010011100001000001100101",
			1043 => "0000001001000000001110100000000100",
			1044 => "00000000000000000001000001100101",
			1045 => "0000000100000000001111101000000100",
			1046 => "00000000000000000001000001100101",
			1047 => "00000001001010110001000001100101",
			1048 => "11111111001000010001000001100101",
			1049 => "0000000110000000001101111100011100",
			1050 => "0000001101000000001010111100001100",
			1051 => "0000001001000000000110000000001000",
			1052 => "0000001010000000000110011100000100",
			1053 => "00000000000000000001000010100001",
			1054 => "00000000000011100001000010100001",
			1055 => "11111111100110110001000010100001",
			1056 => "0000000100000000001011110000000100",
			1057 => "00000000000000000001000010100001",
			1058 => "0000001001000000001110100000000100",
			1059 => "00000000000000000001000010100001",
			1060 => "0000000110000000000001111000000100",
			1061 => "00000000000000000001000010100001",
			1062 => "00000000100100010001000010100001",
			1063 => "11111111011001110001000010100001",
			1064 => "0000001001000000001100110100011100",
			1065 => "0000000011000000000001110100001000",
			1066 => "0000001111000000001101111000000100",
			1067 => "00000001010111100001000011110101",
			1068 => "00000000000000000001000011110101",
			1069 => "0000000101000000000011011100001000",
			1070 => "0000001001000000000000011000000100",
			1071 => "00000000000000000001000011110101",
			1072 => "11111111001100010001000011110101",
			1073 => "0000000101000000001010111000001000",
			1074 => "0000001010000000000110011100000100",
			1075 => "00000000000000000001000011110101",
			1076 => "00000001001101010001000011110101",
			1077 => "11111111010111110001000011110101",
			1078 => "0000001101000000001010011100000100",
			1079 => "11111110011101000001000011110101",
			1080 => "0000000110000000001101111100001000",
			1081 => "0000000000000000001001101000000100",
			1082 => "11111111110111000001000011110101",
			1083 => "00000001101000000001000011110101",
			1084 => "11111110101100010001000011110101",
			1085 => "0000001101000000001001110100001100",
			1086 => "0000000100000000000100111000001000",
			1087 => "0000001001000000000000011000000100",
			1088 => "00000000000000000001000100111001",
			1089 => "11111111001001100001000100111001",
			1090 => "00000000000000000001000100111001",
			1091 => "0000001100000000000100001000010100",
			1092 => "0000001010000000000001010000010000",
			1093 => "0000000100000000001111101000000100",
			1094 => "00000000000000000001000100111001",
			1095 => "0000000001000000001101101000001000",
			1096 => "0000001100000000000100000000000100",
			1097 => "00000000000000000001000100111001",
			1098 => "00000000100110100001000100111001",
			1099 => "00000000000000000001000100111001",
			1100 => "00000000000000000001000100111001",
			1101 => "00000000000000000001000100111001",
			1102 => "0000000100000000000011011000000100",
			1103 => "11111110011111100001000101110101",
			1104 => "0000001100000000000011011100011000",
			1105 => "0000001101000000001010111100010000",
			1106 => "0000000100000000000101100000001000",
			1107 => "0000000001000000001100100000000100",
			1108 => "00000000000000000001000101110101",
			1109 => "11111110111101110001000101110101",
			1110 => "0000001111000000001010111000000100",
			1111 => "00000001001011010001000101110101",
			1112 => "00000000000000000001000101110101",
			1113 => "0000000010000000001110110100000100",
			1114 => "00000001010110110001000101110101",
			1115 => "00000000000000000001000101110101",
			1116 => "11111111010011110001000101110101",
			1117 => "0000000110000000001101111100100000",
			1118 => "0000000101000000001100101000010000",
			1119 => "0000001111000000001010111000001100",
			1120 => "0000001010000000000110011100000100",
			1121 => "00000000000000000001000110111001",
			1122 => "0000000110000000000111101000000100",
			1123 => "00000000000000000001000110111001",
			1124 => "00000000101111000001000110111001",
			1125 => "11111110111100010001000110111001",
			1126 => "0000000100000000001111101000000100",
			1127 => "00000000000000000001000110111001",
			1128 => "0000000001000000000000011000000100",
			1129 => "00000000000000000001000110111001",
			1130 => "0000001011000000001000111000000100",
			1131 => "00000000000000000001000110111001",
			1132 => "00000001010100110001000110111001",
			1133 => "11111110110010000001000110111001",
			1134 => "0000001110000000000101000100010000",
			1135 => "0000001111000000001010111000001100",
			1136 => "0000000100000000000101001100000100",
			1137 => "00000000000000000001001000001101",
			1138 => "0000001010000000000010101000000100",
			1139 => "00000000101000000001001000001101",
			1140 => "00000000000000000001001000001101",
			1141 => "00000000000000000001001000001101",
			1142 => "0000001101000000001010011100001000",
			1143 => "0000000001000000001100100000000100",
			1144 => "00000000000000000001001000001101",
			1145 => "11111110101000010001001000001101",
			1146 => "0000001100000000000100001000010000",
			1147 => "0000001010000000001001000100001100",
			1148 => "0000000100000000001011110000000100",
			1149 => "00000000000000000001001000001101",
			1150 => "0000000001000000001101011100000100",
			1151 => "00000000111101110001001000001101",
			1152 => "00000000000000000001001000001101",
			1153 => "00000000000000000001001000001101",
			1154 => "11111111100101100001001000001101",
			1155 => "0000000110000000001101111100100000",
			1156 => "0000000011000000000100011000010100",
			1157 => "0000001010000000000110011100000100",
			1158 => "11111111010111000001001001010001",
			1159 => "0000000010000000000111100000001100",
			1160 => "0000000100000000001011100100000100",
			1161 => "00000000000000000001001001010001",
			1162 => "0000000000000000000001001000000100",
			1163 => "00000000011110110001001001010001",
			1164 => "00000000000000000001001001010001",
			1165 => "00000000000000000001001001010001",
			1166 => "0000000100000000001111101000000100",
			1167 => "00000000000000000001001001010001",
			1168 => "0000000101000000000111001000000100",
			1169 => "00000000000000000001001001010001",
			1170 => "00000000111100010001001001010001",
			1171 => "11111111001110000001001001010001",
			1172 => "0000000011000000000111000000001100",
			1173 => "0000001000000000000100000000001000",
			1174 => "0000000110000000000111101000000100",
			1175 => "00000000111100100001001010101101",
			1176 => "00000010001101010001001010101101",
			1177 => "11111110100000010001001010101101",
			1178 => "0000001111000000001101010100010000",
			1179 => "0000001100000000001100001000001100",
			1180 => "0000000100000000001101000000000100",
			1181 => "11111110100111000001001010101101",
			1182 => "0000000110000000000001111000000100",
			1183 => "00000010000011110001001010101101",
			1184 => "00000011011110010001001010101101",
			1185 => "11111110011000110001001010101101",
			1186 => "0000000100000000000011011000000100",
			1187 => "11111110010111010001001010101101",
			1188 => "0000000110000000001101111100001100",
			1189 => "0000000110000000000001111000000100",
			1190 => "11111110011010010001001010101101",
			1191 => "0000000100000000001111011000000100",
			1192 => "00000101000100010001001010101101",
			1193 => "11111110011111110001001010101101",
			1194 => "11111110010111110001001010101101",
			1195 => "0000001110000000000001010100011000",
			1196 => "0000000110000000001101111100010000",
			1197 => "0000001111000000001010111000001100",
			1198 => "0000000100000000000101001100000100",
			1199 => "00000000000000000001001100001001",
			1200 => "0000001000000000001011000100000100",
			1201 => "00000001100110100001001100001001",
			1202 => "00000000000000000001001100001001",
			1203 => "11111111110100110001001100001001",
			1204 => "0000000110000000001101111100000100",
			1205 => "00000000000000000001001100001001",
			1206 => "11111111010101010001001100001001",
			1207 => "0000000100000000000011011000000100",
			1208 => "11111110011010000001001100001001",
			1209 => "0000000110000000001101111100010000",
			1210 => "0000000011000000001100101100001100",
			1211 => "0000001111000000001101010100001000",
			1212 => "0000000100000000001101100100000100",
			1213 => "00000000111110100001001100001001",
			1214 => "00000000000000000001001100001001",
			1215 => "11111110101111000001001100001001",
			1216 => "00000001110011110001001100001001",
			1217 => "11111110100010000001001100001001",
			1218 => "0000001101000000001001110100011000",
			1219 => "0000000100000000000100111000001000",
			1220 => "0000000001000000001100100000000100",
			1221 => "00000000000000000001001101100101",
			1222 => "11111110100110100001001101100101",
			1223 => "0000000010000000000011001000001100",
			1224 => "0000000100000000000101100000000100",
			1225 => "00000000000000000001001101100101",
			1226 => "0000000101000000001110110000000100",
			1227 => "00000000110011000001001101100101",
			1228 => "00000000000000000001001101100101",
			1229 => "00000000000000000001001101100101",
			1230 => "0000001100000000000100001000010100",
			1231 => "0000001010000000000001010000010000",
			1232 => "0000000100000000001111101000000100",
			1233 => "00000000000000000001001101100101",
			1234 => "0000000001000000001101101000001000",
			1235 => "0000001100000000000100000000000100",
			1236 => "00000000000000000001001101100101",
			1237 => "00000001001011100001001101100101",
			1238 => "00000000000000000001001101100101",
			1239 => "00000000000000000001001101100101",
			1240 => "11111111100111110001001101100101",
			1241 => "0000000100000000000011011000001100",
			1242 => "0000001000000000000110011000001000",
			1243 => "0000000000000000001001101000000100",
			1244 => "11111111001000110001001110110001",
			1245 => "00000001011101110001001110110001",
			1246 => "11111110011100100001001110110001",
			1247 => "0000000110000000001101111100011000",
			1248 => "0000000111000000001110001100010100",
			1249 => "0000000110000000001110010100000100",
			1250 => "00000000000000000001001110110001",
			1251 => "0000000001000000000000011000001000",
			1252 => "0000000010000000000011001000000100",
			1253 => "00000001100000110001001110110001",
			1254 => "00000000000000000001001110110001",
			1255 => "0000000001000000000110000000000100",
			1256 => "11111111101010100001001110110001",
			1257 => "00000000110011010001001110110001",
			1258 => "11111111111101010001001110110001",
			1259 => "11111110110100000001001110110001",
			1260 => "0000000001000000000000011000010100",
			1261 => "0000000101000000001010111000010000",
			1262 => "0000000100000000001011100100000100",
			1263 => "11111111110011110001010000010101",
			1264 => "0000001010000000000110011100000100",
			1265 => "00000000000000000001010000010101",
			1266 => "0000001111000000001010011100000100",
			1267 => "00000001011001110001010000010101",
			1268 => "00000000000000000001010000010101",
			1269 => "11111111000000000001010000010101",
			1270 => "0000001000000000000110011000001100",
			1271 => "0000001111000000000111010100000100",
			1272 => "11111110111100000001010000010101",
			1273 => "0000001101000000001110010000000100",
			1274 => "00000001101010100001010000010101",
			1275 => "00000000000000000001010000010101",
			1276 => "0000000100000000001101110100000100",
			1277 => "11111110011011110001010000010101",
			1278 => "0000000100000000000000100000000100",
			1279 => "00000000010011100001010000010101",
			1280 => "0000000100000000000001100100001000",
			1281 => "0000000100000000000000101100000100",
			1282 => "11111111111010110001010000010101",
			1283 => "00000000000000000001010000010101",
			1284 => "11111110111011010001010000010101",
			1285 => "0000000011000000000111000000001100",
			1286 => "0000000110000000001101111100001000",
			1287 => "0000000110000000000111101000000100",
			1288 => "00000000000000000001010010000001",
			1289 => "00000001101010010001010010000001",
			1290 => "11111110111110100001010010000001",
			1291 => "0000000100000000000011011000001100",
			1292 => "0000001000000000000110011000001000",
			1293 => "0000000100000000001000100000000100",
			1294 => "11111110011101010001010010000001",
			1295 => "00001000011100010001010010000001",
			1296 => "11111110011001010001010010000001",
			1297 => "0000000010000000001110000100010000",
			1298 => "0000001011000000001100001000001000",
			1299 => "0000001111000000001010111100000100",
			1300 => "00000001010110000001010010000001",
			1301 => "11111110101110000001010010000001",
			1302 => "0000001001000000001100100000000100",
			1303 => "11111111011001000001010010000001",
			1304 => "00000010111101110001010010000001",
			1305 => "0000000110000000001101111100001100",
			1306 => "0000000110000000000001111000000100",
			1307 => "11111110100010000001010010000001",
			1308 => "0000000100000000001111110100000100",
			1309 => "00000001110011010001010010000001",
			1310 => "11111111011000000001010010000001",
			1311 => "11111110011010110001010010000001",
			1312 => "0000000011000000000111000000010000",
			1313 => "0000000110000000001101111100001000",
			1314 => "0000000110000000000111101000000100",
			1315 => "00000000000000000001010011110101",
			1316 => "00000001101000110001010011110101",
			1317 => "0000000011000000001010101100000100",
			1318 => "00000000000000000001010011110101",
			1319 => "11111111000000000001010011110101",
			1320 => "0000000100000000000011011000001100",
			1321 => "0000000000000000001011010100001000",
			1322 => "0000000100000000001101101100000100",
			1323 => "11111110011101110001010011110101",
			1324 => "00000100011001000001010011110101",
			1325 => "11111110011001100001010011110101",
			1326 => "0000000000000000000011010000001000",
			1327 => "0000001100000000001100110000000100",
			1328 => "00000011010001000001010011110101",
			1329 => "00000000000000000001010011110101",
			1330 => "0000000110000000001101111100010100",
			1331 => "0000000110000000000001111000001000",
			1332 => "0000001111000000001010111100000100",
			1333 => "00000000100010000001010011110101",
			1334 => "11111110100101000001010011110101",
			1335 => "0000000111000000001101111000001000",
			1336 => "0000000111000000001011000100000100",
			1337 => "00000000000000000001010011110101",
			1338 => "00000001110010100001010011110101",
			1339 => "11111111001110110001010011110101",
			1340 => "11111110011011110001010011110101",
			1341 => "0000000011000000000111000000010100",
			1342 => "0000000110000000001101111100001100",
			1343 => "0000000110000000000111101000000100",
			1344 => "00000000000000000001010101101001",
			1345 => "0000001010000000000111000100000100",
			1346 => "00000001101001000001010101101001",
			1347 => "00000000000000000001010101101001",
			1348 => "0000000011000000001010101100000100",
			1349 => "00000000000000000001010101101001",
			1350 => "11111111000011100001010101101001",
			1351 => "0000000110000000001101111100100100",
			1352 => "0000001101000000001010011100011000",
			1353 => "0000001010000000000001010100001000",
			1354 => "0000001111000000000110000100000100",
			1355 => "00000000000000000001010101101001",
			1356 => "11111110011010000001010101101001",
			1357 => "0000000000000000001110110000001100",
			1358 => "0000001111000000001110110000000100",
			1359 => "00000001011001100001010101101001",
			1360 => "0000001111000000001000011000000100",
			1361 => "11111111100010110001010101101001",
			1362 => "00000000110011010001010101101001",
			1363 => "11111111011110110001010101101001",
			1364 => "0000000000000000001011010100000100",
			1365 => "11111110100100010001010101101001",
			1366 => "0000001111000000001011011100000100",
			1367 => "11111111011100000001010101101001",
			1368 => "00000011011001000001010101101001",
			1369 => "11111110011001110001010101101001",
			1370 => "0000000011000000001000101100011000",
			1371 => "0000000110000000001110010100000100",
			1372 => "11111110100111010001010111100101",
			1373 => "0000000110000000001101111100010000",
			1374 => "0000000100000000001111111000001100",
			1375 => "0000001111000000001110110000001000",
			1376 => "0000001101000000000011011100000100",
			1377 => "00000001101010100001010111100101",
			1378 => "00000010111111000001010111100101",
			1379 => "00000000000000000001010111100101",
			1380 => "11111111110101000001010111100101",
			1381 => "11111110110011100001010111100101",
			1382 => "0000001111000000001010111000010000",
			1383 => "0000001100000000001100001000001100",
			1384 => "0000000001000000001100100000001000",
			1385 => "0000000110000000000111101000000100",
			1386 => "00000000000000000001010111100101",
			1387 => "00000010001010110001010111100101",
			1388 => "11111110110110100001010111100101",
			1389 => "11111110011110010001010111100101",
			1390 => "0000000100000000001101110100000100",
			1391 => "11111110011010100001010111100101",
			1392 => "0000000110000000001101111100010000",
			1393 => "0000001001000000001110100000000100",
			1394 => "11111110011101100001010111100101",
			1395 => "0000001111000000000001101000000100",
			1396 => "11111110101001100001010111100101",
			1397 => "0000000110000000001110010100000100",
			1398 => "00000000000000000001010111100101",
			1399 => "00000010110101010001010111100101",
			1400 => "11111110011011000001010111100101",
			1401 => "0000000011000000001000101100010100",
			1402 => "0000001000000000000100000000010000",
			1403 => "0000000100000000000101100000000100",
			1404 => "11111111000101000001011001101001",
			1405 => "0000001111000000001010111000001000",
			1406 => "0000001011000000001011000100000100",
			1407 => "00000001101011100001011001101001",
			1408 => "00000011000000110001011001101001",
			1409 => "11111111011100010001011001101001",
			1410 => "11111110110011100001011001101001",
			1411 => "0000001111000000001010111000010000",
			1412 => "0000001100000000001100001000001100",
			1413 => "0000000001000000001100100000001000",
			1414 => "0000001100000000001010000000000100",
			1415 => "00000000000000000001011001101001",
			1416 => "00000010010010010001011001101001",
			1417 => "11111110110100000001011001101001",
			1418 => "11111110011101010001011001101001",
			1419 => "0000000100000000001101110100000100",
			1420 => "11111110011010010001011001101001",
			1421 => "0000000100000000000000100000001100",
			1422 => "0000001001000000000110101000000100",
			1423 => "11111111000110110001011001101001",
			1424 => "0000000001000000000110101000000100",
			1425 => "00000011001100010001011001101001",
			1426 => "00000000000000000001011001101001",
			1427 => "0000000100000000000001100100001100",
			1428 => "0000001001000000001011101000000100",
			1429 => "11111110101010100001011001101001",
			1430 => "0000001001000000001101011000000100",
			1431 => "00000001100100000001011001101001",
			1432 => "11111111010100010001011001101001",
			1433 => "11111110100101110001011001101001",
			1434 => "0000001110000000000001010100010100",
			1435 => "0000000110000000001101111100010000",
			1436 => "0000000110000000001110010100000100",
			1437 => "11111111110010000001011011100101",
			1438 => "0000000010000000001100010100001000",
			1439 => "0000000000000000000111100000000100",
			1440 => "00000001101000000001011011100101",
			1441 => "00000000000000000001011011100101",
			1442 => "00000000000000000001011011100101",
			1443 => "11111111001000100001011011100101",
			1444 => "0000000100000000000011011000001100",
			1445 => "0000000110000000001110010100001000",
			1446 => "0000000110000000001011111100000100",
			1447 => "11111110101010000001011011100101",
			1448 => "00000000010100110001011011100101",
			1449 => "11111110011001110001011011100101",
			1450 => "0000000110000000001101111100011100",
			1451 => "0000001110000000001100001000011000",
			1452 => "0000000100000000000100111000001100",
			1453 => "0000000011000000000011111100001000",
			1454 => "0000001110000000001001101000000100",
			1455 => "00000000000000000001011011100101",
			1456 => "00000000000111110001011011100101",
			1457 => "11111110101011100001011011100101",
			1458 => "0000000101000000001000000000001000",
			1459 => "0000000111000000000111111000000100",
			1460 => "00000000000000000001011011100101",
			1461 => "00000001100100100001011011100101",
			1462 => "11111111001110000001011011100101",
			1463 => "00000010010000100001011011100101",
			1464 => "11111110011110100001011011100101",
			1465 => "0000000011000000000111000000010000",
			1466 => "0000000110000000001101111100001100",
			1467 => "0000001111000000001010111000001000",
			1468 => "0000001100000000000100000000000100",
			1469 => "00000001101110010001011101111011",
			1470 => "00000000100000110001011101111011",
			1471 => "11111111111010000001011101111011",
			1472 => "11111110101011100001011101111011",
			1473 => "0000001111000000001010111000010100",
			1474 => "0000000101000000001010111100010000",
			1475 => "0000000100000000001011100100000100",
			1476 => "11111110101110110001011101111011",
			1477 => "0000000101000000001000111000000100",
			1478 => "11111111110101110001011101111011",
			1479 => "0000001111000000000000001100000100",
			1480 => "00000001011110100001011101111011",
			1481 => "00000011001100110001011101111011",
			1482 => "11111110011011110001011101111011",
			1483 => "0000000100000000000011011000001100",
			1484 => "0000000110000000001110010100001000",
			1485 => "0000000110000000001011111100000100",
			1486 => "11111110100000100001011101111011",
			1487 => "00000001011101100001011101111011",
			1488 => "11111110011001110001011101111011",
			1489 => "0000001000000000001111001000001100",
			1490 => "0000000001000000001110100000000100",
			1491 => "11111110110101000001011101111011",
			1492 => "0000001011000000000111001000000100",
			1493 => "00000100001011010001011101111011",
			1494 => "11111111001011010001011101111011",
			1495 => "0000000110000000001101111100001100",
			1496 => "0000000101000000001100101000000100",
			1497 => "11111110011100100001011101111011",
			1498 => "0000000101000000001010011100000100",
			1499 => "00000010100011100001011101111011",
			1500 => "11111110101101100001011101111011",
			1501 => "11111110011001110001011101111011",
			1502 => "00000000000000000001011101111101",
			1503 => "00000000000000000001011110000001",
			1504 => "00000000000000000001011110000101",
			1505 => "00000000000000000001011110001001",
			1506 => "00000000000000000001011110001101",
			1507 => "00000000000000000001011110010001",
			1508 => "00000000000000000001011110010101",
			1509 => "00000000000000000001011110011001",
			1510 => "00000000000000000001011110011101",
			1511 => "00000000000000000001011110100001",
			1512 => "00000000000000000001011110100101",
			1513 => "00000000000000000001011110101001",
			1514 => "00000000000000000001011110101101",
			1515 => "00000000000000000001011110110001",
			1516 => "00000000000000000001011110110101",
			1517 => "00000000000000000001011110111001",
			1518 => "00000000000000000001011110111101",
			1519 => "00000000000000000001011111000001",
			1520 => "00000000000000000001011111000101",
			1521 => "00000000000000000001011111001001",
			1522 => "00000000000000000001011111001101",
			1523 => "00000000000000000001011111010001",
			1524 => "00000000000000000001011111010101",
			1525 => "00000000000000000001011111011001",
			1526 => "00000000000000000001011111011101",
			1527 => "00000000000000000001011111100001",
			1528 => "00000000000000000001011111100101",
			1529 => "00000000000000000001011111101001",
			1530 => "00000000000000000001011111101101",
			1531 => "0000000010000000000111100000000100",
			1532 => "00000000000000000001011111111001",
			1533 => "11111111111101100001011111111001",
			1534 => "0000001110000000001010110000000100",
			1535 => "00000000000000000001100000000101",
			1536 => "11111111110101110001100000000101",
			1537 => "0000000010000000001100100100000100",
			1538 => "00000000000000000001100000010001",
			1539 => "11111111111001100001100000010001",
			1540 => "0000000010000000001100100100000100",
			1541 => "00000000000000000001100000011101",
			1542 => "11111111111110010001100000011101",
			1543 => "0000000110000000001101111100001000",
			1544 => "0000000110000000000111101000000100",
			1545 => "00000000000000000001100000110001",
			1546 => "00000000000100110001100000110001",
			1547 => "11111111111001100001100000110001",
			1548 => "0000000001000000000000011000000100",
			1549 => "00000000000000000001100001000101",
			1550 => "0000001101000000001001110100000100",
			1551 => "11111111100010000001100001000101",
			1552 => "00000000000000000001100001000101",
			1553 => "0000000110000000001101111100001000",
			1554 => "0000000110000000001011111100000100",
			1555 => "00000000000000000001100001011001",
			1556 => "00000000000101100001100001011001",
			1557 => "00000000000000000001100001011001",
			1558 => "0000000100000000001011100100001000",
			1559 => "0000000011000000000100011000000100",
			1560 => "11111111110001010001100001101101",
			1561 => "00000000000000000001100001101101",
			1562 => "00000000000000000001100001101101",
			1563 => "0000000110000000001101111100001000",
			1564 => "0000000110000000001011111100000100",
			1565 => "00000000000000000001100010000001",
			1566 => "00000000000011110001100010000001",
			1567 => "00000000000000000001100010000001",
			1568 => "0000000010000000001100100100000100",
			1569 => "00000000000000000001100010010101",
			1570 => "0000000011000000000111000000000100",
			1571 => "00000000000000000001100010010101",
			1572 => "11111111111001000001100010010101",
			1573 => "0000000110000000001101111100001000",
			1574 => "0000000110000000001011111100000100",
			1575 => "00000000000000000001100010101001",
			1576 => "00000000000011110001100010101001",
			1577 => "00000000000000000001100010101001",
			1578 => "0000000110000000001101111100001000",
			1579 => "0000000110000000001011111100000100",
			1580 => "00000000000000000001100010111101",
			1581 => "00000000001000100001100010111101",
			1582 => "00000000000000000001100010111101",
			1583 => "0000000110000000001101111100001000",
			1584 => "0000000110000000001011111100000100",
			1585 => "00000000000000000001100011010001",
			1586 => "00000000000011110001100011010001",
			1587 => "00000000000000000001100011010001",
			1588 => "0000000110000000001101111100001000",
			1589 => "0000000110000000001011111100000100",
			1590 => "00000000000000000001100011100101",
			1591 => "00000000000111010001100011100101",
			1592 => "00000000000000000001100011100101",
			1593 => "0000000010000000000111100000001000",
			1594 => "0000000010000000000000110100000100",
			1595 => "00000000000000000001100100000001",
			1596 => "00000000000011010001100100000001",
			1597 => "0000000010000000001000001100000100",
			1598 => "11111111101101010001100100000001",
			1599 => "00000000000000000001100100000001",
			1600 => "0000000100000000000101100000001100",
			1601 => "0000001111000000000011011100000100",
			1602 => "00000000000000000001100100011101",
			1603 => "0000000101000000000110100100000100",
			1604 => "11111111001111000001100100011101",
			1605 => "00000000000000000001100100011101",
			1606 => "00000000000000000001100100011101",
			1607 => "0000000110000000001101111100001100",
			1608 => "0000000110000000001011111100000100",
			1609 => "00000000000000000001100100111001",
			1610 => "0000000110000000001101111100000100",
			1611 => "00000000001001110001100100111001",
			1612 => "00000000000000000001100100111001",
			1613 => "11111111111000100001100100111001",
			1614 => "0000000010000000000111100000001100",
			1615 => "0000000110000000001011111100000100",
			1616 => "00000000000000000001100101011101",
			1617 => "0000000110000000001101111100000100",
			1618 => "00000000001000100001100101011101",
			1619 => "00000000000000000001100101011101",
			1620 => "0000000010000000001000001100000100",
			1621 => "11111111101111100001100101011101",
			1622 => "00000000000000000001100101011101",
			1623 => "0000000100000000000101100000010000",
			1624 => "0000000010000000000111010000000100",
			1625 => "00000000000000000001100110000001",
			1626 => "0000001011000000000000001100001000",
			1627 => "0000000001000000001110011100000100",
			1628 => "00000000000000000001100110000001",
			1629 => "11111111001101010001100110000001",
			1630 => "00000000000000000001100110000001",
			1631 => "00000000000000000001100110000001",
			1632 => "0000000100000000000011011000000100",
			1633 => "11111111101001000001100110100101",
			1634 => "0000000111000000000110000100001100",
			1635 => "0000000110000000001101111100001000",
			1636 => "0000000110000000001110010100000100",
			1637 => "00000000000000000001100110100101",
			1638 => "00000000001100100001100110100101",
			1639 => "00000000000000000001100110100101",
			1640 => "00000000000000000001100110100101",
			1641 => "0000000110000000001101111100010000",
			1642 => "0000000100000000001111101000000100",
			1643 => "00000000000000000001100111010001",
			1644 => "0000000110000000001011111100000100",
			1645 => "00000000000000000001100111010001",
			1646 => "0000001000000000000100010100000100",
			1647 => "00000000001011110001100111010001",
			1648 => "00000000000000000001100111010001",
			1649 => "0000000100000000001010010000000100",
			1650 => "11111111101010010001100111010001",
			1651 => "00000000000000000001100111010001",
			1652 => "0000001101000000001001110100001000",
			1653 => "0000000011000000000001110100000100",
			1654 => "00000000000000000001100111111101",
			1655 => "11111111101111110001100111111101",
			1656 => "0000000110000000001101111100001100",
			1657 => "0000000011000000000100011000000100",
			1658 => "00000000000000000001100111111101",
			1659 => "0000000110000000001011111100000100",
			1660 => "00000000000000000001100111111101",
			1661 => "00000000011011010001100111111101",
			1662 => "00000000000000000001100111111101",
			1663 => "0000000100000000000011011000001100",
			1664 => "0000001000000000000110011000001000",
			1665 => "0000000100000000001000100000000100",
			1666 => "11111110110101000001101000110001",
			1667 => "00000010011010010001101000110001",
			1668 => "11111110011011000001101000110001",
			1669 => "0000000110000000001101111100001100",
			1670 => "0000000111000000001110001100001000",
			1671 => "0000000110000000001110010100000100",
			1672 => "11111111111010000001101000110001",
			1673 => "00000001011101110001101000110001",
			1674 => "11111111001101000001101000110001",
			1675 => "11111110100111100001101000110001",
			1676 => "0000000100000000000011011000001000",
			1677 => "0000000110000000001110010100000100",
			1678 => "00000000000000000001101001100101",
			1679 => "11111110110100100001101001100101",
			1680 => "0000000110000000001101111100010000",
			1681 => "0000001100000000001100110000001100",
			1682 => "0000000110000000000111101000000100",
			1683 => "00000000000000000001101001100101",
			1684 => "0000001000000000001011000100000100",
			1685 => "00000000110001110001101001100101",
			1686 => "00000000000000000001101001100101",
			1687 => "00000000000000000001101001100101",
			1688 => "00000000000000000001101001100101",
			1689 => "0000000100000000000011011000000100",
			1690 => "11111110011110100001101010010001",
			1691 => "0000000110000000001101111100010000",
			1692 => "0000000111000000001110001100001100",
			1693 => "0000000110000000001110010100000100",
			1694 => "00000000000000000001101010010001",
			1695 => "0000000010000000001110110100000100",
			1696 => "00000001001010010001101010010001",
			1697 => "00000000000000000001101010010001",
			1698 => "11111111111010110001101010010001",
			1699 => "11111111000001010001101010010001",
			1700 => "0000000100000000000011011000000100",
			1701 => "11111110111001110001101010111101",
			1702 => "0000001100000000000011011100010000",
			1703 => "0000000110000000001101111100001100",
			1704 => "0000000110000000000111101000000100",
			1705 => "00000000000000000001101010111101",
			1706 => "0000001000000000001011000100000100",
			1707 => "00000000100100110001101010111101",
			1708 => "00000000000000000001101010111101",
			1709 => "00000000000000000001101010111101",
			1710 => "00000000000000000001101010111101",
			1711 => "0000000011000000001010101100001000",
			1712 => "0000000110000000001101111100000100",
			1713 => "11101100101000110001101011111001",
			1714 => "11010011001100010001101011111001",
			1715 => "0000000011000000000111000000001000",
			1716 => "0000000000000000000011100000000100",
			1717 => "11100101111111100001101011111001",
			1718 => "11010010111000010001101011111001",
			1719 => "0000001111000000000001111100001100",
			1720 => "0000001011000000000000101000001000",
			1721 => "0000000001000000001100100000000100",
			1722 => "11101011101110010001101011111001",
			1723 => "11010011000000010001101011111001",
			1724 => "11010010110101000001101011111001",
			1725 => "11010010110101010001101011111001",
			1726 => "0000000100000000000011011000001000",
			1727 => "0000000110000000001110010100000100",
			1728 => "00000000000000000001101100111101",
			1729 => "11111110110010110001101100111101",
			1730 => "0000000010000000000111100000010000",
			1731 => "0000000110000000001101111100001100",
			1732 => "0000000000000000000001001000001000",
			1733 => "0000000110000000000111101000000100",
			1734 => "00000000000000000001101100111101",
			1735 => "00000000110011100001101100111101",
			1736 => "00000000000000000001101100111101",
			1737 => "00000000000000000001101100111101",
			1738 => "0000001000000000000110001000000100",
			1739 => "00000000000000000001101100111101",
			1740 => "0000000011000000000111000000000100",
			1741 => "00000000000000000001101100111101",
			1742 => "11111111101001110001101100111101",
			1743 => "0000000001000000000000011000010100",
			1744 => "0000000101000000001010111000010000",
			1745 => "0000000110000000001101111100001100",
			1746 => "0000000110000000001110010100000100",
			1747 => "11111111100010110001101110001001",
			1748 => "0000000010000000000011001000000100",
			1749 => "00000001101001110001101110001001",
			1750 => "00000000000000000001101110001001",
			1751 => "11111111010011110001101110001001",
			1752 => "11111110101011100001101110001001",
			1753 => "0000001000000000000110011000001000",
			1754 => "0000000100000000001000100000000100",
			1755 => "11111110101100100001101110001001",
			1756 => "00000011110001000001101110001001",
			1757 => "0000000100000000000011011000000100",
			1758 => "11111110011010100001101110001001",
			1759 => "0000000100000000000001101100000100",
			1760 => "00000000001101010001101110001001",
			1761 => "11111110111001100001101110001001",
			1762 => "0000000100000000000011011000001100",
			1763 => "0000001000000000000110011000001000",
			1764 => "0000000100000000001111100100000100",
			1765 => "00000000000000000001101111010101",
			1766 => "00000000101010110001101111010101",
			1767 => "11111110101110110001101111010101",
			1768 => "0000001110000000000111111000010000",
			1769 => "0000001111000000001010111000001100",
			1770 => "0000000101000000001110110000001000",
			1771 => "0000000001000000001100100000000100",
			1772 => "00000000100110000001101111010101",
			1773 => "00000000000000000001101111010101",
			1774 => "00000000000000000001101111010101",
			1775 => "11111111100100100001101111010101",
			1776 => "0000000010000000001110110100001000",
			1777 => "0000001000000000001000101100000100",
			1778 => "00000001000101110001101111010101",
			1779 => "00000000000000000001101111010101",
			1780 => "00000000000000000001101111010101",
			1781 => "0000000110000000001101111100011100",
			1782 => "0000001101000000001010111100010000",
			1783 => "0000001111000000001010111000001100",
			1784 => "0000001010000000000110011100000100",
			1785 => "00000000000000000001110000010001",
			1786 => "0000000110000000000111101000000100",
			1787 => "00000000000000000001110000010001",
			1788 => "00000000101011000001110000010001",
			1789 => "11111111000000100001110000010001",
			1790 => "0000000100000000001111101000000100",
			1791 => "00000000000000000001110000010001",
			1792 => "0000000100000000000101001100000100",
			1793 => "00000001001111110001110000010001",
			1794 => "00000000000000000001110000010001",
			1795 => "11111110110101110001110000010001",
			1796 => "0000000110000000001101111100011100",
			1797 => "0000001101000000001010111100010000",
			1798 => "0000001111000000001010111000001100",
			1799 => "0000001001000000000110000000001000",
			1800 => "0000000110000000001110010100000100",
			1801 => "00000000000000000001110001001101",
			1802 => "00000000010000000001110001001101",
			1803 => "00000000000000000001110001001101",
			1804 => "11111111011010110001110001001101",
			1805 => "0000001001000000001110100000000100",
			1806 => "00000000000000000001110001001101",
			1807 => "0000000100000000001111101000000100",
			1808 => "00000000000000000001110001001101",
			1809 => "00000000111111110001110001001101",
			1810 => "11111111010000110001110001001101",
			1811 => "0000000100000000000011011000001100",
			1812 => "0000001000000000000110011000001000",
			1813 => "0000000000000000001001101000000100",
			1814 => "11111111001101010001110010100001",
			1815 => "00000001001011010001110010100001",
			1816 => "11111110011101100001110010100001",
			1817 => "0000000010000000000111100000010000",
			1818 => "0000000100000000001011100100001000",
			1819 => "0000000000000000000100000000000100",
			1820 => "00000000011101100001110010100001",
			1821 => "11111111101011100001110010100001",
			1822 => "0000000000000000000001001000000100",
			1823 => "00000001010111000001110010100001",
			1824 => "00000000000000000001110010100001",
			1825 => "0000000000000000000011010000001000",
			1826 => "0000001101000000001011011100000100",
			1827 => "00000000000000000001110010100001",
			1828 => "00000000100100100001110010100001",
			1829 => "0000000011000000000111000000000100",
			1830 => "00000000000000000001110010100001",
			1831 => "11111111000100100001110010100001",
			1832 => "0000000110000000000001111000100000",
			1833 => "0000000011000000000111000000001100",
			1834 => "0000000110000000000111101000000100",
			1835 => "00000000000000000001110011111101",
			1836 => "0000000000000000000100000100000100",
			1837 => "00000000011110110001110011111101",
			1838 => "00000000000000000001110011111101",
			1839 => "0000000011000000000100011000001100",
			1840 => "0000001111000000000101101100000100",
			1841 => "00000000000000000001110011111101",
			1842 => "0000000001000000001110011100000100",
			1843 => "00000000000000000001110011111101",
			1844 => "11111111010101100001110011111101",
			1845 => "0000000000000000001011010100000100",
			1846 => "00000000000000000001110011111101",
			1847 => "00000000100100010001110011111101",
			1848 => "0000001101000000001011011100001000",
			1849 => "0000000011000000000111000100000100",
			1850 => "00000000000000000001110011111101",
			1851 => "11111110101110110001110011111101",
			1852 => "0000000101000000000100000100000100",
			1853 => "00000000000000000001110011111101",
			1854 => "11111111101111010001110011111101",
			1855 => "0000000100000000000011011000001100",
			1856 => "0000001000000000000110011000001000",
			1857 => "0000000100000000001000100000000100",
			1858 => "11111111010011000001110101001001",
			1859 => "00000001001011000001110101001001",
			1860 => "11111110011101000001110101001001",
			1861 => "0000001100000000000011011100011000",
			1862 => "0000000100000000001011100100001100",
			1863 => "0000000111000000001101100000001000",
			1864 => "0000000001000000001100100000000100",
			1865 => "00000000000000000001110101001001",
			1866 => "11111111000000110001110101001001",
			1867 => "00000001001001100001110101001001",
			1868 => "0000000010000000000011001000001000",
			1869 => "0000001010000000000110011100000100",
			1870 => "00000000000000000001110101001001",
			1871 => "00000001010010110001110101001001",
			1872 => "00000000000000000001110101001001",
			1873 => "11111111000100100001110101001001",
			1874 => "0000000110000000001101111100011100",
			1875 => "0000000011000000000100011000010100",
			1876 => "0000000001000000000000011000010000",
			1877 => "0000000101000000000011100000001100",
			1878 => "0000000110000000001110010100000100",
			1879 => "00000000000000000001110110000101",
			1880 => "0000000010000000000011001000000100",
			1881 => "00000001000000000001110110000101",
			1882 => "00000000000000000001110110000101",
			1883 => "00000000000000000001110110000101",
			1884 => "11111110110100110001110110000101",
			1885 => "0000000100000000001111101000000100",
			1886 => "00000000000000000001110110000101",
			1887 => "00000001010101110001110110000101",
			1888 => "11111110100111010001110110000101",
			1889 => "0000000110000000001101111100100000",
			1890 => "0000001101000000001010111100010000",
			1891 => "0000001001000000000110000000001100",
			1892 => "0000000010000000000011001000001000",
			1893 => "0000001010000000000110011100000100",
			1894 => "00000000000000000001110111001001",
			1895 => "00000000001010010001110111001001",
			1896 => "00000000000000000001110111001001",
			1897 => "11111111100101010001110111001001",
			1898 => "0000000100000000001011110000000100",
			1899 => "00000000000000000001110111001001",
			1900 => "0000001001000000001110100000000100",
			1901 => "00000000000000000001110111001001",
			1902 => "0000000110000000000001111000000100",
			1903 => "00000000000000000001110111001001",
			1904 => "00000000100111010001110111001001",
			1905 => "11111111010111100001110111001001",
			1906 => "0000000110000000001101111100100000",
			1907 => "0000001101000000001010111100010100",
			1908 => "0000001111000000001010111000010000",
			1909 => "0000001010000000000110011100000100",
			1910 => "00000000000000000001111000001101",
			1911 => "0000000110000000001101111100001000",
			1912 => "0000000110000000000111101000000100",
			1913 => "00000000000000000001111000001101",
			1914 => "00000000010100010001111000001101",
			1915 => "00000000000000000001111000001101",
			1916 => "11111111001111000001111000001101",
			1917 => "0000001001000000001110100000000100",
			1918 => "00000000000000000001111000001101",
			1919 => "0000000100000000001111101000000100",
			1920 => "00000000000000000001111000001101",
			1921 => "00000001010010110001111000001101",
			1922 => "11111111000010110001111000001101",
			1923 => "0000000110000000001101111100100000",
			1924 => "0000000011000000000100011000010100",
			1925 => "0000000001000000000000011000010000",
			1926 => "0000000101000000000100011000001100",
			1927 => "0000000010000000000011001000001000",
			1928 => "0000001010000000000110011100000100",
			1929 => "00000000000000000001111001010001",
			1930 => "00000000011101000001111001010001",
			1931 => "00000000000000000001111001010001",
			1932 => "00000000000000000001111001010001",
			1933 => "11111111011101000001111001010001",
			1934 => "0000000000000000001011010100000100",
			1935 => "00000000000000000001111001010001",
			1936 => "0000001101000000001001001000000100",
			1937 => "00000000000000000001111001010001",
			1938 => "00000000101110110001111001010001",
			1939 => "11111111011000110001111001010001",
			1940 => "0000001110000000000001010100001100",
			1941 => "0000001010000000001000101100001000",
			1942 => "0000001111000000001010111100000100",
			1943 => "00000010000100110001111010101101",
			1944 => "11111110011111110001111010101101",
			1945 => "11111110011101000001111010101101",
			1946 => "0000001111000000001101010100010000",
			1947 => "0000001100000000001100001000001100",
			1948 => "0000000100000000001010101000000100",
			1949 => "11111110011000010001111010101101",
			1950 => "0000000111000000000100010100000100",
			1951 => "00000010000000000001111010101101",
			1952 => "00000011010000110001111010101101",
			1953 => "11111110011001100001111010101101",
			1954 => "0000000100000000000011011000000100",
			1955 => "11111110010111100001111010101101",
			1956 => "0000000110000000001101111100001100",
			1957 => "0000000110000000000001111000000100",
			1958 => "11111110011011110001111010101101",
			1959 => "0000000100000000001111011000000100",
			1960 => "00000011011101010001111010101101",
			1961 => "11111110100001100001111010101101",
			1962 => "11111110011000000001111010101101",
			1963 => "0000001110000000000001010100011000",
			1964 => "0000000110000000001101111100010000",
			1965 => "0000001111000000001010111000001100",
			1966 => "0000000110000000000111101000000100",
			1967 => "00000000000000000001111100001001",
			1968 => "0000001000000000001011000100000100",
			1969 => "00000001100110000001111100001001",
			1970 => "00000000000000000001111100001001",
			1971 => "11111111111011010001111100001001",
			1972 => "0000000110000000001101111100000100",
			1973 => "00000000000000000001111100001001",
			1974 => "11111111011010100001111100001001",
			1975 => "0000000100000000000011011000000100",
			1976 => "11111110011010010001111100001001",
			1977 => "0000000110000000001101111100010000",
			1978 => "0000001110000000001100001000001100",
			1979 => "0000001111000000001101010100001000",
			1980 => "0000000100000000001101100100000100",
			1981 => "00000000111001010001111100001001",
			1982 => "00000000000000000001111100001001",
			1983 => "11111110110010000001111100001001",
			1984 => "00000001101101100001111100001001",
			1985 => "11111110100011010001111100001001",
			1986 => "0000000100000000000011011000001100",
			1987 => "0000001000000000000110011000001000",
			1988 => "0000000000000000001011010100000100",
			1989 => "11111110110110110001111101010101",
			1990 => "00000010010001110001111101010101",
			1991 => "11111110011011000001111101010101",
			1992 => "0000000110000000001101111100011000",
			1993 => "0000000111000000001110001100010100",
			1994 => "0000000110000000001110010100000100",
			1995 => "00000000000000000001111101010101",
			1996 => "0000000001000000000000011000001000",
			1997 => "0000000010000000000011001000000100",
			1998 => "00000001100110010001111101010101",
			1999 => "00000000000000000001111101010101",
			2000 => "0000000001000000000110000000000100",
			2001 => "11111111101011110001111101010101",
			2002 => "00000000111111010001111101010101",
			2003 => "11111111010000110001111101010101",
			2004 => "11111110101001100001111101010101",
			2005 => "0000000110000000001101111100100100",
			2006 => "0000000011000000000100011000011000",
			2007 => "0000000100000000001101000000001000",
			2008 => "0000001001000000000000011000000100",
			2009 => "00000000000000000001111110100001",
			2010 => "11111110101111100001111110100001",
			2011 => "0000000101000000000100011000001100",
			2012 => "0000000110000000000111101000000100",
			2013 => "00000000000000000001111110100001",
			2014 => "0000000000000000000100000100000100",
			2015 => "00000001000001010001111110100001",
			2016 => "00000000000000000001111110100001",
			2017 => "00000000000000000001111110100001",
			2018 => "0000000100000000001111101000000100",
			2019 => "00000000000000000001111110100001",
			2020 => "0000001101000000001011000000000100",
			2021 => "00000000000000000001111110100001",
			2022 => "00000001011111110001111110100001",
			2023 => "11111110100100110001111110100001",
			2024 => "0000000011000000000111000000010000",
			2025 => "0000000100000000001011011000000100",
			2026 => "11111111011010100001111111111101",
			2027 => "0000001010000000000010101000001000",
			2028 => "0000000110000000000111101000000100",
			2029 => "00000000000000000001111111111101",
			2030 => "00000001100100000001111111111101",
			2031 => "00000000000000000001111111111101",
			2032 => "0000001010000000001010100100001000",
			2033 => "0000000100000000001111101000000100",
			2034 => "11111110101111010001111111111101",
			2035 => "00000011010100000001111111111101",
			2036 => "0000000100000000000011011000000100",
			2037 => "11111110011010110001111111111101",
			2038 => "0000000110000000001101111100010000",
			2039 => "0000001110000000000111111000001100",
			2040 => "0000001111000000000111001000001000",
			2041 => "0000000010000000001100100100000100",
			2042 => "00000000111111100001111111111101",
			2043 => "00000000000000000001111111111101",
			2044 => "11111110110001010001111111111101",
			2045 => "00000001110001010001111111111101",
			2046 => "11111110100101100001111111111101",
			2047 => "0000000100000000000011011000010000",
			2048 => "0000000110000000001110010100001100",
			2049 => "0000000010000000001110101000000100",
			2050 => "00000000000000000010000001011001",
			2051 => "0000000011000000000001111100000100",
			2052 => "00000000000000000010000001011001",
			2053 => "00000000011000000010000001011001",
			2054 => "11111110100001010010000001011001",
			2055 => "0000000110000000001101111100011100",
			2056 => "0000000111000000001110001100011000",
			2057 => "0000000100000000000000101100001100",
			2058 => "0000001010000000001001000100001000",
			2059 => "0000001010000000001000010100000100",
			2060 => "00000000000000000010000001011001",
			2061 => "00000000100001110010000001011001",
			2062 => "11111111101001110010000001011001",
			2063 => "0000000110000000001110010100000100",
			2064 => "00000000000000000010000001011001",
			2065 => "0000000010000000001110110100000100",
			2066 => "00000001001000000010000001011001",
			2067 => "00000000000000000010000001011001",
			2068 => "00000000000000000010000001011001",
			2069 => "11111111001100110010000001011001",
			2070 => "0000001110000000000101000100010000",
			2071 => "0000001111000000001010111000001100",
			2072 => "0000000110000000001101111100001000",
			2073 => "0000000011000000000111000000000100",
			2074 => "00000001100111100010000011000101",
			2075 => "00000000000000000010000011000101",
			2076 => "00000000000000000010000011000101",
			2077 => "11111111111001110010000011000101",
			2078 => "0000000100000000000011011000001100",
			2079 => "0000000110000000001110010100001000",
			2080 => "0000000110000000001011111100000100",
			2081 => "11111110101100010010000011000101",
			2082 => "00000000010100100010000011000101",
			2083 => "11111110011010000010000011000101",
			2084 => "0000000110000000001101111100011000",
			2085 => "0000001110000000001100001000010100",
			2086 => "0000001111000000000111001000001000",
			2087 => "0000000000000000001000011000000100",
			2088 => "00000001011010110010000011000101",
			2089 => "11111111110110100010000011000101",
			2090 => "0000000100000000001010010000000100",
			2091 => "11111110101011100010000011000101",
			2092 => "0000000010000000001100010100000100",
			2093 => "00000000100110110010000011000101",
			2094 => "11111111110001110010000011000101",
			2095 => "00000010000111000010000011000101",
			2096 => "11111110011111000010000011000101",
			2097 => "0000000011000000000111000000010000",
			2098 => "0000000110000000001101111100001000",
			2099 => "0000000110000000000111101000000100",
			2100 => "00000000000000000010000101000001",
			2101 => "00000001101000000010000101000001",
			2102 => "0000000011000000001010101100000100",
			2103 => "00000000000000000010000101000001",
			2104 => "11111111000111010010000101000001",
			2105 => "0000000100000000000011011000001100",
			2106 => "0000001000000000000110011000001000",
			2107 => "0000000000000000001001101000000100",
			2108 => "11111110100000110010000101000001",
			2109 => "00000011000001000010000101000001",
			2110 => "11111110011001110010000101000001",
			2111 => "0000001000000000001111001000010000",
			2112 => "0000000010000000001110110100001100",
			2113 => "0000001111000000001011011100000100",
			2114 => "00000000000000000010000101000001",
			2115 => "0000000101000000001000111100000100",
			2116 => "00000000000000000010000101000001",
			2117 => "00000010100000100010000101000001",
			2118 => "11111111110101110010000101000001",
			2119 => "0000000110000000001101111100010000",
			2120 => "0000001000000000001000110000000100",
			2121 => "11111110101100110010000101000001",
			2122 => "0000000010000000001001011100001000",
			2123 => "0000000000000000001001001000000100",
			2124 => "00000001010011000010000101000001",
			2125 => "00000000000000000010000101000001",
			2126 => "11111111010001000010000101000001",
			2127 => "11111110011100110010000101000001",
			2128 => "0000001110000000000001110000010000",
			2129 => "0000000110000000001101111100001100",
			2130 => "0000001111000000001010111100001000",
			2131 => "0000000000000000000001000000000100",
			2132 => "00000001110000100010000111000101",
			2133 => "11111111001000110010000111000101",
			2134 => "11111110101010000010000111000101",
			2135 => "11111110100000010010000111000101",
			2136 => "0000001111000000001010111000001100",
			2137 => "0000000101000000001010111100001000",
			2138 => "0000000100000000001011100100000100",
			2139 => "11111110100110110010000111000101",
			2140 => "00000010110101100010000111000101",
			2141 => "11111110011011100010000111000101",
			2142 => "0000000100000000000011011000001100",
			2143 => "0000000110000000001110010100001000",
			2144 => "0000000110000000001011111100000100",
			2145 => "11111110011111010010000111000101",
			2146 => "00000001100110010010000111000101",
			2147 => "11111110011001100010000111000101",
			2148 => "0000001000000000001111001000001100",
			2149 => "0000000101000000000110100100000100",
			2150 => "11111110110000110010000111000101",
			2151 => "0000001011000000000111001000000100",
			2152 => "00000101010001110010000111000101",
			2153 => "11111111000110110010000111000101",
			2154 => "0000000110000000001101111100001100",
			2155 => "0000000101000000001100101000000100",
			2156 => "11111110011011110010000111000101",
			2157 => "0000000101000000001010011100000100",
			2158 => "00000011000100000010000111000101",
			2159 => "11111110101010100010000111000101",
			2160 => "11111110011001100010000111000101",
			2161 => "0000000011000000000111000000010100",
			2162 => "0000000100000000001011011000000100",
			2163 => "11111111110000000010001001010001",
			2164 => "0000001010000000000010101000001100",
			2165 => "0000001100000000000000101000001000",
			2166 => "0000001111000000000111001000000100",
			2167 => "00000001101001110010001001010001",
			2168 => "00000000000000000010001001010001",
			2169 => "00000010111100000010001001010001",
			2170 => "11111111010011010010001001010001",
			2171 => "0000000100000000000011011000001100",
			2172 => "0000001010000000001010100100001000",
			2173 => "0000000100000000001111101000000100",
			2174 => "11111110011100100010001001010001",
			2175 => "00010000110001000010001001010001",
			2176 => "11111110011001010010001001010001",
			2177 => "0000000010000000001110000100010000",
			2178 => "0000001011000000001100001000001000",
			2179 => "0000001111000000001010111100000100",
			2180 => "00000001011010110010001001010001",
			2181 => "11111110101011010010001001010001",
			2182 => "0000001100000000000110000100000100",
			2183 => "00000011010110110010001001010001",
			2184 => "11111111010010100010001001010001",
			2185 => "0000000010000000001010001000010100",
			2186 => "0000000010000000001001011100001100",
			2187 => "0000000010000000000101001000001000",
			2188 => "0000001100000000000111111000000100",
			2189 => "11111111101101000010001001010001",
			2190 => "00000000000110110010001001010001",
			2191 => "11111110011110010010001001010001",
			2192 => "0000001010000000001100000100000100",
			2193 => "00000010010010100010001001010001",
			2194 => "00000000000000000010001001010001",
			2195 => "11111110011010110010001001010001",
			2196 => "0000001110000000000001010100010000",
			2197 => "0000000110000000001101111100001100",
			2198 => "0000001111000000001010111100001000",
			2199 => "0000000000000000000111100000000100",
			2200 => "00000001111001110010001011011101",
			2201 => "11111110111111100010001011011101",
			2202 => "11111110100010100010001011011101",
			2203 => "11111110011101010010001011011101",
			2204 => "0000001111000000001010111000010000",
			2205 => "0000000111000000000000101000001100",
			2206 => "0000000001000000001100100000001000",
			2207 => "0000001111000000000000001100000100",
			2208 => "00000001110100110010001011011101",
			2209 => "00000011111100010010001011011101",
			2210 => "11111110011001100010001011011101",
			2211 => "11111110011010000010001011011101",
			2212 => "0000000100000000000011011000001100",
			2213 => "0000000110000000001110010100001000",
			2214 => "0000000110000000001011111100000100",
			2215 => "11111110011100110010001011011101",
			2216 => "00000010010011110010001011011101",
			2217 => "11111110011000000010001011011101",
			2218 => "0000000010000000000111100000001000",
			2219 => "0000000110000000001101111100000100",
			2220 => "00000010000000000010001011011101",
			2221 => "11111111011011010010001011011101",
			2222 => "0000000010000000001110110100010000",
			2223 => "0000000010000000001110110100001000",
			2224 => "0000000100000000001010010000000100",
			2225 => "11111110011010100010001011011101",
			2226 => "11111111101010110010001011011101",
			2227 => "0000000100000000000001001100000100",
			2228 => "00000110010110100010001011011101",
			2229 => "11111110111001010010001011011101",
			2230 => "11111110011000110010001011011101",
			2231 => "0000000011000000001000101100010100",
			2232 => "0000000110000000001101111100010000",
			2233 => "0000000110000000001110010100000100",
			2234 => "11111110010101100010001101111011",
			2235 => "0000000000000000000101001000001000",
			2236 => "0000001111000000000001111100000100",
			2237 => "00000001111110110010001101111011",
			2238 => "00000000001100100010001101111011",
			2239 => "11111111000000000010001101111011",
			2240 => "11111110011100100010001101111011",
			2241 => "0000001111000000001010111000010000",
			2242 => "0000001101000000001100101100001100",
			2243 => "0000000001000000001100100000001000",
			2244 => "0000001111000000000001111100000100",
			2245 => "00000001111000110010001101111011",
			2246 => "00000111000001110010001101111011",
			2247 => "11111110100100110010001101111011",
			2248 => "11111110011001100010001101111011",
			2249 => "0000000100000000000011011000001100",
			2250 => "0000000110000000001110010100001000",
			2251 => "0000000110000000001011111100000100",
			2252 => "11111110011011110010001101111011",
			2253 => "00000010111010100010001101111011",
			2254 => "11111110010111110010001101111011",
			2255 => "0000000010000000000111100000001000",
			2256 => "0000000110000000001101111100000100",
			2257 => "00000010011011010010001101111011",
			2258 => "11111111010110100010001101111011",
			2259 => "0000000100000000000001101100001100",
			2260 => "0000000010000000001110110100000100",
			2261 => "11111110110000110010001101111011",
			2262 => "0000000110000000001011001100000100",
			2263 => "00000100101001110010001101111011",
			2264 => "11111111010101010010001101111011",
			2265 => "0000000110000000001101111100001000",
			2266 => "0000000110000000001101111100000100",
			2267 => "11111110011010000010001101111011",
			2268 => "00000001011011100010001101111011",
			2269 => "11111110011000100010001101111011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(736, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(1502, initial_addr_3'length));
	end generate gen_rom_6;

	gen_rom_7: if SELECT_ROM = 7 generate
		bank <= (
			0 => "0000000100000000000110110001101000",
			1 => "0000001001000000001100011000111000",
			2 => "0000001111000000001110110100101000",
			3 => "0000000100000000001010000100001000",
			4 => "0000000111000000000100010100000100",
			5 => "00000000000000000000000100010101",
			6 => "11111110000011110000000100010101",
			7 => "0000001001000000000110101000010000",
			8 => "0000001100000000000100010100001000",
			9 => "0000001001000000000010001100000100",
			10 => "11111111101101010000000100010101",
			11 => "00000000001001110000000100010101",
			12 => "0000001110000000000100010100000100",
			13 => "11111111110111000000000100010101",
			14 => "11111110011110000000000100010101",
			15 => "0000000001000000001110100000001000",
			16 => "0000001110000000001100110000000100",
			17 => "00000001110101000000000100010101",
			18 => "11111111011110110000000100010101",
			19 => "0000000110000000000111101000000100",
			20 => "00000001001110100000000100010101",
			21 => "00000000001001010000000100010101",
			22 => "0000000101000000001000011000001000",
			23 => "0000001001000000001011111100000100",
			24 => "00000010000000100000000100010101",
			25 => "11111110010010000000000100010101",
			26 => "0000000010000000000101010100000100",
			27 => "00000010010100110000000100010101",
			28 => "11111111001011010000000100010101",
			29 => "0000000110000000001001111100011100",
			30 => "0000001010000000000001010000000100",
			31 => "11111110011001000000000100010101",
			32 => "0000001100000000000100011000001100",
			33 => "0000000010000000000110001100001000",
			34 => "0000000110000000000100111100000100",
			35 => "11111111101110010000000100010101",
			36 => "11111110010010100000000100010101",
			37 => "00000000000000000000000100010101",
			38 => "0000001111000000000101000000001000",
			39 => "0000000100000000001011100000000100",
			40 => "00000001001010010000000100010101",
			41 => "11111111001111100000000100010101",
			42 => "11111110011100000000000100010101",
			43 => "0000001110000000000010110000001100",
			44 => "0000000100000000001110111000000100",
			45 => "11111111000101000000000100010101",
			46 => "0000001100000000001000000000000100",
			47 => "00000000101010100000000100010101",
			48 => "00000010000000100000000100010101",
			49 => "0000001100000000000001011000000100",
			50 => "11111110100001100000000100010101",
			51 => "00000000110100100000000100010101",
			52 => "0000000110000000001011001100001100",
			53 => "0000000100000000000011111000000100",
			54 => "11111101110000110000000100010101",
			55 => "0000000100000000001110011000000100",
			56 => "00000000000000000000000100010101",
			57 => "11111110011011110000000100010101",
			58 => "0000000010000000000010000100001000",
			59 => "0000000001000000001110011100000100",
			60 => "11111111110011010000000100010101",
			61 => "00000001100100100000000100010101",
			62 => "0000001010000000001100000100001100",
			63 => "0000001000000000001111000100000100",
			64 => "11111110101111100000000100010101",
			65 => "0000000100000000000101100000000100",
			66 => "00000001111110010000000100010101",
			67 => "00000000000000000000000100010101",
			68 => "11111110100011110000000100010101",
			69 => "0000000111000000001100101000111100",
			70 => "0000000001000000001100100000001000",
			71 => "0000000110000000001011001100000100",
			72 => "11111110011000010000001000011001",
			73 => "11111111100101010000001000011001",
			74 => "0000000110000000000001000100000100",
			75 => "11111110011000000000001000011001",
			76 => "0000000110000000000100111100100000",
			77 => "0000001110000000000100010100010000",
			78 => "0000000101000000000101101100001000",
			79 => "0000000011000000001011000100000100",
			80 => "00000000111010100000001000011001",
			81 => "00000000010101000000001000011001",
			82 => "0000000110000000000001111000000100",
			83 => "00000001101011110000001000011001",
			84 => "00000000111000010000001000011001",
			85 => "0000001111000000001011011100001000",
			86 => "0000000110000000000111101000000100",
			87 => "00000001000011000000001000011001",
			88 => "11111111010110110000001000011001",
			89 => "0000001100000000000100000000000100",
			90 => "00000000011000110000001000011001",
			91 => "00000000111000110000001000011001",
			92 => "0000001100000000001100110000001100",
			93 => "0000001010000000001001101000001000",
			94 => "0000001011000000000111001000000100",
			95 => "11111110001111100000001000011001",
			96 => "11111111000101100000001000011001",
			97 => "00000001000011000000001000011001",
			98 => "00000001011111100000001000011001",
			99 => "0000001000000000001001101000010000",
			100 => "0000000001000000001011101000001100",
			101 => "0000000001000000001011101000000100",
			102 => "11111110011110100000001000011001",
			103 => "0000000101000000000001011000000100",
			104 => "11111110111010010000001000011001",
			105 => "00000010101010010000001000011001",
			106 => "11111110010111010000001000011001",
			107 => "0000001000000000000010011000101100",
			108 => "0000001110000000001101101100010100",
			109 => "0000001001000000000111101100010000",
			110 => "0000001111000000001100010000001000",
			111 => "0000001101000000000001011000000100",
			112 => "00000001011101000000001000011001",
			113 => "11111110010011000000001000011001",
			114 => "0000000110000000000100111100000100",
			115 => "00000011001000110000001000011001",
			116 => "00000000111011100000001000011001",
			117 => "11111110010110000000001000011001",
			118 => "0000000110000000001001111100001000",
			119 => "0000001000000000001001101000000100",
			120 => "00000000100001100000001000011001",
			121 => "11111110010011000000001000011001",
			122 => "0000001100000000000111010000001000",
			123 => "0000001010000000000110011100000100",
			124 => "11111110001110010000001000011001",
			125 => "00000000000100110000001000011001",
			126 => "0000001111000000001010110100000100",
			127 => "00000011011100000000001000011001",
			128 => "11111111111010100000001000011001",
			129 => "0000001000000000000000110000001000",
			130 => "0000001000000000000000110000000100",
			131 => "11111110011010110000001000011001",
			132 => "00000001010000000000001000011001",
			133 => "11111110010111110000001000011001",
			134 => "0000001100000000000000001101100000",
			135 => "0000000001000000000000011000010000",
			136 => "0000000010000000000001001000001000",
			137 => "0000000110000000000001111000000100",
			138 => "11111110110010110000001100111101",
			139 => "00000001111000110000001100111101",
			140 => "0000000110000000001011001100000100",
			141 => "11111110011000010000001100111101",
			142 => "00000000000000000000001100111101",
			143 => "0000000100000000000000010000010000",
			144 => "0000001110000000001000111000000100",
			145 => "11111111100000100000001100111101",
			146 => "0000001011000000001110001100000100",
			147 => "11111110000101110000001100111101",
			148 => "0000001011000000001101111000000100",
			149 => "00000000000000000000001100111101",
			150 => "11111110011011010000001100111101",
			151 => "0000001100000000000000101000100000",
			152 => "0000001100000000000100010100010000",
			153 => "0000001100000000000100010100001000",
			154 => "0000000011000000000100010100000100",
			155 => "00000000101111100000001100111101",
			156 => "00000000001010010000001100111101",
			157 => "0000000100000000000001101100000100",
			158 => "00000000111011010000001100111101",
			159 => "11111110000011100000001100111101",
			160 => "0000000100000000000100001100001000",
			161 => "0000001100000000000100010100000100",
			162 => "11111111001001000000001100111101",
			163 => "11111111111110100000001100111101",
			164 => "0000001100000000000100010100000100",
			165 => "00000000000000000000001100111101",
			166 => "00000001010010110000001100111101",
			167 => "0000001100000000000000101000010000",
			168 => "0000001010000000000001010000001000",
			169 => "0000000010000000000010000000000100",
			170 => "00000001011100010000001100111101",
			171 => "00000011101001100000001100111101",
			172 => "0000000100000000000010111000000100",
			173 => "11111110101100010000001100111101",
			174 => "00000000111100110000001100111101",
			175 => "0000001100000000000000101000001000",
			176 => "0000001111000000000101110100000100",
			177 => "00000000010111000000001100111101",
			178 => "11111101110011010000001100111101",
			179 => "0000001110000000001001110000000100",
			180 => "00000001000001000000001100111101",
			181 => "00000000010011000000001100111101",
			182 => "0000001000000000001001101000001000",
			183 => "0000001110000000000100000100000100",
			184 => "00000001010101110000001100111101",
			185 => "11111110011010100000001100111101",
			186 => "0000000100000000000110110000101000",
			187 => "0000001000000000000110001000010000",
			188 => "0000000010000000000101000000001100",
			189 => "0000000100000000001001001100001000",
			190 => "0000000100000000000010111000000100",
			191 => "11111111100101110000001100111101",
			192 => "00000011100111110000001100111101",
			193 => "11111110100010100000001100111101",
			194 => "11111110011001110000001100111101",
			195 => "0000000100000000000011101100001100",
			196 => "0000000100000000000101010100000100",
			197 => "11111111101111000000001100111101",
			198 => "0000001100000000000111001000000100",
			199 => "00000000110110110000001100111101",
			200 => "00000010010100110000001100111101",
			201 => "0000001000000000000001110100000100",
			202 => "11111110001010010000001100111101",
			203 => "0000000110000000000101010000000100",
			204 => "11111110010010100000001100111101",
			205 => "00000001000111110000001100111101",
			206 => "11111110011001000000001100111101",
			207 => "0000000111000000001101111001100100",
			208 => "0000000100000000000001100101001000",
			209 => "0000000110000000000001000100001000",
			210 => "0000000110000000000001000100000100",
			211 => "11111110010100000000010010000001",
			212 => "11111111101011000000010010000001",
			213 => "0000001110000000001000111100100000",
			214 => "0000001011000000001100001000010000",
			215 => "0000000011000000000100000000001000",
			216 => "0000000111000000000111111000000100",
			217 => "00000000100010100000010010000001",
			218 => "00000001101010110000010010000001",
			219 => "0000001111000000000010001000000100",
			220 => "00000000101100110000010010000001",
			221 => "00000001100101100000010010000001",
			222 => "0000000100000000000101010100001000",
			223 => "0000000110000000000100110100000100",
			224 => "00000001101111100000010010000001",
			225 => "00000000001111000000010010000001",
			226 => "0000001001000000000111100100000100",
			227 => "00000001110000010000010010000001",
			228 => "00000010010111010000010010000001",
			229 => "0000000100000000000010111000010000",
			230 => "0000000111000000001000111000001000",
			231 => "0000000110000000001100011000000100",
			232 => "00000000010010010000010010000001",
			233 => "11111110111101000000010010000001",
			234 => "0000001001000000000001111000000100",
			235 => "00000001001011110000010010000001",
			236 => "11111110101001000000010010000001",
			237 => "0000000110000000001011001100001000",
			238 => "0000001001000000001101101000000100",
			239 => "00000000111001100000010010000001",
			240 => "00000001101101010000010010000001",
			241 => "0000000111000000001101100000000100",
			242 => "11111111001010110000010010000001",
			243 => "00000001010100110000010010000001",
			244 => "0000000110000000000100110100001000",
			245 => "0000001101000000001100101100000100",
			246 => "11111110010010000000010010000001",
			247 => "11111111010111000000010010000001",
			248 => "0000000101000000000100001000001100",
			249 => "0000000110000000001100011000000100",
			250 => "11111111011001110000010010000001",
			251 => "0000000000000000001101111000000100",
			252 => "00000000110100100000010010000001",
			253 => "00000010011100010000010010000001",
			254 => "0000001111000000000110010000000100",
			255 => "11111110001110100000010010000001",
			256 => "00000001101010010000010010000001",
			257 => "0000001000000000001001101000001100",
			258 => "0000000111000000000001111100001000",
			259 => "0000000111000000000001111100000100",
			260 => "11111110010110010000010010000001",
			261 => "00000010000001000000010010000001",
			262 => "11111110010001110000010010000001",
			263 => "0000000100000000000010010000110000",
			264 => "0000001000000000001111001000011000",
			265 => "0000001111000000001000000100001100",
			266 => "0000000100000000000100001100001000",
			267 => "0000000100000000000011001100000100",
			268 => "11111111100111100000010010000001",
			269 => "00000100011011100000010010000001",
			270 => "11111110010110000000010010000001",
			271 => "0000001000000000001001101000000100",
			272 => "00000000000000000000010010000001",
			273 => "0000000111000000000111110000000100",
			274 => "11111110010001100000010010000001",
			275 => "11111111111010100000010010000001",
			276 => "0000001111000000000000010100010000",
			277 => "0000000100000000001001001100001000",
			278 => "0000001010000000000110011100000100",
			279 => "00000000011010000000010010000001",
			280 => "11111110001111110000010010000001",
			281 => "0000000000000000000000111000000100",
			282 => "00000101000011000000010010000001",
			283 => "00000001100111100000010010000001",
			284 => "0000000110000000000100101100000100",
			285 => "11111110000101010000010010000001",
			286 => "00000001101101100000010010000001",
			287 => "11111110010010110000010010000001",
			288 => "0000000111000000001110001101100100",
			289 => "0000000100000000000110110001000100",
			290 => "0000000110000000000001000100000100",
			291 => "11111110011000110000010111001101",
			292 => "0000000100000000000100001100100000",
			293 => "0000001010000000001010110000010000",
			294 => "0000000010000000000010000000001000",
			295 => "0000000110000000000100110100000100",
			296 => "00000000100011110000010111001101",
			297 => "00000000000111100000010111001101",
			298 => "0000000110000000001010011000000100",
			299 => "00000001111111000000010111001101",
			300 => "00000000100100010000010111001101",
			301 => "0000000010000000001100010100001000",
			302 => "0000001001000000001101101000000100",
			303 => "11111111111110000000010111001101",
			304 => "00000001100100000000010111001101",
			305 => "0000001100000000000100000000000100",
			306 => "11111111000001010000010111001101",
			307 => "00000000100101100000010111001101",
			308 => "0000001001000000001001111000010000",
			309 => "0000000011000000001000111000001000",
			310 => "0000000011000000000000111000000100",
			311 => "00000001011000110000010111001101",
			312 => "00000000010110000000010111001101",
			313 => "0000001011000000000100010100000100",
			314 => "00000001000010000000010111001101",
			315 => "11111110101001010000010111001101",
			316 => "0000000101000000001101010100001000",
			317 => "0000000011000000001001110000000100",
			318 => "00000001011011010000010111001101",
			319 => "00000000110110110000010111001101",
			320 => "0000001111000000000010000000000100",
			321 => "11111111100100010000010111001101",
			322 => "00000001110110000000010111001101",
			323 => "0000000001000000001110100000011000",
			324 => "0000001001000000001110100000010100",
			325 => "0000000001000000001100100000000100",
			326 => "11111110011000010000010111001101",
			327 => "0000000101000000001000111100001000",
			328 => "0000000100000000001110011000000100",
			329 => "11111110000101000000010111001101",
			330 => "00000000000000000000010111001101",
			331 => "0000000010000000001001011100000100",
			332 => "00000001010000100000010111001101",
			333 => "11111110111010000000010111001101",
			334 => "11111101011110100000010111001101",
			335 => "0000000100000000000001001100000100",
			336 => "00000000011000110000010111001101",
			337 => "11111110011100000000010111001101",
			338 => "0000001000000000001001101000010000",
			339 => "0000000001000000001011101000001100",
			340 => "0000000001000000001011101000000100",
			341 => "11111110001110010000010111001101",
			342 => "0000001011000000000100011000000100",
			343 => "11111110111100010000010111001101",
			344 => "00000010011110110000010111001101",
			345 => "11111110010111110000010111001101",
			346 => "0000000100000000000010010000100100",
			347 => "0000001010000000000001010100011100",
			348 => "0000000110000000000100111100001100",
			349 => "0000000110000000000100111100001000",
			350 => "0000000001000000001101101000000100",
			351 => "00000001101110010000010111001101",
			352 => "11111110100111010000010111001101",
			353 => "00000010111011000000010111001101",
			354 => "0000000111000000001111011100001000",
			355 => "0000001000000000001001101000000100",
			356 => "00000000001101010000010111001101",
			357 => "11111110100000000000010111001101",
			358 => "0000000100000000000000010100000100",
			359 => "00000001111111000000010111001101",
			360 => "11111111011001110000010111001101",
			361 => "0000001010000000000001110000000100",
			362 => "00000000111100000000010111001101",
			363 => "00000010000101000000010111001101",
			364 => "0000000100000000000000000000001100",
			365 => "0000001000000000000000110000000100",
			366 => "11111110101011110000010111001101",
			367 => "0000001010000000000001110100000100",
			368 => "00000001100000100000010111001101",
			369 => "11111110110100110000010111001101",
			370 => "11111110011000000000010111001101",
			371 => "0000000111000000001110001101111100",
			372 => "0000000001000000000000011000010000",
			373 => "0000000010000000000001001000001000",
			374 => "0000000100000000000101001100000100",
			375 => "00000001011101010000011101011001",
			376 => "11111110101111100000011101011001",
			377 => "0000001010000000000010101000000100",
			378 => "11111110010111110000011101011001",
			379 => "00000000000000000000011101011001",
			380 => "0000000111000000000100010100111100",
			381 => "0000000011000000000000101000100000",
			382 => "0000000101000000001000111100010000",
			383 => "0000000011000000001010000000001000",
			384 => "0000000000000000001100001000000100",
			385 => "11111111111110000000011101011001",
			386 => "00000001011101100000011101011001",
			387 => "0000000101000000001000111100000100",
			388 => "11111111011101010000011101011001",
			389 => "11111101010010110000011101011001",
			390 => "0000001010000000000101000100001000",
			391 => "0000001001000000001100110100000100",
			392 => "00000000000000000000011101011001",
			393 => "00000001010111000000011101011001",
			394 => "0000001110000000000111000000000100",
			395 => "00000000011010010000011101011001",
			396 => "11111101100100010000011101011001",
			397 => "0000001001000000000010001100001100",
			398 => "0000001100000000000100010100001000",
			399 => "0000001110000000000010111100000100",
			400 => "00000000000010100000011101011001",
			401 => "11111101110000110000011101011001",
			402 => "00000001000111010000011101011001",
			403 => "0000000011000000001000111000001000",
			404 => "0000001011000000000111111000000100",
			405 => "11111110100000100000011101011001",
			406 => "00000000100010000000011101011001",
			407 => "0000000010000000001110010000000100",
			408 => "11111110111000010000011101011001",
			409 => "00000000001111000000011101011001",
			410 => "0000000100000000000000010000010000",
			411 => "0000001110000000001000111000000100",
			412 => "11111111111111100000011101011001",
			413 => "0000000111000000000101101100000100",
			414 => "11111110000001100000011101011001",
			415 => "0000000111000000000101101100000100",
			416 => "00000000010001110000011101011001",
			417 => "11111110011110100000011101011001",
			418 => "0000001010000000000111110100010000",
			419 => "0000001101000000000110000100001000",
			420 => "0000001110000000001010000000000100",
			421 => "00000000100110110000011101011001",
			422 => "11111100110001110000011101011001",
			423 => "0000000100000000001011101100000100",
			424 => "00000000011011110000011101011001",
			425 => "00000001110110000000011101011001",
			426 => "0000001110000000001000111000001000",
			427 => "0000001001000000000111100100000100",
			428 => "00000000011110000000011101011001",
			429 => "00000001001011110000011101011001",
			430 => "0000000010000000000100101000000100",
			431 => "11111111101110100000011101011001",
			432 => "00000000011010000000011101011001",
			433 => "0000001010000000000001010000011000",
			434 => "0000001110000000001010001100001100",
			435 => "0000001101000000000101100100001000",
			436 => "0000001110000000001011000000000100",
			437 => "00000000000000000000011101011001",
			438 => "11111110010100110000011101011001",
			439 => "00000010000100000000011101011001",
			440 => "0000001001000000000001111000001000",
			441 => "0000001001000000000001111000000100",
			442 => "11111110000011100000011101011001",
			443 => "00000000110101110000011101011001",
			444 => "11111110011001010000011101011001",
			445 => "0000000100000000000001001100101000",
			446 => "0000001010000000000001010100011100",
			447 => "0000000010000000001000101000001100",
			448 => "0000000100000000000011011000001000",
			449 => "0000001111000000001100010000000100",
			450 => "00000000101010000000011101011001",
			451 => "00000010110110000000011101011001",
			452 => "11111110010000000000011101011001",
			453 => "0000000111000000001111011100001000",
			454 => "0000001001000000000101010000000100",
			455 => "11111111110000000000011101011001",
			456 => "11111110010010010000011101011001",
			457 => "0000001111000000000010111000000100",
			458 => "00000001010000100000011101011001",
			459 => "11111111001100100000011101011001",
			460 => "0000001010000000001100000100001000",
			461 => "0000001111000000000000010100000100",
			462 => "00000001101100010000011101011001",
			463 => "11111110100110010000011101011001",
			464 => "00000011000001000000011101011001",
			465 => "0000000100000000000000000000001000",
			466 => "0000000100000000001010101000000100",
			467 => "11111110011100100000011101011001",
			468 => "00000000000000000000011101011001",
			469 => "11111110011000100000011101011001",
			470 => "0000000100000000000000101110011000",
			471 => "0000000101000000000100011000111100",
			472 => "0000000111000000001101100000101000",
			473 => "0000000001000000000110101000100000",
			474 => "0000001111000000001011011100010000",
			475 => "0000001110000000000000111000001000",
			476 => "0000001011000000000100010100000100",
			477 => "11111111111010000000100100000101",
			478 => "00000000011111010000100100000101",
			479 => "0000001010000000000001010000000100",
			480 => "11111111111001100000100100000101",
			481 => "11111111001100010000100100000101",
			482 => "0000000110000000000100110100001000",
			483 => "0000000101000000000100001000000100",
			484 => "00000000010001000000100100000101",
			485 => "00000001011000010000100100000101",
			486 => "0000001100000000001010000000000100",
			487 => "00000001011001000000100100000101",
			488 => "00000000000000110000100100000101",
			489 => "0000000100000000001000000100000100",
			490 => "00000010111101000000100100000101",
			491 => "00000000000011100000100100000101",
			492 => "0000001111000000001110000100001100",
			493 => "0000000110000000001100011000001000",
			494 => "0000001110000000001101111000000100",
			495 => "00000001011000110000100100000101",
			496 => "11111110101100100000100100000101",
			497 => "00000001111111100000100100000101",
			498 => "0000001100000000001000111000000100",
			499 => "11111110111001000000100100000101",
			500 => "00000001101010000000100100000101",
			501 => "0000001010000000000110011000101100",
			502 => "0000000010000000000101110000011100",
			503 => "0000000010000000001111010000001100",
			504 => "0000001111000000000101110100001000",
			505 => "0000001111000000000110110100000100",
			506 => "11111110111011110000100100000101",
			507 => "00000000111001100000100100000101",
			508 => "11111110010111110000100100000101",
			509 => "0000000010000000000010011100001000",
			510 => "0000000110000000000111101000000100",
			511 => "00000000000000000000100100000101",
			512 => "00000010100101110000100100000101",
			513 => "0000000010000000000101110000000100",
			514 => "11111110110000110000100100000101",
			515 => "00000010000111110000100100000101",
			516 => "0000000101000000000011100000000100",
			517 => "11111101101111000000100100000101",
			518 => "0000000101000000001000000000000100",
			519 => "00000001100101000000100100000101",
			520 => "0000001000000000001011010100000100",
			521 => "11111110111100000000100100000101",
			522 => "11111100101010110000100100000101",
			523 => "0000001100000000001000111000010100",
			524 => "0000001110000000000001101000000100",
			525 => "11111101111100110000100100000101",
			526 => "0000000110000000001001100100001000",
			527 => "0000000001000000000111100100000100",
			528 => "00000001000001000000100100000101",
			529 => "11111110100110100000100100000101",
			530 => "0000001111000000001100010000000100",
			531 => "11111110010110100000100100000101",
			532 => "00000000001011110000100100000101",
			533 => "0000000000000000000010111100010000",
			534 => "0000001111000000000101000000001000",
			535 => "0000000100000000000010111000000100",
			536 => "00000000110110010000100100000101",
			537 => "00000010100100000000100100000101",
			538 => "0000001010000000001100011100000100",
			539 => "11111110101001000000100100000101",
			540 => "00000001010100010000100100000101",
			541 => "0000001100000000001000111000000100",
			542 => "00000001101010010000100100000101",
			543 => "0000001100000000001100110000000100",
			544 => "11111111011110110000100100000101",
			545 => "00000000100011100000100100000101",
			546 => "0000001000000000001101010000100000",
			547 => "0000000001000000000110000000001100",
			548 => "0000000100000000000110110000001000",
			549 => "0000000001000000000000011000000100",
			550 => "11111111100100100000100100000101",
			551 => "00000001011101010000100100000101",
			552 => "11111110101100010000100100000101",
			553 => "0000001100000000000000101000000100",
			554 => "11111100010101010000100100000101",
			555 => "0000000000000000001100001000000100",
			556 => "11111110010111010000100100000101",
			557 => "0000000110000000001011001100000100",
			558 => "00000000101111110000100100000101",
			559 => "0000000001000000001011101000000100",
			560 => "11111111000101100000100100000101",
			561 => "00000000000000000000100100000101",
			562 => "0000000100000000000101100000011000",
			563 => "0000000000000000000011011100001000",
			564 => "0000000001000000001011101000000100",
			565 => "11111101110010010000100100000101",
			566 => "00000000011100010000100100000101",
			567 => "0000001101000000001000111000000100",
			568 => "11111111000000010000100100000101",
			569 => "0000001011000000000000101000000100",
			570 => "00000001101000110000100100000101",
			571 => "0000000111000000001000111000000100",
			572 => "11111110111111000000100100000101",
			573 => "00000000111100000000100100000101",
			574 => "0000001100000000000000111000000100",
			575 => "00000000000000000000100100000101",
			576 => "11111110100011010000100100000101",
			577 => "0000000100000000000110110010011100",
			578 => "0000001001000000001100011001101000",
			579 => "0000000010000000001001010000111000",
			580 => "0000001110000000001000111000011000",
			581 => "0000001101000000001100101000001100",
			582 => "0000000111000000000100000000001000",
			583 => "0000000110000000000111101000000100",
			584 => "00000000011011010000101010011001",
			585 => "11111111111101000000101010011001",
			586 => "11111101011101010000101010011001",
			587 => "0000000001000000000010001100001000",
			588 => "0000000010000000001111010000000100",
			589 => "00000001101110100000101010011001",
			590 => "11111111101110000000101010011001",
			591 => "11111110111001110000101010011001",
			592 => "0000001001000000000111100100010000",
			593 => "0000000011000000001100101100001000",
			594 => "0000001001000000000110101000000100",
			595 => "11111110001001110000101010011001",
			596 => "00000001010101100000101010011001",
			597 => "0000000101000000000110000100000100",
			598 => "00000000110110110000101010011001",
			599 => "11111110001111000000101010011001",
			600 => "0000000101000000001101111000001000",
			601 => "0000001110000000000101101100000100",
			602 => "00000010110001100000101010011001",
			603 => "00000000000000000000101010011001",
			604 => "0000000000000000000010011000000100",
			605 => "00000000000000000000101010011001",
			606 => "11111110011000010000101010011001",
			607 => "0000000010000000000010011100010000",
			608 => "0000000110000000000001111000000100",
			609 => "00000000011011110000101010011001",
			610 => "0000000000000000000010111100000100",
			611 => "00000100001111100000101010011001",
			612 => "0000000111000000001100001000000100",
			613 => "00000010010110110000101010011001",
			614 => "11111111111111100000101010011001",
			615 => "0000001000000000000111000000010000",
			616 => "0000000001000000000110000000001000",
			617 => "0000000101000000001000111000000100",
			618 => "11111101010010110000101010011001",
			619 => "11111111001100110000101010011001",
			620 => "0000001000000000000110001000000100",
			621 => "00000000011010110000101010011001",
			622 => "00000000000110110000101010011001",
			623 => "0000001111000000000101100100001000",
			624 => "0000001011000000001011000100000100",
			625 => "00000001101010100000101010011001",
			626 => "11111110011110110000101010011001",
			627 => "0000000110000000001011001100000100",
			628 => "00000001101000000000101010011001",
			629 => "00000000001001000000101010011001",
			630 => "0000000110000000001001111100100000",
			631 => "0000001000000000001001101000000100",
			632 => "11111110011001000000101010011001",
			633 => "0000000111000000000110100100001100",
			634 => "0000000010000000001100001100001000",
			635 => "0000000110000000000100111100000100",
			636 => "11111111011000000000101010011001",
			637 => "11111110001111000000101010011001",
			638 => "00000000000101110000101010011001",
			639 => "0000000010000000001100001100001000",
			640 => "0000001001000000000100101100000100",
			641 => "00000001100000010000101010011001",
			642 => "00000000000000000000101010011001",
			643 => "0000001001000000000100101100000100",
			644 => "11111111100110000000101010011001",
			645 => "11111110011000000000101010011001",
			646 => "0000001110000000000010110000001100",
			647 => "0000000100000000001110111000000100",
			648 => "11111111000001010000101010011001",
			649 => "0000000111000000001111011100000100",
			650 => "00000000110000000000101010011001",
			651 => "00000010001001010000101010011001",
			652 => "0000000111000000001001010100000100",
			653 => "11111110100010000000101010011001",
			654 => "00000000111000110000101010011001",
			655 => "0000000110000000001011001100010100",
			656 => "0000000100000000000011111000000100",
			657 => "11111101101011010000101010011001",
			658 => "0000000100000000001101000000001000",
			659 => "0000001001000000000110000000000100",
			660 => "00000000000000000000101010011001",
			661 => "00000000010001010000101010011001",
			662 => "0000000001000000000000011000000100",
			663 => "11111110011010100000101010011001",
			664 => "11111111101101010000101010011001",
			665 => "0000000010000000000010000100001000",
			666 => "0000000001000000001110011100000100",
			667 => "11111111101100110000101010011001",
			668 => "00000001101010000000101010011001",
			669 => "0000001000000000000010011000010000",
			670 => "0000001000000000001111000100000100",
			671 => "11111110101010110000101010011001",
			672 => "0000000010000000000010010100000100",
			673 => "11111111110110110000101010011001",
			674 => "0000000001000000001011101000000100",
			675 => "00000010000011000000101010011001",
			676 => "00000000000000000000101010011001",
			677 => "11111110100001100000101010011001",
			678 => "0000000100000000001011101100011000",
			679 => "0000000110000000000001111000010100",
			680 => "0000001001000000001101101000001000",
			681 => "0000000101000000001100101100000100",
			682 => "11111101101001110000110000000101",
			683 => "11111111001101000000110000000101",
			684 => "0000000000000000001011010100000100",
			685 => "11111110011101010000110000000101",
			686 => "0000000111000000000100000000000100",
			687 => "00000000011000110000110000000101",
			688 => "00000001100010110000110000000101",
			689 => "11111110001110110000110000000101",
			690 => "0000000100000000000011011001011000",
			691 => "0000000000000000001100001000110100",
			692 => "0000000101000000001000111100010100",
			693 => "0000000101000000001000111100010000",
			694 => "0000000010000000001110000100001000",
			695 => "0000000110000000000001111000000100",
			696 => "11111111100101010000110000000101",
			697 => "00000001100001100000110000000101",
			698 => "0000000011000000000100010100000100",
			699 => "11111110111111100000110000000101",
			700 => "11111101001011110000110000000101",
			701 => "11111100111100010000110000000101",
			702 => "0000001011000000000111111000010000",
			703 => "0000000100000000000000010100001000",
			704 => "0000000011000000000100000000000100",
			705 => "00000001100011010000110000000101",
			706 => "11111111111011010000110000000101",
			707 => "0000000111000000000111111000000100",
			708 => "11111111001010000000110000000101",
			709 => "00000001010100100000110000000101",
			710 => "0000001011000000000111111000001000",
			711 => "0000001100000000000111111000000100",
			712 => "11111100101111100000110000000101",
			713 => "00000000100110010000110000000101",
			714 => "0000001001000000000110101000000100",
			715 => "11111111111010010000110000000101",
			716 => "00000000000111100000110000000101",
			717 => "0000001110000000000000101000011000",
			718 => "0000001011000000000111111000001100",
			719 => "0000000101000000001000111100001000",
			720 => "0000000101000000001000111100000100",
			721 => "00000001110001000000110000000101",
			722 => "00000000101000000000110000000101",
			723 => "11111110111011000000110000000101",
			724 => "0000001010000000000001010100001000",
			725 => "0000000111000000000000101000000100",
			726 => "00000001110101010000110000000101",
			727 => "00000001000011100000110000000101",
			728 => "00000000000010010000110000000101",
			729 => "0000001110000000000100000000000100",
			730 => "11111101010100010000110000000101",
			731 => "0000000001000000000010001100000100",
			732 => "00000001101100010000110000000101",
			733 => "11111111100100100000110000000101",
			734 => "0000001111000000001001010100100100",
			735 => "0000001110000000001011000100100000",
			736 => "0000000111000000000111111000010000",
			737 => "0000001010000000001001101000001000",
			738 => "0000001011000000001110111100000100",
			739 => "11111110011111110000110000000101",
			740 => "11111100111100010000110000000101",
			741 => "0000000101000000000100000000000100",
			742 => "11111111000011100000110000000101",
			743 => "00000000000000000000110000000101",
			744 => "0000001100000000000111111000001000",
			745 => "0000000100000000000110110000000100",
			746 => "00000001100001110000110000000101",
			747 => "11111111001000110000110000000101",
			748 => "0000000010000000000011001000000100",
			749 => "11111110110101100000110000000101",
			750 => "00000000110001110000110000000101",
			751 => "11111100101011100000110000000101",
			752 => "0000000111000000001101111000010100",
			753 => "0000000010000000001100010000001000",
			754 => "0000000011000000001101111000000100",
			755 => "00000001110100100000110000000101",
			756 => "11111110000010000000110000000101",
			757 => "0000000000000000001100001000000100",
			758 => "11111111011011100000110000000101",
			759 => "0000000100000000000001001100000100",
			760 => "00000001110011100000110000000101",
			761 => "11111111100001010000110000000101",
			762 => "0000000000000000000100010100000100",
			763 => "11111110011011010000110000000101",
			764 => "0000000001000000001001011000001000",
			765 => "0000000011000000001101000100000100",
			766 => "00000000011010100000110000000101",
			767 => "11111110101111100000110000000101",
			768 => "00000001001011110000110000000101",
			769 => "0000001000000000000111000001110000",
			770 => "0000000010000000000010110100101100",
			771 => "0000000110000000001101111100101000",
			772 => "0000001010000000001000010100010100",
			773 => "0000000010000000001110101100001100",
			774 => "0000000110000000000001111000001000",
			775 => "0000000100000000001011110000000100",
			776 => "11111111101011010000110110001001",
			777 => "00000000111100000000110110001001",
			778 => "11111111000011000000110110001001",
			779 => "0000000110000000000111101000000100",
			780 => "11111111010111010000110110001001",
			781 => "11111101110100000000110110001001",
			782 => "0000001101000000000110000100010000",
			783 => "0000000110000000000001111000001000",
			784 => "0000001101000000000011011100000100",
			785 => "00000000000000000000110110001001",
			786 => "00000001100100110000110110001001",
			787 => "0000000110000000001101111100000100",
			788 => "11111110110010110000110110001001",
			789 => "00000000000111110000110110001001",
			790 => "00000001111110100000110110001001",
			791 => "11111110000011010000110110001001",
			792 => "0000000010000000000010110100001000",
			793 => "0000001111000000001000011000000100",
			794 => "00000001101001000000110110001001",
			795 => "00000000011000010000110110001001",
			796 => "0000000100000000000010110000011100",
			797 => "0000000011000000001000111000001100",
			798 => "0000001111000000000100000100001000",
			799 => "0000001110000000000000110000000100",
			800 => "00000001000101010000110110001001",
			801 => "11111111011010100000110110001001",
			802 => "00000001111101000000110110001001",
			803 => "0000001101000000000101101100001000",
			804 => "0000000110000000000111101000000100",
			805 => "11111110000101010000110110001001",
			806 => "11111111011111100000110110001001",
			807 => "0000000011000000000110000100000100",
			808 => "00000000100110100000110110001001",
			809 => "00000000000010100000110110001001",
			810 => "0000000100000000000010110000010000",
			811 => "0000001001000000000111100100001000",
			812 => "0000000110000000000111101000000100",
			813 => "00000001011101000000110110001001",
			814 => "11111110100000000000110110001001",
			815 => "0000001101000000001101111000000100",
			816 => "00000001000001010000110110001001",
			817 => "11111111011011110000110110001001",
			818 => "0000000100000000001000001000001000",
			819 => "0000001100000000000011011100000100",
			820 => "00000001110000100000110110001001",
			821 => "11111110001101100000110110001001",
			822 => "0000000101000000001010111100000100",
			823 => "00000000000001010000110110001001",
			824 => "11111111101101000000110110001001",
			825 => "0000001010000000000101000100010000",
			826 => "0000000110000000001010011000001000",
			827 => "0000000001000000000000011000000100",
			828 => "00000000000000000000110110001001",
			829 => "00000001100100010000110110001001",
			830 => "0000000010000000001100010100000100",
			831 => "11111111000010100000110110001001",
			832 => "00000000111111010000110110001001",
			833 => "0000001100000000000000110000001000",
			834 => "0000001010000000001011010100000100",
			835 => "11111101110101010000110110001001",
			836 => "00000000000000000000110110001001",
			837 => "0000000110000000001100011000100000",
			838 => "0000000111000000000100010100010000",
			839 => "0000000111000000000111111000001000",
			840 => "0000001110000000001100011100000100",
			841 => "00000000110010010000110110001001",
			842 => "11111110011000100000110110001001",
			843 => "0000000001000000000000011000000100",
			844 => "00000000000000000000110110001001",
			845 => "00000001101000110000110110001001",
			846 => "0000000010000000000111111100001000",
			847 => "0000001000000000000010111100000100",
			848 => "11111110000010100000110110001001",
			849 => "00000000000000000000110110001001",
			850 => "0000001100000000000110000100000100",
			851 => "00000000001100100000110110001001",
			852 => "00000000000000000000110110001001",
			853 => "0000000100000000001011100000001100",
			854 => "0000000100000000000011101100001000",
			855 => "0000000110000000001011001100000100",
			856 => "00000001010011100000110110001001",
			857 => "11111111011011000000110110001001",
			858 => "11111110000110110000110110001001",
			859 => "0000000100000000000110110000001000",
			860 => "0000001000000000001000101100000100",
			861 => "00000000000000000000110110001001",
			862 => "00000001001101010000110110001001",
			863 => "0000001000000000000011010000000100",
			864 => "11111111010100100000110110001001",
			865 => "00000000100010100000110110001001",
			866 => "0000000111000000001101111010011000",
			867 => "0000000001000000000000011000100000",
			868 => "0000000001000000001100100000000100",
			869 => "11111110010110110000111100111101",
			870 => "0000000011000000000000111000001100",
			871 => "0000001011000000001110111100000100",
			872 => "11111110111101010000111100111101",
			873 => "0000000010000000001110101000000100",
			874 => "00000010001110010000111100111101",
			875 => "00000000000000000000111100111101",
			876 => "0000001010000000001100011100001100",
			877 => "0000001000000000000010101000001000",
			878 => "0000000010000000001101000100000100",
			879 => "11111111101101110000111100111101",
			880 => "11111110001001100000111100111101",
			881 => "00000000000000000000111100111101",
			882 => "11111101010101100000111100111101",
			883 => "0000001110000000000000001101000000",
			884 => "0000000111000000001100001000100000",
			885 => "0000000011000000001001110000010000",
			886 => "0000000111000000000111111000001000",
			887 => "0000000010000000000001000000000100",
			888 => "00000000100010000000111100111101",
			889 => "11111110110000000000111100111101",
			890 => "0000000011000000000111111000000100",
			891 => "00000001011110010000111100111101",
			892 => "00000000110101100000111100111101",
			893 => "0000000010000000000101110000001000",
			894 => "0000001110000000001100001000000100",
			895 => "00000000010000100000111100111101",
			896 => "11111111100001000000111100111101",
			897 => "0000001100000000001110111100000100",
			898 => "11111111010001000000111100111101",
			899 => "00000000110000000000111100111101",
			900 => "0000000111000000001100001000010000",
			901 => "0000001010000000001100011100001000",
			902 => "0000001101000000000000001100000100",
			903 => "00000001101010100000111100111101",
			904 => "00000010101101110000111100111101",
			905 => "0000000100000000000100001100000100",
			906 => "11111111110000100000111100111101",
			907 => "00000001011100000000111100111101",
			908 => "0000000111000000000100000000001000",
			909 => "0000000101000000000100001000000100",
			910 => "00000000000010110000111100111101",
			911 => "00000001110010010000111100111101",
			912 => "0000001110000000001000111000000100",
			913 => "00000001011011100000111100111101",
			914 => "00000000110011000000111100111101",
			915 => "0000000010000000000011001000011100",
			916 => "0000000110000000001010011000010000",
			917 => "0000001010000000001000010100001000",
			918 => "0000000100000000001000000100000100",
			919 => "11111111001110110000111100111101",
			920 => "00000010111001000000111100111101",
			921 => "0000001100000000000100000000000100",
			922 => "11111110000101100000111100111101",
			923 => "00000000000000000000111100111101",
			924 => "0000000010000000000101110000000100",
			925 => "00000011001001010000111100111101",
			926 => "0000001011000000001101100000000100",
			927 => "11111111000000000000111100111101",
			928 => "00000000111101000000111100111101",
			929 => "0000000110000000001100011000001100",
			930 => "0000000001000000001100110100000100",
			931 => "11111101111101100000111100111101",
			932 => "0000001011000000000101101100000100",
			933 => "00000011010101000000111100111101",
			934 => "00000000000100010000111100111101",
			935 => "0000001100000000001000111000001000",
			936 => "0000000110000000001001100100000100",
			937 => "00000000001101110000111100111101",
			938 => "11111110111111100000111100111101",
			939 => "0000000001000000001011101000000100",
			940 => "00000001010001110000111100111101",
			941 => "11111110011001010000111100111101",
			942 => "0000001000000000001001101000001100",
			943 => "0000000001000000001011101000001000",
			944 => "0000000001000000001011101000000100",
			945 => "11111110011110000000111100111101",
			946 => "00000010001101100000111100111101",
			947 => "11111110010111000000111100111101",
			948 => "0000000100000000000010010000101000",
			949 => "0000001000000000000001110100011000",
			950 => "0000001110000000001011110000001100",
			951 => "0000000100000000001011100000001000",
			952 => "0000000100000000001000001000000100",
			953 => "11111111000011010000111100111101",
			954 => "00000001110011000000111100111101",
			955 => "11111110001001010000111100111101",
			956 => "0000000110000000001001111100000100",
			957 => "11111110010101000000111100111101",
			958 => "0000000110000000000100101100000100",
			959 => "00000000101000110000111100111101",
			960 => "11111110010111000000111100111101",
			961 => "0000000100000000001101110100001000",
			962 => "0000000111000000001111011100000100",
			963 => "00000001000100010000111100111101",
			964 => "00000010011010010000111100111101",
			965 => "0000001000000000001010101100000100",
			966 => "11111110000101110000111100111101",
			967 => "00000001110100010000111100111101",
			968 => "0000000100000000000000000000001100",
			969 => "0000001000000000000000110000000100",
			970 => "11111110100100110000111100111101",
			971 => "0000001010000000000001110100000100",
			972 => "00000001100110000000111100111101",
			973 => "11111110101000110000111100111101",
			974 => "11111110010110110000111100111101",
			975 => "0000001101000000001011000010011100",
			976 => "0000000111000000000111111001000000",
			977 => "0000000111000000001110111100101000",
			978 => "0000001100000000001010000000010000",
			979 => "0000001011000000000111111000001100",
			980 => "0000000100000000001011100000001000",
			981 => "0000000000000000000011111100000100",
			982 => "11111110000100100001000100011001",
			983 => "00000001111011100001000100011001",
			984 => "11111110011001010001000100011001",
			985 => "11111101011001010001000100011001",
			986 => "0000000100000000000011010100001000",
			987 => "0000000010000000000101001000000100",
			988 => "00000001110100100001000100011001",
			989 => "11111111000100000001000100011001",
			990 => "0000001010000000000110011100001000",
			991 => "0000000101000000001000111000000100",
			992 => "00000000101110010001000100011001",
			993 => "11111101000010110001000100011001",
			994 => "0000000011000000000010011000000100",
			995 => "11111110101101000001000100011001",
			996 => "00000001101011100001000100011001",
			997 => "0000001010000000001010110000010000",
			998 => "0000000110000000001011111100001000",
			999 => "0000001111000000000111010000000100",
			1000 => "00000001100000000001000100011001",
			1001 => "11111111100011000001000100011001",
			1002 => "0000000001000000001110100000000100",
			1003 => "11111100011110000001000100011001",
			1004 => "11111110100111100001000100011001",
			1005 => "0000001000000000000111000000000100",
			1006 => "00000001001100010001000100011001",
			1007 => "11111110011100110001000100011001",
			1008 => "0000001010000000001001000100111000",
			1009 => "0000000010000000001110000100011100",
			1010 => "0000000101000000000011011100001100",
			1011 => "0000000011000000001000111000001000",
			1012 => "0000000111000000000100010100000100",
			1013 => "11111110000111110001000100011001",
			1014 => "00000000011010010001000100011001",
			1015 => "11111100001010100001000100011001",
			1016 => "0000000011000000001101100000001000",
			1017 => "0000000101000000000101101100000100",
			1018 => "00000000010000100001000100011001",
			1019 => "00000001010101000001000100011001",
			1020 => "0000001000000000000001110000000100",
			1021 => "00000000010111000001000100011001",
			1022 => "11111111001110100001000100011001",
			1023 => "0000000100000000001100001100010000",
			1024 => "0000001010000000001000010100001000",
			1025 => "0000000100000000001011110000000100",
			1026 => "00000000000010100001000100011001",
			1027 => "00000001101100110001000100011001",
			1028 => "0000000100000000000010010100000100",
			1029 => "00000011000100110001000100011001",
			1030 => "11111111010111110001000100011001",
			1031 => "0000001000000000000001110000000100",
			1032 => "11111101111001000001000100011001",
			1033 => "0000001111000000001011011100000100",
			1034 => "00000000000110100001000100011001",
			1035 => "00000001011011010001000100011001",
			1036 => "0000000000000000001111000100000100",
			1037 => "00000011000100000001000100011001",
			1038 => "0000000100000000000010110000010000",
			1039 => "0000000111000000000100010100001000",
			1040 => "0000000010000000000010011100000100",
			1041 => "00000000001011110001000100011001",
			1042 => "00000011000000100001000100011001",
			1043 => "0000000101000000001010111000000100",
			1044 => "11111111011001100001000100011001",
			1045 => "00000001111001000001000100011001",
			1046 => "0000000111000000001100001000001000",
			1047 => "0000000111000000001100001000000100",
			1048 => "00000000001001000001000100011001",
			1049 => "11111111010010000001000100011001",
			1050 => "0000000111000000001100001000000100",
			1051 => "00000000110101100001000100011001",
			1052 => "00000000001100000001000100011001",
			1053 => "0000000000000000000111000000011000",
			1054 => "0000000101000000001000000000010000",
			1055 => "0000000111000000001101100000001000",
			1056 => "0000001101000000001001001000000100",
			1057 => "11111111010010010001000100011001",
			1058 => "00000000101011010001000100011001",
			1059 => "0000000000000000001010100000000100",
			1060 => "11111111011110010001000100011001",
			1061 => "00000010000110100001000100011001",
			1062 => "0000001000000000000001110000000100",
			1063 => "11111110011000110001000100011001",
			1064 => "00000000001011000001000100011001",
			1065 => "0000000100000000000000000000111000",
			1066 => "0000001011000000001100101100011100",
			1067 => "0000000011000000000100000100001100",
			1068 => "0000000001000000001001111000000100",
			1069 => "11111110110110110001000100011001",
			1070 => "0000001111000000000111100000000100",
			1071 => "00000000010001010001000100011001",
			1072 => "00000001011101110001000100011001",
			1073 => "0000001010000000000001010000001000",
			1074 => "0000001111000000001001010000000100",
			1075 => "11111110001010100001000100011001",
			1076 => "00000001101000100001000100011001",
			1077 => "0000000110000000001011001100000100",
			1078 => "11111100111111010001000100011001",
			1079 => "11111110001111100001000100011001",
			1080 => "0000000011000000000100000100001100",
			1081 => "0000000101000000001001001000001000",
			1082 => "0000000011000000001010001100000100",
			1083 => "00000000001010010001000100011001",
			1084 => "11111101111011010001000100011001",
			1085 => "11111101001110100001000100011001",
			1086 => "0000000110000000000100111100001000",
			1087 => "0000000111000000001101100000000100",
			1088 => "11111111011000100001000100011001",
			1089 => "00000000110011100001000100011001",
			1090 => "0000001000000000001001101000000100",
			1091 => "11111110011100000001000100011001",
			1092 => "11111111110100010001000100011001",
			1093 => "11111110011010100001000100011001",
			1094 => "0000000100000000000001001110111100",
			1095 => "0000000011000000001011000101010000",
			1096 => "0000000110000000000001111000100100",
			1097 => "0000000010000000000010110100010000",
			1098 => "0000001011000000001110111100000100",
			1099 => "11111101100111110001001010111101",
			1100 => "0000000100000000001110000000000100",
			1101 => "11111111011011010001001010111101",
			1102 => "0000001100000000001110111100000100",
			1103 => "00000000010000010001001010111101",
			1104 => "00000001101111010001001010111101",
			1105 => "0000001000000000000110001000001100",
			1106 => "0000001011000000000111111000001000",
			1107 => "0000000011000000000100010100000100",
			1108 => "00000000001111000001001010111101",
			1109 => "11111100010010100001001010111101",
			1110 => "11111100100000000001001010111101",
			1111 => "0000001100000000000000111000000100",
			1112 => "00000000000000000001001010111101",
			1113 => "00000001101010000001001010111101",
			1114 => "0000000100000000000000010100011000",
			1115 => "0000001111000000000001101000010000",
			1116 => "0000000110000000001101111100001000",
			1117 => "0000000010000000000110100000000100",
			1118 => "00000001111000110001001010111101",
			1119 => "00000000100001110001001010111101",
			1120 => "0000001110000000001000110000000100",
			1121 => "00000001001100110001001010111101",
			1122 => "11111111001111110001001010111101",
			1123 => "0000001000000000000110001000000100",
			1124 => "00000000110101110001001010111101",
			1125 => "00000001111101010001001010111101",
			1126 => "0000000000000000000111111000001000",
			1127 => "0000001110000000001111000100000100",
			1128 => "00000000000000000001001010111101",
			1129 => "11111100001110110001001010111101",
			1130 => "0000001111000000000001011000001000",
			1131 => "0000000010000000000101110000000100",
			1132 => "00000000011111000001001010111101",
			1133 => "11111110010111110001001010111101",
			1134 => "00000010000101010001001010111101",
			1135 => "0000000101000000000011011100101100",
			1136 => "0000001110000000000010011000001100",
			1137 => "0000000101000000001001110000001000",
			1138 => "0000000011000000001100001000000100",
			1139 => "00000000110011010001001010111101",
			1140 => "11111101111100110001001010111101",
			1141 => "11111010011001010001001010111101",
			1142 => "0000000001000000001110100000010000",
			1143 => "0000000001000000000110000000001000",
			1144 => "0000000000000000001011000100000100",
			1145 => "11111110011110110001001010111101",
			1146 => "00000000100011110001001010111101",
			1147 => "0000000110000000000100110100000100",
			1148 => "00000000101011110001001010111101",
			1149 => "11111101101100100001001010111101",
			1150 => "0000001011000000000100010100001000",
			1151 => "0000000111000000000111111000000100",
			1152 => "00000000000000000001001010111101",
			1153 => "11111100001010100001001010111101",
			1154 => "0000000011000000001000111000000100",
			1155 => "00000001001001000001001010111101",
			1156 => "11111110110110100001001010111101",
			1157 => "0000001011000000001011000100100000",
			1158 => "0000001011000000000100010100010000",
			1159 => "0000000100000000000101010100001000",
			1160 => "0000000110000000000001111000000100",
			1161 => "00000001000000110001001010111101",
			1162 => "11111101110100010001001010111101",
			1163 => "0000001011000000000111111000000100",
			1164 => "00000001111010010001001010111101",
			1165 => "00000000011110000001001010111101",
			1166 => "0000001100000000001110111100001000",
			1167 => "0000001010000000000110011000000100",
			1168 => "00000001111001000001001010111101",
			1169 => "11111110000101000001001010111101",
			1170 => "0000001111000000000101110100000100",
			1171 => "00000000111111000001001010111101",
			1172 => "00000010010101100001001010111101",
			1173 => "0000000111000000000100010100010000",
			1174 => "0000001111000000001010010100001000",
			1175 => "0000000101000000001101100000000100",
			1176 => "00000000100111100001001010111101",
			1177 => "11111110100101010001001010111101",
			1178 => "0000000010000000000011001000000100",
			1179 => "00000011011010100001001010111101",
			1180 => "11111111100110010001001010111101",
			1181 => "0000000011000000001100001000001000",
			1182 => "0000001111000000001000011000000100",
			1183 => "11111101001110000001001010111101",
			1184 => "11111111111101110001001010111101",
			1185 => "0000000011000000000100000000000100",
			1186 => "00000001000010100001001010111101",
			1187 => "00000000000101010001001010111101",
			1188 => "0000000111000000001100001000010100",
			1189 => "0000001100000000000111111000001100",
			1190 => "0000000101000000001001110000000100",
			1191 => "11111110100101110001001010111101",
			1192 => "0000000101000000000011011100000100",
			1193 => "00000000101000110001001010111101",
			1194 => "11111110010010000001001010111101",
			1195 => "0000000010000000001111010000000100",
			1196 => "11111111100010100001001010111101",
			1197 => "00000001001110110001001010111101",
			1198 => "11111110011010010001001010111101",
			1199 => "0000001100000000000100000010010000",
			1200 => "0000000111000000001001110001100100",
			1201 => "0000000101000000001010111100110000",
			1202 => "0000001100000000000100000000010100",
			1203 => "0000001001000000001111001100010000",
			1204 => "0000001001000000000110101000001000",
			1205 => "0000000011000000000011011100000100",
			1206 => "00000000000010010001010011010001",
			1207 => "11111111100101010001010011010001",
			1208 => "0000000001000000001110100000000100",
			1209 => "00000001101001010001010011010001",
			1210 => "00000000000101000001010011010001",
			1211 => "00000001111000110001010011010001",
			1212 => "0000001011000000001000111000010000",
			1213 => "0000001010000000001010110000001000",
			1214 => "0000001000000000001011010100000100",
			1215 => "11111111100111000001010011010001",
			1216 => "00000001111101110001010011010001",
			1217 => "0000000100000000000100001100000100",
			1218 => "11111101101111110001010011010001",
			1219 => "00000001011000110001010011010001",
			1220 => "0000001000000000000001110100001000",
			1221 => "0000001010000000001001000100000100",
			1222 => "00000000000010010001010011010001",
			1223 => "00000010001110100001010011010001",
			1224 => "11111111111111000001010011010001",
			1225 => "0000001001000000001101011100100000",
			1226 => "0000001011000000001101100000010000",
			1227 => "0000001100000000000100000000001000",
			1228 => "0000000111000000000100000000000100",
			1229 => "11111110010110010001010011010001",
			1230 => "00000000000000000001010011010001",
			1231 => "0000000111000000001000111000000100",
			1232 => "00000010010001110001010011010001",
			1233 => "11111110111010010001010011010001",
			1234 => "0000001111000000001110101100001000",
			1235 => "0000001001000000001011101000000100",
			1236 => "11111110111010010001010011010001",
			1237 => "00000001000011010001010011010001",
			1238 => "0000001011000000001100110000000100",
			1239 => "11111101101101010001010011010001",
			1240 => "11111111010010010001010011010001",
			1241 => "0000001100000000000000101000000100",
			1242 => "00000010010100000001010011010001",
			1243 => "0000001110000000001000000000001000",
			1244 => "0000000010000000000010000000000100",
			1245 => "11111111111011100001010011010001",
			1246 => "00000010001011100001010011010001",
			1247 => "0000000010000000001110110100000100",
			1248 => "11111110100000010001010011010001",
			1249 => "00000000110101110001010011010001",
			1250 => "0000001000000000000001110100100100",
			1251 => "0000000101000000001010111000001100",
			1252 => "0000000010000000000101110000000100",
			1253 => "11111111010110000001010011010001",
			1254 => "0000001000000000000111000100000100",
			1255 => "00000010001101110001010011010001",
			1256 => "00000001000000110001010011010001",
			1257 => "0000001101000000000110100100001100",
			1258 => "0000001010000000001010110000001000",
			1259 => "0000001011000000001100101100000100",
			1260 => "00000001000011100001010011010001",
			1261 => "11111110001000010001010011010001",
			1262 => "11111110100101010001010011010001",
			1263 => "0000001001000000001011111100001000",
			1264 => "0000000010000000001100010000000100",
			1265 => "00000000110110100001010011010001",
			1266 => "00000010001010110001010011010001",
			1267 => "11111111101100010001010011010001",
			1268 => "0000001000000000000010101000000100",
			1269 => "11111101101001100001010011010001",
			1270 => "00000000101011100001010011010001",
			1271 => "0000001100000000000100000000100000",
			1272 => "0000000101000000001010111000011000",
			1273 => "0000001101000000000001111100001000",
			1274 => "0000001111000000001110101100000100",
			1275 => "11111110110101110001010011010001",
			1276 => "00000000110111010001010011010001",
			1277 => "0000001010000000001100011100001100",
			1278 => "0000000001000000001001111000001000",
			1279 => "0000000010000000000100101000000100",
			1280 => "11111111000111000001010011010001",
			1281 => "11111101100011110001010011010001",
			1282 => "11111111100101110001010011010001",
			1283 => "11111111101110010001010011010001",
			1284 => "0000001110000000001000011000000100",
			1285 => "00000001111011110001010011010001",
			1286 => "11111110111011000001010011010001",
			1287 => "0000001100000000001000111100100100",
			1288 => "0000001100000000001000111100010100",
			1289 => "0000000111000000001001110000001100",
			1290 => "0000001111000000000100010000000100",
			1291 => "00000010010101010001010011010001",
			1292 => "0000000010000000001010001000000100",
			1293 => "11111110111001100001010011010001",
			1294 => "00000000101011000001010011010001",
			1295 => "0000001000000000000111000100000100",
			1296 => "11111101101100000001010011010001",
			1297 => "00000000100101010001010011010001",
			1298 => "0000001000000000001011010100001000",
			1299 => "0000001010000000000110011000000100",
			1300 => "00000001111110110001010011010001",
			1301 => "11111101100100110001010011010001",
			1302 => "0000000010000000001100000000000100",
			1303 => "00000010001011110001010011010001",
			1304 => "00000000000000000001010011010001",
			1305 => "0000000001000000000010001100011000",
			1306 => "0000001111000000000010001000001100",
			1307 => "0000001111000000001011011100001000",
			1308 => "0000001111000000001011011100000100",
			1309 => "11111111010110100001010011010001",
			1310 => "00000000001010010001010011010001",
			1311 => "11111110001010100001010011010001",
			1312 => "0000000101000000001110110000001000",
			1313 => "0000000111000000001000111000000100",
			1314 => "00000001000110100001010011010001",
			1315 => "00000010011000010001010011010001",
			1316 => "00000000000000000001010011010001",
			1317 => "0000000001000000001001111000010000",
			1318 => "0000001100000000001000111000001000",
			1319 => "0000000001000000000010001100000100",
			1320 => "11111111100101110001010011010001",
			1321 => "11111110010110000001010011010001",
			1322 => "0000001110000000000001111100000100",
			1323 => "11111111100101100001010011010001",
			1324 => "00000001100100010001010011010001",
			1325 => "0000001010000000000001010000001000",
			1326 => "0000001110000000000101100100000100",
			1327 => "11111110110110010001010011010001",
			1328 => "00000000000000000001010011010001",
			1329 => "0000001101000000001000000000000100",
			1330 => "00000001001111010001010011010001",
			1331 => "11111111110100110001010011010001",
			1332 => "0000000000000000001100001010110000",
			1333 => "0000001010000000001100011101010100",
			1334 => "0000000010000000000010110100101000",
			1335 => "0000000010000000000001001000010100",
			1336 => "0000000000000000001000110000001100",
			1337 => "0000001011000000001011000100000100",
			1338 => "11111110000100100001011011110101",
			1339 => "0000001100000000000100010100000100",
			1340 => "00000000111110010001011011110101",
			1341 => "11111110100101110001011011110101",
			1342 => "0000001100000000001010000000000100",
			1343 => "00000000000000000001011011110101",
			1344 => "00000001101000100001011011110101",
			1345 => "0000001000000000000001110100010000",
			1346 => "0000001010000000001000010100001000",
			1347 => "0000000010000000001110101100000100",
			1348 => "11111111101001100001011011110101",
			1349 => "11111101111101000001011011110101",
			1350 => "0000001010000000001001000100000100",
			1351 => "00000001010111000001011011110101",
			1352 => "11111111100011110001011011110101",
			1353 => "11111101101101100001011011110101",
			1354 => "0000001000000000000010101000100000",
			1355 => "0000000100000000000010100100010000",
			1356 => "0000000011000000001000111100001000",
			1357 => "0000001011000000000100010100000100",
			1358 => "11111111111001110001011011110101",
			1359 => "00000000011100110001011011110101",
			1360 => "0000001101000000001100101100000100",
			1361 => "11111111101111000001011011110101",
			1362 => "00000000000101100001011011110101",
			1363 => "0000001101000000000011011100001000",
			1364 => "0000000000000000001011000100000100",
			1365 => "00000000000000000001011011110101",
			1366 => "00000001101101110001011011110101",
			1367 => "0000000110000000000100110100000100",
			1368 => "11111110001111110001011011110101",
			1369 => "11111111111011110001011011110101",
			1370 => "0000001101000000000011011100000100",
			1371 => "11111111100000100001011011110101",
			1372 => "0000000011000000001000111000000100",
			1373 => "00000001000000100001011011110101",
			1374 => "00000010000010010001011011110101",
			1375 => "0000001001000000000111100100101100",
			1376 => "0000000011000000000101101100011000",
			1377 => "0000001001000000000110101000010000",
			1378 => "0000000100000000000011110100001000",
			1379 => "0000000000000000001011000100000100",
			1380 => "11111101111010010001011011110101",
			1381 => "11111111110101000001011011110101",
			1382 => "0000001100000000000100010100000100",
			1383 => "00000001000011110001011011110101",
			1384 => "11111111000111000001011011110101",
			1385 => "0000001001000000000111100100000100",
			1386 => "00000001100100000001011011110101",
			1387 => "00000000000101100001011011110101",
			1388 => "0000001110000000000000101000001000",
			1389 => "0000001110000000001011000100000100",
			1390 => "11111111100000000001011011110101",
			1391 => "11111100110010000001011011110101",
			1392 => "0000001110000000000100000000000100",
			1393 => "00000001101001000001011011110101",
			1394 => "0000001010000000000110011100000100",
			1395 => "11111110101011000001011011110101",
			1396 => "00000000110110100001011011110101",
			1397 => "0000000110000000001101011000011000",
			1398 => "0000000011000000000001111100001100",
			1399 => "0000001110000000001100110000001000",
			1400 => "0000001100000000000000101000000100",
			1401 => "00000001100110110001011011110101",
			1402 => "11111111110011000001011011110101",
			1403 => "11111110000001010001011011110101",
			1404 => "0000001111000000001101000100000100",
			1405 => "00000001111010110001011011110101",
			1406 => "0000001101000000000001111100000100",
			1407 => "00000001011111010001011011110101",
			1408 => "11111111101001000001011011110101",
			1409 => "0000000111000000001000111000001100",
			1410 => "0000000011000000001010111100000100",
			1411 => "00000000111110000001011011110101",
			1412 => "0000001101000000001010111100000100",
			1413 => "11111110000001010001011011110101",
			1414 => "11111111010101010001011011110101",
			1415 => "0000001101000000000111001000000100",
			1416 => "00000001011101010001011011110101",
			1417 => "0000000100000000000010100100000100",
			1418 => "11111111010010000001011011110101",
			1419 => "00000000010100110001011011110101",
			1420 => "0000001100000000000111111000101100",
			1421 => "0000000011000000000100000000101000",
			1422 => "0000000011000000000100010100011100",
			1423 => "0000001010000000000110011100001100",
			1424 => "0000001100000000000000111000000100",
			1425 => "00000000000000000001011011110101",
			1426 => "0000000110000000001101111100000100",
			1427 => "00000000000000000001011011110101",
			1428 => "00000001100101110001011011110101",
			1429 => "0000001101000000001000111100001000",
			1430 => "0000001100000000001010000000000100",
			1431 => "11111111111111010001011011110101",
			1432 => "11111101011000000001011011110101",
			1433 => "0000000011000000000000111000000100",
			1434 => "00000001000000010001011011110101",
			1435 => "11111111011010000001011011110101",
			1436 => "0000000000000000000100000000000100",
			1437 => "00000000000000000001011011110101",
			1438 => "0000001101000000001000111000000100",
			1439 => "00000000011111110001011011110101",
			1440 => "11111101101010000001011011110101",
			1441 => "00000001101011010001011011110101",
			1442 => "0000000111000000000100010100010000",
			1443 => "0000001001000000001100110100001100",
			1444 => "0000001111000000000100011000001000",
			1445 => "0000001001000000000000011000000100",
			1446 => "00000000000000000001011011110101",
			1447 => "00000001011110110001011011110101",
			1448 => "11111110010101100001011011110101",
			1449 => "00000001100110010001011011110101",
			1450 => "0000001011000000000000101000010100",
			1451 => "0000001001000000000110101000001100",
			1452 => "0000000100000000000011011000000100",
			1453 => "00000001100010010001011011110101",
			1454 => "0000000110000000000100110100000100",
			1455 => "00000001000011010001011011110101",
			1456 => "11111111001101110001011011110101",
			1457 => "0000000010000000000011001000000100",
			1458 => "11111101001000110001011011110101",
			1459 => "00000000000000000001011011110101",
			1460 => "0000001101000000001110001100000100",
			1461 => "00000001101000100001011011110101",
			1462 => "0000001001000000000110101000001000",
			1463 => "0000000110000000001101111100000100",
			1464 => "00000000000100100001011011110101",
			1465 => "11111110100011100001011011110101",
			1466 => "0000001000000000000111000000000100",
			1467 => "00000000000000000001011011110101",
			1468 => "00000001000100010001011011110101",
			1469 => "0000001110000000000101101110011000",
			1470 => "0000001111000000000101100101011100",
			1471 => "0000000110000000000111101000101000",
			1472 => "0000001101000000000110000100011000",
			1473 => "0000000011000000001000111000010000",
			1474 => "0000000000000000000011111100001000",
			1475 => "0000001000000000000101000100000100",
			1476 => "11111101111001000001100101010001",
			1477 => "00000001011010010001100101010001",
			1478 => "0000000111000000000100010100000100",
			1479 => "11111111001111110001100101010001",
			1480 => "00000001100100110001100101010001",
			1481 => "0000001110000000001110111100000100",
			1482 => "11111110110100010001100101010001",
			1483 => "11111101011011010001100101010001",
			1484 => "0000000101000000000101101100000100",
			1485 => "00000000000110010001100101010001",
			1486 => "0000000000000000001001101000000100",
			1487 => "00000000000000000001100101010001",
			1488 => "0000001000000000001100000100000100",
			1489 => "00000001101111010001100101010001",
			1490 => "00000000100011000001100101010001",
			1491 => "0000000011000000001100110000100000",
			1492 => "0000001011000000001100001000010000",
			1493 => "0000000101000000001101100000001000",
			1494 => "0000001011000000000100010100000100",
			1495 => "11111111110011000001100101010001",
			1496 => "00000000110000010001100101010001",
			1497 => "0000000101000000001101100000000100",
			1498 => "11111110110111110001100101010001",
			1499 => "11111111101100100001100101010001",
			1500 => "0000001111000000000100000100001000",
			1501 => "0000000000000000000011010000000100",
			1502 => "11111110111101010001100101010001",
			1503 => "00000000010111010001100101010001",
			1504 => "0000000001000000001110100000000100",
			1505 => "00000000010001100001100101010001",
			1506 => "00000001100011110001100101010001",
			1507 => "0000000010000000001111010000010000",
			1508 => "0000000010000000000111100000001000",
			1509 => "0000000010000000001101000100000100",
			1510 => "11111110110011000001100101010001",
			1511 => "00000000000000000001100101010001",
			1512 => "0000000101000000001110001100000100",
			1513 => "11111101010110110001100101010001",
			1514 => "11111110100000100001100101010001",
			1515 => "00000000111101010001100101010001",
			1516 => "0000001000000000000111000000101100",
			1517 => "0000000100000000000011011000011100",
			1518 => "0000001101000000000011011100001100",
			1519 => "0000000100000000001001001100000100",
			1520 => "11111100111010110001100101010001",
			1521 => "0000000100000000000011010100000100",
			1522 => "00000001000010010001100101010001",
			1523 => "11111110101101000001100101010001",
			1524 => "0000000011000000001001110000001000",
			1525 => "0000000000000000000000101000000100",
			1526 => "00000000111000000001100101010001",
			1527 => "11111111100010000001100101010001",
			1528 => "0000000000000000000000110000000100",
			1529 => "00000000010001010001100101010001",
			1530 => "11111111111100100001100101010001",
			1531 => "0000001111000000001010010100001000",
			1532 => "0000000111000000000111111000000100",
			1533 => "00000000000000000001100101010001",
			1534 => "11111100110010000001100101010001",
			1535 => "0000001000000000000001110100000100",
			1536 => "00000000000000000001100101010001",
			1537 => "00000001010111000001100101010001",
			1538 => "0000000100000000000001001100001000",
			1539 => "0000000010000000000010000100000100",
			1540 => "00000001101011110001100101010001",
			1541 => "00000000101011110001100101010001",
			1542 => "0000000101000000001101111000000100",
			1543 => "00000000000000000001100101010001",
			1544 => "11111110010101000001100101010001",
			1545 => "0000000011000000000111001001001000",
			1546 => "0000001100000000000000101000100000",
			1547 => "0000001100000000000100010100010000",
			1548 => "0000001111000000001110101000001100",
			1549 => "0000000100000000001100111000000100",
			1550 => "00000110011111110001100101010001",
			1551 => "0000001111000000001101000100000100",
			1552 => "11111111011001110001100101010001",
			1553 => "11111101011011110001100101010001",
			1554 => "00000001111101110001100101010001",
			1555 => "0000001100000000000100010100001000",
			1556 => "0000000100000000001100001100000100",
			1557 => "11111111010100010001100101010001",
			1558 => "11111101100011000001100101010001",
			1559 => "0000001111000000001110101100000100",
			1560 => "11111110001111100001100101010001",
			1561 => "11111111111010100001100101010001",
			1562 => "0000001011000000001000111100010100",
			1563 => "0000001000000000001001101000000100",
			1564 => "11111110011010000001100101010001",
			1565 => "0000001110000000001100101100001000",
			1566 => "0000001000000000000110001000000100",
			1567 => "00000001001000110001100101010001",
			1568 => "11111111001111010001100101010001",
			1569 => "0000001100000000000000101000000100",
			1570 => "11111111110110110001100101010001",
			1571 => "00000010110100010001100101010001",
			1572 => "0000000010000000001100100100001000",
			1573 => "0000000110000000001101011100000100",
			1574 => "00000000000000000001100101010001",
			1575 => "00000011110010110001100101010001",
			1576 => "0000001100000000000000101000000100",
			1577 => "00000000111000010001100101010001",
			1578 => "0000001110000000000000001100000100",
			1579 => "11111111011100110001100101010001",
			1580 => "11111101101011010001100101010001",
			1581 => "0000000011000000000111001000010100",
			1582 => "0000000000000000001010000000001100",
			1583 => "0000001101000000000001111100000100",
			1584 => "00000011001111000001100101010001",
			1585 => "0000000100000000000010110000000100",
			1586 => "11111111011101110001100101010001",
			1587 => "00000010011001000001100101010001",
			1588 => "0000001111000000000010110100000100",
			1589 => "11111110101000000001100101010001",
			1590 => "00000001111000000001100101010001",
			1591 => "0000000110000000001010011000100000",
			1592 => "0000000010000000000010000100010000",
			1593 => "0000000100000000001110111000001000",
			1594 => "0000000110000000000100110100000100",
			1595 => "00000000011011000001100101010001",
			1596 => "11111111100110010001100101010001",
			1597 => "0000000100000000000011010100000100",
			1598 => "00000001001110110001100101010001",
			1599 => "11111111001011110001100101010001",
			1600 => "0000000111000000000100000000001000",
			1601 => "0000001101000000000100001000000100",
			1602 => "00000000101000110001100101010001",
			1603 => "00000010100001110001100101010001",
			1604 => "0000000110000000001010011000000100",
			1605 => "11111111111001000001100101010001",
			1606 => "00000001100001100001100101010001",
			1607 => "0000000101000000000100001000001100",
			1608 => "0000000010000000000110111100001000",
			1609 => "0000001110000000001010111100000100",
			1610 => "11111110000101010001100101010001",
			1611 => "11111111101101010001100101010001",
			1612 => "00000000101000100001100101010001",
			1613 => "0000001111000000000001000000001000",
			1614 => "0000000010000000000010000100000100",
			1615 => "00000000000110010001100101010001",
			1616 => "00000001100010100001100101010001",
			1617 => "0000001110000000000100000100000100",
			1618 => "11111111001000110001100101010001",
			1619 => "00000000000000110001100101010001",
			1620 => "0000001101000000001011000010111100",
			1621 => "0000001111000000000101100101000100",
			1622 => "0000001110000000000100000000110100",
			1623 => "0000000100000000000110110000100000",
			1624 => "0000000011000000000000110000010000",
			1625 => "0000000111000000000111111000001000",
			1626 => "0000000011000000000011111100000100",
			1627 => "00000001011010000001101101010101",
			1628 => "11111111101110100001101101010101",
			1629 => "0000001111000000001010111000000100",
			1630 => "00000000111011100001101101010101",
			1631 => "00000001110111000001101101010101",
			1632 => "0000000111000000001100001000001000",
			1633 => "0000001100000000000100010100000100",
			1634 => "00000000000000010001101101010101",
			1635 => "11111111010011110001101101010101",
			1636 => "0000000111000000001100001000000100",
			1637 => "00000001100100110001101101010101",
			1638 => "00000000000101000001101101010101",
			1639 => "0000000110000000001010011000001100",
			1640 => "0000000100000000000011111000000100",
			1641 => "11111101101000000001101101010101",
			1642 => "0000000100000000000101100000000100",
			1643 => "00000000010110100001101101010101",
			1644 => "11111110011011010001101101010101",
			1645 => "0000001010000000001000110000000100",
			1646 => "00000001010010100001101101010101",
			1647 => "00000000000000000001101101010101",
			1648 => "0000000110000000000111101000001000",
			1649 => "0000000010000000000001001000000100",
			1650 => "11111101111011010001101101010101",
			1651 => "00000001100000010001101101010101",
			1652 => "0000001100000000000100010100000100",
			1653 => "11111111111000010001101101010101",
			1654 => "11111101101111010001101101010101",
			1655 => "0000001010000000000110011000111100",
			1656 => "0000000010000000000100101000100000",
			1657 => "0000000011000000000110000100010000",
			1658 => "0000001001000000000110101000001000",
			1659 => "0000000011000000001101100000000100",
			1660 => "00000000100010100001101101010101",
			1661 => "11111110011000100001101101010101",
			1662 => "0000001100000000000111111000000100",
			1663 => "00000011000111110001101101010101",
			1664 => "00000001001110010001101101010101",
			1665 => "0000001001000000000110101000001000",
			1666 => "0000001111000000000101110100000100",
			1667 => "11111101110101000001101101010101",
			1668 => "11111111110111000001101101010101",
			1669 => "0000001010000000001000010100000100",
			1670 => "00000000101000010001101101010101",
			1671 => "11111111110011000001101101010101",
			1672 => "0000000010000000000100101000001100",
			1673 => "0000000011000000000100001000001000",
			1674 => "0000000100000000001000001000000100",
			1675 => "00000100010101000001101101010101",
			1676 => "00000001100110010001101101010101",
			1677 => "00000000011011010001101101010101",
			1678 => "0000000110000000000001111000001000",
			1679 => "0000001110000000001001110000000100",
			1680 => "00000000000000000001101101010101",
			1681 => "11111110011011010001101101010101",
			1682 => "0000001100000000001000111100000100",
			1683 => "00000000111111010001101101010101",
			1684 => "11111110110111010001101101010101",
			1685 => "0000001110000000000100010100011100",
			1686 => "0000001100000000001110111100010000",
			1687 => "0000000110000000000100110100001000",
			1688 => "0000001111000000000110110100000100",
			1689 => "00000000101010000001101101010101",
			1690 => "11111110010101100001101101010101",
			1691 => "0000000010000000000011001000000100",
			1692 => "00000001100100010001101101010101",
			1693 => "11111111000100100001101101010101",
			1694 => "0000000000000000000000111000000100",
			1695 => "11111111001101110001101101010101",
			1696 => "0000001010000000000001010000000100",
			1697 => "00000001101000110001101101010101",
			1698 => "00000000101011110001101101010101",
			1699 => "0000001001000000000110101000010000",
			1700 => "0000001111000000000111110000001000",
			1701 => "0000000011000000001101100000000100",
			1702 => "00000000011011100001101101010101",
			1703 => "11111110011111010001101101010101",
			1704 => "0000001010000000000001010000000100",
			1705 => "00000001011001110001101101010101",
			1706 => "11111111100111010001101101010101",
			1707 => "0000001110000000001100001000001000",
			1708 => "0000000110000000000100110100000100",
			1709 => "00000010010000010001101101010101",
			1710 => "00000000111000000001101101010101",
			1711 => "0000000100000000000011010100000100",
			1712 => "00000000000000010001101101010101",
			1713 => "00000000101100000001101101010101",
			1714 => "0000000000000000000111000000010100",
			1715 => "0000001011000000000000001100010000",
			1716 => "0000001000000000001100011100001100",
			1717 => "0000000111000000000101101100000100",
			1718 => "11111110011010110001101101010101",
			1719 => "0000000111000000000101101100000100",
			1720 => "00000000101011100001101101010101",
			1721 => "11111111000100100001101101010101",
			1722 => "00000000011001000001101101010101",
			1723 => "11111110011000000001101101010101",
			1724 => "0000000100000000000000000000110000",
			1725 => "0000001001000000001101011100010100",
			1726 => "0000001100000000001000111000001100",
			1727 => "0000001101000000001000000000000100",
			1728 => "11111111100110000001101101010101",
			1729 => "0000000111000000001101100000000100",
			1730 => "11111110111011000001101101010101",
			1731 => "11111101001000000001101101010101",
			1732 => "0000000110000000001101011000000100",
			1733 => "11111111010001110001101101010101",
			1734 => "00000001110010010001101101010101",
			1735 => "0000000111000000001101100000001100",
			1736 => "0000001110000000000001101000000100",
			1737 => "00000001111111000001101101010101",
			1738 => "0000000100000000000011110000000100",
			1739 => "11111101110010010001101101010101",
			1740 => "11111111101101100001101101010101",
			1741 => "0000001110000000000011100000001000",
			1742 => "0000001010000000001010110000000100",
			1743 => "11111101001001100001101101010101",
			1744 => "00000000000000000001101101010101",
			1745 => "0000001101000000001001001000000100",
			1746 => "00000001110110010001101101010101",
			1747 => "00000000000000100001101101010101",
			1748 => "11111110011011000001101101010101",
			1749 => "0000001100000000000111111010001000",
			1750 => "0000001001000000000110101001001100",
			1751 => "0000000011000000001001110000110000",
			1752 => "0000000111000000001011000100100000",
			1753 => "0000000000000000000010111100010000",
			1754 => "0000000101000000000011011100001000",
			1755 => "0000000100000000000101000000000100",
			1756 => "11111110101110010001110110110001",
			1757 => "11111010110111110001110110110001",
			1758 => "0000001100000000000111111000000100",
			1759 => "00000001101000100001110110110001",
			1760 => "11111111111001110001110110110001",
			1761 => "0000000001000000000110000000001000",
			1762 => "0000000011000000000011010000000100",
			1763 => "00000000111100110001110110110001",
			1764 => "11111111000001010001110110110001",
			1765 => "0000000011000000001011000100000100",
			1766 => "00000000110001000001110110110001",
			1767 => "11111111111101100001110110110001",
			1768 => "0000001100000000000111111000000100",
			1769 => "00000001110010100001110110110001",
			1770 => "0000000110000000001101111100001000",
			1771 => "0000000110000000000001111000000100",
			1772 => "00000001001011100001110110110001",
			1773 => "11111111000100100001110110110001",
			1774 => "00000001101110100001110110110001",
			1775 => "0000001000000000000010101000011000",
			1776 => "0000001110000000000111111000001100",
			1777 => "0000001100000000000111111000001000",
			1778 => "0000000010000000000011001000000100",
			1779 => "11111111110000000001110110110001",
			1780 => "11111101010100010001110110110001",
			1781 => "11111101010101000001110110110001",
			1782 => "0000000100000000001111100000001000",
			1783 => "0000000000000000000011010000000100",
			1784 => "11111101001011010001110110110001",
			1785 => "11111111111110100001110110110001",
			1786 => "11111101000110000001110110110001",
			1787 => "00000001011001110001110110110001",
			1788 => "0000000101000000001100110000010100",
			1789 => "0000001011000000000000101000010000",
			1790 => "0000001110000000001000111100001100",
			1791 => "0000001110000000001110111100000100",
			1792 => "11111111111100100001110110110001",
			1793 => "0000000110000000001101111100000100",
			1794 => "00000001000000100001110110110001",
			1795 => "00000010010001010001110110110001",
			1796 => "11111111101110010001110110110001",
			1797 => "00000011001010010001110110110001",
			1798 => "0000001100000000001110111100010000",
			1799 => "0000001010000000001001000100000100",
			1800 => "00000001001111010001110110110001",
			1801 => "0000001100000000001010000000000100",
			1802 => "00000000001101010001110110110001",
			1803 => "0000000011000000000110000100000100",
			1804 => "11111101001001110001110110110001",
			1805 => "11111110101111000001110110110001",
			1806 => "0000000111000000001100001000010000",
			1807 => "0000001110000000001001110000001000",
			1808 => "0000001001000000000111100100000100",
			1809 => "00000000101100110001110110110001",
			1810 => "00000010111000110001110110110001",
			1811 => "0000000011000000000100001000000100",
			1812 => "11111111011001010001110110110001",
			1813 => "00000001000100000001110110110001",
			1814 => "0000000101000000001110001100000100",
			1815 => "11111101101001110001110110110001",
			1816 => "00000000000000000001110110110001",
			1817 => "0000001100000000000100010100110100",
			1818 => "0000001010000000001001000100010100",
			1819 => "0000000111000000000100010100000100",
			1820 => "11111101111001100001110110110001",
			1821 => "0000000001000000001110100000001000",
			1822 => "0000000110000000000001111000000100",
			1823 => "00000000010000100001110110110001",
			1824 => "00000010100101110001110110110001",
			1825 => "0000001100000000000111111000000100",
			1826 => "00000000000001010001110110110001",
			1827 => "11111101110011000001110110110001",
			1828 => "0000000010000000000011001000011000",
			1829 => "0000000111000000000100010100001100",
			1830 => "0000001011000000001110111100000100",
			1831 => "00000001111001000001110110110001",
			1832 => "0000000011000000000000110000000100",
			1833 => "11111110000110100001110110110001",
			1834 => "00000000111000000001110110110001",
			1835 => "0000000001000000000110000000000100",
			1836 => "00000001000111010001110110110001",
			1837 => "0000001110000000000100010100000100",
			1838 => "11111110001110100001110110110001",
			1839 => "11111101010100100001110110110001",
			1840 => "0000000110000000001100011000000100",
			1841 => "00000001000011110001110110110001",
			1842 => "11111110100110100001110110110001",
			1843 => "0000000011000000001100110000111000",
			1844 => "0000001001000000000110101000011100",
			1845 => "0000000001000000001110100000010000",
			1846 => "0000000101000000000101101100001000",
			1847 => "0000000011000000000011011100000100",
			1848 => "00000000001000000001110110110001",
			1849 => "11111110111111010001110110110001",
			1850 => "0000000010000000000111100000000100",
			1851 => "11111111110100100001110110110001",
			1852 => "00000000111100110001110110110001",
			1853 => "0000000110000000001100011000001000",
			1854 => "0000000111000000001100001000000100",
			1855 => "00000000001100110001110110110001",
			1856 => "11111110100101100001110110110001",
			1857 => "00000001110011000001110110110001",
			1858 => "0000001000000000001011010100001100",
			1859 => "0000000100000000001100001100001000",
			1860 => "0000000010000000000110100000000100",
			1861 => "00000000000100110001110110110001",
			1862 => "00000001111100000001110110110001",
			1863 => "11111110010010010001110110110001",
			1864 => "0000000100000000001110111000001000",
			1865 => "0000000100000000000010111000000100",
			1866 => "00000010111010110001110110110001",
			1867 => "00000001110010000001110110110001",
			1868 => "0000000110000000001010011000000100",
			1869 => "11111111111001000001110110110001",
			1870 => "00000001100110110001110110110001",
			1871 => "0000001001000000000111100100011100",
			1872 => "0000000011000000001101111000010000",
			1873 => "0000000010000000001100010100001000",
			1874 => "0000000011000000001100110000000100",
			1875 => "11111110010010110001110110110001",
			1876 => "11111111101001110001110110110001",
			1877 => "0000001010000000000110011100000100",
			1878 => "00000001111000000001110110110001",
			1879 => "11111111100110000001110110110001",
			1880 => "0000000100000000001011100000001000",
			1881 => "0000001010000000001100011100000100",
			1882 => "11111110110100010001110110110001",
			1883 => "11111100000010110001110110110001",
			1884 => "00000001100110110001110110110001",
			1885 => "0000000001000000001100110100010000",
			1886 => "0000000011000000000000001100001000",
			1887 => "0000000010000000001001010000000100",
			1888 => "00000000000000000001110110110001",
			1889 => "00000001011100000001110110110001",
			1890 => "0000001011000000001100001000000100",
			1891 => "00000001010111110001110110110001",
			1892 => "11111111000110000001110110110001",
			1893 => "0000001001000000000111100100001000",
			1894 => "0000001000000000000111000100000100",
			1895 => "11111111001101100001110110110001",
			1896 => "00000000010111100001110110110001",
			1897 => "0000001011000000000100000000000100",
			1898 => "00000001000110110001110110110001",
			1899 => "00000000000101000001110110110001",
			1900 => "0000001110000000000101101110100000",
			1901 => "0000001111000000000101100101011100",
			1902 => "0000000110000000000111101000101000",
			1903 => "0000001101000000000110000100011000",
			1904 => "0000000011000000001000111000010000",
			1905 => "0000000101000000001000111000001000",
			1906 => "0000001111000000001011000000000100",
			1907 => "00000000000001010010000000010101",
			1908 => "11111100111000100010000000010101",
			1909 => "0000001010000000001001000100000100",
			1910 => "00000000111110000010000000010101",
			1911 => "11111110111011000010000000010101",
			1912 => "0000000000000000001101010000000100",
			1913 => "11111100100110010010000000010101",
			1914 => "11111110000111110010000000010101",
			1915 => "0000000101000000000101101100000100",
			1916 => "00000000000000000010000000010101",
			1917 => "0000000000000000001001101000000100",
			1918 => "11111111111101100010000000010101",
			1919 => "0000001111000000000000011100000100",
			1920 => "00000001110010100010000000010101",
			1921 => "00000000111010000010000000010101",
			1922 => "0000000011000000001100110000100000",
			1923 => "0000001011000000001100001000010000",
			1924 => "0000000101000000001101100000001000",
			1925 => "0000000101000000000011011100000100",
			1926 => "11111111110111100010000000010101",
			1927 => "00000001000001010010000000010101",
			1928 => "0000001110000000001011000100000100",
			1929 => "11111111011001100010000000010101",
			1930 => "00000001001000110010000000010101",
			1931 => "0000001111000000000111010000001000",
			1932 => "0000000011000000001001110000000100",
			1933 => "00000000000100010010000000010101",
			1934 => "11111101011111100010000000010101",
			1935 => "0000000011000000001001110000000100",
			1936 => "00000001101010110010000000010101",
			1937 => "00000000011100010010000000010101",
			1938 => "0000001101000000001101010100010000",
			1939 => "0000000001000000001100110100001000",
			1940 => "0000001101000000001100101000000100",
			1941 => "11111110111110010010000000010101",
			1942 => "00000000101010000010000000010101",
			1943 => "0000000001000000000010001100000100",
			1944 => "11111110010111110010000000010101",
			1945 => "11111101010011100010000000010101",
			1946 => "00000000101010000010000000010101",
			1947 => "0000001001000000001011101000101100",
			1948 => "0000001011000000001101100000100000",
			1949 => "0000000011000000001001110000010000",
			1950 => "0000001101000000000011011100001000",
			1951 => "0000001111000000000101110100000100",
			1952 => "11111110111000010010000000010101",
			1953 => "00000001101010110010000000010101",
			1954 => "0000000000000000000000101000000100",
			1955 => "00000001000010110010000000010101",
			1956 => "11111111100000000010000000010101",
			1957 => "0000001001000000001001111000001000",
			1958 => "0000001011000000000000101000000100",
			1959 => "11111101111100000010000000010101",
			1960 => "00000001001001010010000000010101",
			1961 => "0000001001000000000110101000000100",
			1962 => "11111111111110110010000000010101",
			1963 => "00000000010110000010000000010101",
			1964 => "0000000111000000001001110000000100",
			1965 => "11111100101111010010000000010101",
			1966 => "0000000101000000000000011100000100",
			1967 => "00000001010000000010000000010101",
			1968 => "00000000000000000010000000010101",
			1969 => "0000000110000000001010011000001000",
			1970 => "0000001110000000001100110000000100",
			1971 => "00000010110100000010000000010101",
			1972 => "00000001000011100010000000010101",
			1973 => "0000001111000000000000110100001000",
			1974 => "0000000011000000001010111100000100",
			1975 => "00000001100100000010000000010101",
			1976 => "00000000000010000010000000010101",
			1977 => "0000000010000000001011101100000100",
			1978 => "11111100001101010010000000010101",
			1979 => "00000000000000000010000000010101",
			1980 => "0000000000000000001111000100111000",
			1981 => "0000001001000000000100110100110000",
			1982 => "0000000100000000001000000100011100",
			1983 => "0000000000000000001101010000001100",
			1984 => "0000000100000000001011110000001000",
			1985 => "0000000110000000001010011000000100",
			1986 => "11111111111101110010000000010101",
			1987 => "00000001101111010010000000010101",
			1988 => "00000010010111100010000000010101",
			1989 => "0000001010000000001001000100001000",
			1990 => "0000000101000000001100101000000100",
			1991 => "11111111011100100010000000010101",
			1992 => "11111110000001000010000000010101",
			1993 => "0000000110000000001001100100000100",
			1994 => "00000001010000100010000000010101",
			1995 => "11111111100110010010000000010101",
			1996 => "0000000110000000001101111100000100",
			1997 => "11111101100101000010000000010101",
			1998 => "0000000010000000001100010100001000",
			1999 => "0000000010000000000100101000000100",
			2000 => "00000001101011000010000000010101",
			2001 => "00000011010001100010000000010101",
			2002 => "0000001110000000000101100100000100",
			2003 => "11111111111100110010000000010101",
			2004 => "00000001001010110010000000010101",
			2005 => "0000001010000000001010110000000100",
			2006 => "11111110011100000010000000010101",
			2007 => "00000000010110010010000000010101",
			2008 => "0000000010000000001110010000100000",
			2009 => "0000000011000000000000001100000100",
			2010 => "00000010110011100010000000010101",
			2011 => "0000000110000000001010011000010000",
			2012 => "0000001101000000000001111100001000",
			2013 => "0000001101000000001100101000000100",
			2014 => "11111110001110100010000000010101",
			2015 => "00000000011011000010000000010101",
			2016 => "0000001010000000000001010000000100",
			2017 => "11111110000010010010000000010101",
			2018 => "11111111110010000010000000010101",
			2019 => "0000001001000000001101101000000100",
			2020 => "00000010110010010010000000010101",
			2021 => "0000001001000000001011101000000100",
			2022 => "11111101100111100010000000010101",
			2023 => "00000000011011100010000000010101",
			2024 => "0000000110000000001100011000011100",
			2025 => "0000001111000000000010110100001100",
			2026 => "0000001011000000001000111100000100",
			2027 => "11111110001110110010000000010101",
			2028 => "0000001111000000001110101100000100",
			2029 => "00000001011111100010000000010101",
			2030 => "11111111110001110010000000010101",
			2031 => "0000001110000000001110001100001000",
			2032 => "0000001010000000000001010000000100",
			2033 => "00000010101010000010000000010101",
			2034 => "00000000010011100010000000010101",
			2035 => "0000000010000000000110010000000100",
			2036 => "11111111110100010010000000010101",
			2037 => "00000001111000100010000000010101",
			2038 => "0000001001000000001011101000010000",
			2039 => "0000001111000000001110101100001000",
			2040 => "0000000100000000001010110100000100",
			2041 => "11111111011011100010000000010101",
			2042 => "00000001010101110010000000010101",
			2043 => "0000000101000000000111001000000100",
			2044 => "11111111001111110010000000010101",
			2045 => "00000001001110110010000000010101",
			2046 => "0000000011000000001011000000001000",
			2047 => "0000000010000000001100010100000100",
			2048 => "00000000011111000010000000010101",
			2049 => "00000010011011000010000000010101",
			2050 => "0000000100000000000101000000000100",
			2051 => "11111110111000110010000000010101",
			2052 => "11111111110111110010000000010101",
			2053 => "0000001000000000001001101010110000",
			2054 => "0000001000000000001001101001011100",
			2055 => "0000001101000000000101101100101000",
			2056 => "0000000111000000000100010100011000",
			2057 => "0000000011000000001000111000010000",
			2058 => "0000000000000000000011111100001000",
			2059 => "0000001011000000000100010100000100",
			2060 => "11111111011101110010001010011001",
			2061 => "00000001101000010010001010011001",
			2062 => "0000001111000000000000011100000100",
			2063 => "11111101101010010010001010011001",
			2064 => "00000001010011010010001010011001",
			2065 => "0000000000000000000011111100000100",
			2066 => "11111101110011100010001010011001",
			2067 => "00000000110110000010001010011001",
			2068 => "0000000010000000001101000100001100",
			2069 => "0000000011000000000100010100000100",
			2070 => "00000000000000000010001010011001",
			2071 => "0000001101000000001100110000000100",
			2072 => "11111100000100110010001010011001",
			2073 => "11111101111100000010001010011001",
			2074 => "00000000100011010010001010011001",
			2075 => "0000000001000000000010001100011100",
			2076 => "0000001011000000001001110000010000",
			2077 => "0000000111000000000100010100001000",
			2078 => "0000000001000000001110100000000100",
			2079 => "00000000101010010010001010011001",
			2080 => "11111101010011110010001010011001",
			2081 => "0000001011000000000000101000000100",
			2082 => "00000001010110010010001010011001",
			2083 => "00000000000011010010001010011001",
			2084 => "0000000010000000001110101000000100",
			2085 => "11111110111100010010001010011001",
			2086 => "0000000100000000001110100100000100",
			2087 => "00000010100101010010001010011001",
			2088 => "00000000110000010010001010011001",
			2089 => "0000001101000000000001111100001000",
			2090 => "0000000101000000000000001100000100",
			2091 => "11111111110010010010001010011001",
			2092 => "11111101011001000010001010011001",
			2093 => "0000000100000000000110001100001000",
			2094 => "0000000000000000001111000100000100",
			2095 => "11111111111111100010001010011001",
			2096 => "11111110010110110010001010011001",
			2097 => "0000001100000000000110000100000100",
			2098 => "00000010101100000010001010011001",
			2099 => "11111110110011010010001010011001",
			2100 => "0000000010000000000101110000110000",
			2101 => "0000000001000000001100110100100000",
			2102 => "0000001111000000000100000100010000",
			2103 => "0000001111000000001111011100001000",
			2104 => "0000000101000000001100110000000100",
			2105 => "00000001101000010010001010011001",
			2106 => "11111111010000100010001010011001",
			2107 => "0000000101000000001101100000000100",
			2108 => "00000000000000000010001010011001",
			2109 => "11111101110000110010001010011001",
			2110 => "0000000011000000001101100000001000",
			2111 => "0000000110000000000001111000000100",
			2112 => "00000000000111000010001010011001",
			2113 => "00000010000010000010001010011001",
			2114 => "0000000111000000001100001000000100",
			2115 => "11111111110011100010001010011001",
			2116 => "00000010000010110010001010011001",
			2117 => "0000001001000000001101101000001100",
			2118 => "0000001000000000001001101000000100",
			2119 => "11111111011010000010001010011001",
			2120 => "0000000011000000001110001100000100",
			2121 => "11111100111010000010001010011001",
			2122 => "11111110011010100010001010011001",
			2123 => "00000001010010000010001010011001",
			2124 => "0000000001000000001001111000010100",
			2125 => "0000000011000000001011000000010000",
			2126 => "0000000001000000000010001100001000",
			2127 => "0000001101000000001100101000000100",
			2128 => "00000000111100010010001010011001",
			2129 => "00000010010110110010001010011001",
			2130 => "0000000001000000000010001100000100",
			2131 => "11111110010011110010001010011001",
			2132 => "00000000001100100010001010011001",
			2133 => "00000100001110010010001010011001",
			2134 => "0000000110000000001010011000000100",
			2135 => "11111110000011110010001010011001",
			2136 => "0000001100000000000100000000000100",
			2137 => "00000010101000100010001010011001",
			2138 => "0000000111000000001001110000000100",
			2139 => "11111111010110000010001010011001",
			2140 => "00000000101001100010001010011001",
			2141 => "0000000010000000000111111101001000",
			2142 => "0000001000000000001011010100010100",
			2143 => "0000001111000000001010010100010000",
			2144 => "0000001100000000001010000000000100",
			2145 => "11111101001100110010001010011001",
			2146 => "0000000000000000000011111100000100",
			2147 => "11111110000001000010001010011001",
			2148 => "0000001000000000001001101000000100",
			2149 => "11111101100101000010001010011001",
			2150 => "00000000010011100010001010011001",
			2151 => "00000000110111100010001010011001",
			2152 => "0000001000000000001011010100010100",
			2153 => "0000001100000000000100010100001100",
			2154 => "0000000010000000000001000000000100",
			2155 => "00000000010111010010001010011001",
			2156 => "0000000011000000001101100000000100",
			2157 => "00000001011110000010001010011001",
			2158 => "00000010101111000010001010011001",
			2159 => "0000001101000000001101111000000100",
			2160 => "11111101001100000010001010011001",
			2161 => "00000001010011110010001010011001",
			2162 => "0000000011000000001101111000010000",
			2163 => "0000001101000000000000001100001000",
			2164 => "0000000111000000000100010100000100",
			2165 => "00000000000000100010001010011001",
			2166 => "11111111101001110010001010011001",
			2167 => "0000001100000000000000101000000100",
			2168 => "11111111111111110010001010011001",
			2169 => "00000001101001010010001010011001",
			2170 => "0000001001000000001011101000001000",
			2171 => "0000001000000000001011010100000100",
			2172 => "00000000011110000010001010011001",
			2173 => "11111110100111000010001010011001",
			2174 => "0000000001000000000010001100000100",
			2175 => "00000001100101010010001010011001",
			2176 => "11111111011001100010001010011001",
			2177 => "0000000010000000000111111100001100",
			2178 => "0000000110000000001100011000001000",
			2179 => "0000001011000000001000111100000100",
			2180 => "00000010001011100010001010011001",
			2181 => "11111111110000100010001010011001",
			2182 => "11111110100000000010001010011001",
			2183 => "0000000100000000000100001100100000",
			2184 => "0000001000000000000001110100010000",
			2185 => "0000000111000000000100000000001000",
			2186 => "0000000111000000000100000000000100",
			2187 => "00000000000000000010001010011001",
			2188 => "00000000110011010010001010011001",
			2189 => "0000000101000000000001111100000100",
			2190 => "11111111001000000010001010011001",
			2191 => "11111111111101010010001010011001",
			2192 => "0000001001000000001101101000001000",
			2193 => "0000001001000000000110101000000100",
			2194 => "00000001010000100010001010011001",
			2195 => "11111101111111000010001010011001",
			2196 => "0000001111000000000110100000000100",
			2197 => "00000001010111010010001010011001",
			2198 => "11111111011000110010001010011001",
			2199 => "0000001000000000001111001000010000",
			2200 => "0000001011000000001000111100001000",
			2201 => "0000000000000000001110111100000100",
			2202 => "11110010011000000010001010011001",
			2203 => "00000000000000000010001010011001",
			2204 => "0000001000000000000110001000000100",
			2205 => "11111101101101000010001010011001",
			2206 => "00000000000000000010001010011001",
			2207 => "0000001100000000000111111000001000",
			2208 => "0000001100000000001010000000000100",
			2209 => "00000000000010010010001010011001",
			2210 => "11111110111010010010001010011001",
			2211 => "0000001000000000000010101000000100",
			2212 => "00000000101100010010001010011001",
			2213 => "00000000000110100010001010011001",
			2214 => "0000000010000000000110010010110000",
			2215 => "0000001100000000000100000001100100",
			2216 => "0000001011000000001000111100110000",
			2217 => "0000001101000000000000001100010100",
			2218 => "0000001001000000001101101000010000",
			2219 => "0000001101000000001101111000001000",
			2220 => "0000001100000000000000101000000100",
			2221 => "00000000000001000010010101000101",
			2222 => "11111111001000100010010101000101",
			2223 => "0000001100000000000111111000000100",
			2224 => "00000001110110010010010101000101",
			2225 => "11111111011011100010010101000101",
			2226 => "00000010001001110010010101000101",
			2227 => "0000000101000000001101111000001100",
			2228 => "0000001001000000000111100100000100",
			2229 => "11111111011010110010010101000101",
			2230 => "0000000100000000000011110000000100",
			2231 => "00000000000001000010010101000101",
			2232 => "00000001111111010010010101000101",
			2233 => "0000001011000000000100000000001000",
			2234 => "0000001101000000001100101000000100",
			2235 => "11111101010110110010010101000101",
			2236 => "00000000000000000010010101000101",
			2237 => "0000001110000000001101100000000100",
			2238 => "00000000111011010010010101000101",
			2239 => "11111111111000010010010101000101",
			2240 => "0000001100000000000000101000010100",
			2241 => "0000000110000000000001111000001000",
			2242 => "0000000100000000001011110000000100",
			2243 => "00000000100100100010010101000101",
			2244 => "00000010000100110010010101000101",
			2245 => "0000000100000000000100001100001000",
			2246 => "0000000000000000001110111100000100",
			2247 => "11111110110111100010010101000101",
			2248 => "00000000100010100010010101000101",
			2249 => "11111100100111110010010101000101",
			2250 => "0000001100000000000000101000010000",
			2251 => "0000000010000000001001011100001000",
			2252 => "0000001110000000001000111000000100",
			2253 => "00000001110011100010010101000101",
			2254 => "11111111000100110010010101000101",
			2255 => "0000001010000000000001010000000100",
			2256 => "00000010101011110010010101000101",
			2257 => "00000000011011110010010101000101",
			2258 => "0000000110000000001101011000001000",
			2259 => "0000001100000000000000101000000100",
			2260 => "11111111000100110010010101000101",
			2261 => "11111111110000100010010101000101",
			2262 => "0000000110000000001101011000000100",
			2263 => "00000010010110000010010101000101",
			2264 => "11111111011100110010010101000101",
			2265 => "0000001100000000000100000000100000",
			2266 => "0000001010000000001010110000010000",
			2267 => "0000000010000000001100010100001100",
			2268 => "0000000110000000001100011000001000",
			2269 => "0000000001000000001100110100000100",
			2270 => "00000010000001010010010101000101",
			2271 => "00000000100110110010010101000101",
			2272 => "00000011111001110010010101000101",
			2273 => "00000000001100100010010101000101",
			2274 => "0000001010000000001100011100001000",
			2275 => "0000001110000000001100101100000100",
			2276 => "11111110011100010010010101000101",
			2277 => "00000000000001000010010101000101",
			2278 => "0000000111000000000100000000000100",
			2279 => "00000000000111100010010101000101",
			2280 => "00000010001011010010010101000101",
			2281 => "0000000110000000001100011000011100",
			2282 => "0000000110000000000100110100001100",
			2283 => "0000000101000000000000001100000100",
			2284 => "11111110101010110010010101000101",
			2285 => "0000000100000000000000010000000100",
			2286 => "11111111000101100010010101000101",
			2287 => "00000001000001000010010101000101",
			2288 => "0000000100000000001001001100001000",
			2289 => "0000000101000000001010111100000100",
			2290 => "00000000000000110010010101000101",
			2291 => "11111110100110000010010101000101",
			2292 => "0000000010000000000010000000000100",
			2293 => "11111101110010110010010101000101",
			2294 => "11111011100110100010010101000101",
			2295 => "0000000110000000001100011000000100",
			2296 => "00000010111111100010010101000101",
			2297 => "0000000101000000000000001100000100",
			2298 => "11111110101100000010010101000101",
			2299 => "0000000001000000000010001100000100",
			2300 => "00000010100000100010010101000101",
			2301 => "00000000000111110010010101000101",
			2302 => "0000001100000000000100000001001100",
			2303 => "0000001001000000001101101000101000",
			2304 => "0000001011000000001001110000100000",
			2305 => "0000000110000000001010011000010000",
			2306 => "0000001110000000001101111000001000",
			2307 => "0000001100000000000100010100000100",
			2308 => "11111111111010000010010101000101",
			2309 => "00000001010101110010010101000101",
			2310 => "0000001100000000000100010100000100",
			2311 => "00000000010001000010010101000101",
			2312 => "11111110001100110010010101000101",
			2313 => "0000000111000000001100001000001000",
			2314 => "0000000011000000000000001100000100",
			2315 => "00000000011010010010010101000101",
			2316 => "11111110010101100010010101000101",
			2317 => "0000000111000000000100000000000100",
			2318 => "00000000110001100010010101000101",
			2319 => "11111111001001010010010101000101",
			2320 => "0000001110000000001110001100000100",
			2321 => "11111111010111000010010101000101",
			2322 => "11111101110100100010010101000101",
			2323 => "0000000011000000000010001000100000",
			2324 => "0000001010000000001010110000010000",
			2325 => "0000000011000000001000000000001000",
			2326 => "0000001001000000001011101000000100",
			2327 => "00000001100000000010010101000101",
			2328 => "00000011001011100010010101000101",
			2329 => "0000000101000000001101010100000100",
			2330 => "11111111101100100010010101000101",
			2331 => "00000001100000100010010101000101",
			2332 => "0000000111000000000100000000001000",
			2333 => "0000001010000000001100011100000100",
			2334 => "11111110101111010010010101000101",
			2335 => "00000000111001100010010101000101",
			2336 => "0000000100000000000100001100000100",
			2337 => "00000000101000110010010101000101",
			2338 => "00000001101100100010010101000101",
			2339 => "11111101111110000010010101000101",
			2340 => "0000000111000000001001110000100100",
			2341 => "0000001110000000001101111000010000",
			2342 => "0000001010000000001010110000000100",
			2343 => "11111110101000000010010101000101",
			2344 => "0000000000000000000100010100000100",
			2345 => "00000010000101100010010101000101",
			2346 => "0000000000000000001011000100000100",
			2347 => "11111111100101000010010101000101",
			2348 => "00000001100001010010010101000101",
			2349 => "0000001010000000000110011000000100",
			2350 => "00000010001101010010010101000101",
			2351 => "0000000100000000001010110100001000",
			2352 => "0000000000000000000000111000000100",
			2353 => "11111110111101110010010101000101",
			2354 => "11111101110100110010010101000101",
			2355 => "0000000100000000000101010100000100",
			2356 => "00000001011001110010010101000101",
			2357 => "11111111010001000010010101000101",
			2358 => "0000000100000000001110100100011000",
			2359 => "0000001001000000001110010100001100",
			2360 => "0000001100000000001000111100000100",
			2361 => "11111110000111010010010101000101",
			2362 => "0000000110000000001001100100000100",
			2363 => "00000000000000000010010101000101",
			2364 => "00000001110001100010010101000101",
			2365 => "0000000101000000001111011100000100",
			2366 => "11111110000001110010010101000101",
			2367 => "0000000101000000000110110100000100",
			2368 => "00000000000010000010010101000101",
			2369 => "11111110100101100010010101000101",
			2370 => "0000000000000000000010111100010000",
			2371 => "0000001001000000001010100000001000",
			2372 => "0000000000000000001000101100000100",
			2373 => "00000101011101100010010101000101",
			2374 => "00000001100010000010010101000101",
			2375 => "0000000111000000000100010000000100",
			2376 => "11111110101110110010010101000101",
			2377 => "00000000011110000010010101000101",
			2378 => "0000001011000000000101101100001000",
			2379 => "0000000000000000001010000000000100",
			2380 => "00000001110111010010010101000101",
			2381 => "00000000000000000010010101000101",
			2382 => "0000001010000000001010110000000100",
			2383 => "11111110111110000010010101000101",
			2384 => "00000000001101100010010101000101",
			2385 => "0000001110000000001100001010111000",
			2386 => "0000001111000000000010001001110000",
			2387 => "0000000100000000000100001100110000",
			2388 => "0000000001000000001110100000011000",
			2389 => "0000001010000000001010110000010000",
			2390 => "0000000110000000001101111100001000",
			2391 => "0000000010000000000101110000000100",
			2392 => "00000000011010010010100000110001",
			2393 => "11111111001011000010100000110001",
			2394 => "0000000000000000000000110000000100",
			2395 => "00000000000000000010100000110001",
			2396 => "00000001100101000010100000110001",
			2397 => "0000001110000000001101010000000100",
			2398 => "11111101101000100010100000110001",
			2399 => "00000000000000000010100000110001",
			2400 => "0000000111000000001011000100001100",
			2401 => "0000000000000000000100010100001000",
			2402 => "0000001101000000001101100000000100",
			2403 => "11111101110111110010100000110001",
			2404 => "11111111110001010010100000110001",
			2405 => "00000001110001010010100000110001",
			2406 => "0000000100000000000100001100001000",
			2407 => "0000001111000000000110110100000100",
			2408 => "00000000001000110010100000110001",
			2409 => "00000000110010010010100000110001",
			2410 => "11111110110010010010100000110001",
			2411 => "0000001000000000000001110100100000",
			2412 => "0000000110000000000001111000010000",
			2413 => "0000000011000000000100010100001000",
			2414 => "0000000011000000000000111000000100",
			2415 => "00000000011010110010100000110001",
			2416 => "11111101010100110010100000110001",
			2417 => "0000000001000000000110000000000100",
			2418 => "00000000000000000010100000110001",
			2419 => "00000001110111100010100000110001",
			2420 => "0000001110000000000000111000001000",
			2421 => "0000001101000000001100110000000100",
			2422 => "11111110100110010010100000110001",
			2423 => "00000001101011010010100000110001",
			2424 => "0000000000000000000111111000000100",
			2425 => "11111111010010010010100000110001",
			2426 => "11111101011001000010100000110001",
			2427 => "0000001101000000001100101100010000",
			2428 => "0000000100000000000010100100001000",
			2429 => "0000000001000000000110000000000100",
			2430 => "11111111010001110010100000110001",
			2431 => "00000000110011000010100000110001",
			2432 => "0000001111000000000110110100000100",
			2433 => "11111111111010110010100000110001",
			2434 => "11111110000000010010100000110001",
			2435 => "0000001010000000001100011100001000",
			2436 => "0000001011000000000100000000000100",
			2437 => "11111101001010110010100000110001",
			2438 => "11111111010110100010100000110001",
			2439 => "0000000100000000000001101100000100",
			2440 => "00000001001001100010100000110001",
			2441 => "11111110001100110010100000110001",
			2442 => "0000001101000000001100101100100100",
			2443 => "0000000011000000000101101100011000",
			2444 => "0000000001000000001100110100010000",
			2445 => "0000001110000000000000101000001000",
			2446 => "0000000010000000001100010100000100",
			2447 => "00000000100011110010100000110001",
			2448 => "11111111011001000010100000110001",
			2449 => "0000000000000000000100010100000100",
			2450 => "00000001101110100010100000110001",
			2451 => "00000000000000010010100000110001",
			2452 => "0000001011000000001100001000000100",
			2453 => "00000000101101100010100000110001",
			2454 => "11111110010010000010100000110001",
			2455 => "0000001111000000000001001000001000",
			2456 => "0000001110000000000000101000000100",
			2457 => "11111100001101100010100000110001",
			2458 => "11111110110001000010100000110001",
			2459 => "00000000000000000010100000110001",
			2460 => "0000000101000000001101111000011000",
			2461 => "0000000101000000000110000100001100",
			2462 => "0000001011000000000100000000001000",
			2463 => "0000000111000000001011000100000100",
			2464 => "11111111101010010010100000110001",
			2465 => "00000001110101110010100000110001",
			2466 => "11111110000101100010100000110001",
			2467 => "0000001000000000001011010100000100",
			2468 => "00000000000000000010100000110001",
			2469 => "0000001000000000001010101100000100",
			2470 => "00000001101011000010100000110001",
			2471 => "00000000011100110010100000110001",
			2472 => "0000000001000000001100110100000100",
			2473 => "11111100110110000010100000110001",
			2474 => "0000000100000000001011100000000100",
			2475 => "00000001101000110010100000110001",
			2476 => "11111111010000000010100000110001",
			2477 => "0000001101000000000000001101011000",
			2478 => "0000000101000000001101111000111000",
			2479 => "0000000001000000001100110100100000",
			2480 => "0000001111000000001011110100010000",
			2481 => "0000001011000000000100000000001000",
			2482 => "0000000010000000000100101000000100",
			2483 => "11111111010011010010100000110001",
			2484 => "11111110000100010010100000110001",
			2485 => "0000001101000000001101111000000100",
			2486 => "00000001011110000010100000110001",
			2487 => "11111111001010100010100000110001",
			2488 => "0000000001000000001100110100001000",
			2489 => "0000000011000000000100001000000100",
			2490 => "00000000010111110010100000110001",
			2491 => "11111110110011010010100000110001",
			2492 => "0000000101000000001110001100000100",
			2493 => "11111111110101010010100000110001",
			2494 => "11111101011110110010100000110001",
			2495 => "0000001110000000001000111000001100",
			2496 => "0000000011000000001110001100000100",
			2497 => "00000010110010110010100000110001",
			2498 => "0000000011000000001101111000000100",
			2499 => "00000000110000010010100000110001",
			2500 => "00000010000101100010100000110001",
			2501 => "0000000100000000000100001100001000",
			2502 => "0000000110000000001010011000000100",
			2503 => "00000000000000000010100000110001",
			2504 => "11111101110011110010100000110001",
			2505 => "00000001111101110010100000110001",
			2506 => "0000000011000000000001111100011000",
			2507 => "0000000001000000001100110100001100",
			2508 => "0000000111000000001100001000000100",
			2509 => "00000000110111110010100000110001",
			2510 => "0000001101000000000000001100000100",
			2511 => "11111101100101100010100000110001",
			2512 => "00000000000000000010100000110001",
			2513 => "0000000100000000000000010100001000",
			2514 => "0000000011000000001101111000000100",
			2515 => "11111111100111110010100000110001",
			2516 => "11111101111111100010100000110001",
			2517 => "11111100101001110010100000110001",
			2518 => "0000001111000000000010110100000100",
			2519 => "00000001000000110010100000110001",
			2520 => "11111111011111010010100000110001",
			2521 => "0000001011000000001000111100101000",
			2522 => "0000000110000000000001111000001000",
			2523 => "0000000001000000001100110100000100",
			2524 => "11111101111101110010100000110001",
			2525 => "00000000000000000010100000110001",
			2526 => "0000001101000000000001111100010000",
			2527 => "0000001011000000001000111100001000",
			2528 => "0000000011000000001101111000000100",
			2529 => "00000001110100110010100000110001",
			2530 => "00000000001001110010100000110001",
			2531 => "0000000011000000001101111000000100",
			2532 => "11111111100000100010100000110001",
			2533 => "00000001100111100010100000110001",
			2534 => "0000001010000000001010110000001000",
			2535 => "0000001000000000000110001000000100",
			2536 => "11111111010110110010100000110001",
			2537 => "00000010001011110010100000110001",
			2538 => "0000000100000000000000010100000100",
			2539 => "11111101110010010010100000110001",
			2540 => "00000000001001110010100000110001",
			2541 => "0000001011000000001000111000100000",
			2542 => "0000001010000000001010110000010000",
			2543 => "0000000010000000001100010100001000",
			2544 => "0000000001000000000010001100000100",
			2545 => "11111111110010100010100000110001",
			2546 => "11111110011001110010100000110001",
			2547 => "0000000011000000000100011000000100",
			2548 => "00000000110110010010100000110001",
			2549 => "00000010101001100010100000110001",
			2550 => "0000000100000000001111100000001000",
			2551 => "0000000101000000000000001100000100",
			2552 => "11111100111111110010100000110001",
			2553 => "11111110101100000010100000110001",
			2554 => "0000000011000000000001111100000100",
			2555 => "11111110111100100010100000110001",
			2556 => "00000000101111110010100000110001",
			2557 => "0000000101000000001100101000010000",
			2558 => "0000000111000000001000111000001000",
			2559 => "0000001000000000000111000100000100",
			2560 => "00000000100100000010100000110001",
			2561 => "11111111010100110010100000110001",
			2562 => "0000001101000000000001111100000100",
			2563 => "00000010111100110010100000110001",
			2564 => "00000001000000000010100000110001",
			2565 => "0000001101000000000001111100001000",
			2566 => "0000000010000000000010000100000100",
			2567 => "11111111000111000010100000110001",
			2568 => "00000010000001100010100000110001",
			2569 => "0000000011000000000100001000000100",
			2570 => "00000001010000110010100000110001",
			2571 => "11111111111101100010100000110001",
			2572 => "0000001111000000000000110111010100",
			2573 => "0000001110000000001010000001110100",
			2574 => "0000001011000000000100010100110100",
			2575 => "0000000001000000001110100000011100",
			2576 => "0000001001000000001001111000010000",
			2577 => "0000001100000000000111111000001000",
			2578 => "0000000111000000000111111000000100",
			2579 => "11111111111000000010101100000111",
			2580 => "00000000110000100010101100000111",
			2581 => "0000001110000000000011111100000100",
			2582 => "11111111110000110010101100000111",
			2583 => "11111110101101110010101100000111",
			2584 => "0000001011000000000100010100001000",
			2585 => "0000001100000000000111111000000100",
			2586 => "00000000010111100010101100000111",
			2587 => "00000001110110100010101100000111",
			2588 => "11111111000010010010101100000111",
			2589 => "0000001100000000000111111000001100",
			2590 => "0000001001000000001001111000000100",
			2591 => "11111110110000100010101100000111",
			2592 => "0000000011000000001100001000000100",
			2593 => "00000001111000010010101100000111",
			2594 => "11111111111101000010101100000111",
			2595 => "0000000111000000001011000100001000",
			2596 => "0000001101000000000101101100000100",
			2597 => "11111101010001000010101100000111",
			2598 => "11111111000111100010101100000111",
			2599 => "00000000101010110010101100000111",
			2600 => "0000000110000000000100110100100000",
			2601 => "0000001110000000000000111000010000",
			2602 => "0000001001000000000010001100001000",
			2603 => "0000000001000000000110000000000100",
			2604 => "00000000110000100010101100000111",
			2605 => "11111100101011010010101100000111",
			2606 => "0000001000000000001011010100000100",
			2607 => "00000000001110110010101100000111",
			2608 => "00000001011000000010101100000111",
			2609 => "0000001001000000001001111000001000",
			2610 => "0000000101000000001101100000000100",
			2611 => "11111111100010100010101100000111",
			2612 => "11111101000101010010101100000111",
			2613 => "0000001111000000000111010000000100",
			2614 => "11111111111010110010101100000111",
			2615 => "00000000110011000010101100000111",
			2616 => "0000001111000000000100000100010000",
			2617 => "0000001111000000001000011000001000",
			2618 => "0000000100000000000000101100000100",
			2619 => "00000001101011110010101100000111",
			2620 => "11111110110000100010101100000111",
			2621 => "0000000111000000001100001000000100",
			2622 => "11111101110011010010101100000111",
			2623 => "00000001011010100010101100000111",
			2624 => "0000001101000000001110001100001000",
			2625 => "0000000101000000001101100000000100",
			2626 => "11111111001010000010101100000111",
			2627 => "00000001100100100010101100000111",
			2628 => "0000001001000000000110101000000100",
			2629 => "11111101101010100010101100000111",
			2630 => "00000001001010100010101100000111",
			2631 => "0000001101000000001100101100100100",
			2632 => "0000001100000000000000101000100000",
			2633 => "0000000011000000000101101100010000",
			2634 => "0000001111000000001011011100001000",
			2635 => "0000001011000000000100010100000100",
			2636 => "00000001000100010010101100000111",
			2637 => "11111111000110110010101100000111",
			2638 => "0000000011000000001001110000000100",
			2639 => "00000000110101100010101100000111",
			2640 => "11111111111000100010101100000111",
			2641 => "0000001111000000000111110000001000",
			2642 => "0000000100000000000010110000000100",
			2643 => "11111111110101100010101100000111",
			2644 => "11111101110111110010101100000111",
			2645 => "0000001000000000000110001000000100",
			2646 => "00000010001101110010101100000111",
			2647 => "11111111010100100010101100000111",
			2648 => "11111101011100110010101100000111",
			2649 => "0000001110000000001101100000100000",
			2650 => "0000001001000000000111100100010000",
			2651 => "0000000001000000001100110100001000",
			2652 => "0000001001000000000110101000000100",
			2653 => "11111111111010000010101100000111",
			2654 => "00000000111100010010101100000111",
			2655 => "0000001100000000000100000000000100",
			2656 => "11111111110101010010101100000111",
			2657 => "11111101100010010010101100000111",
			2658 => "0000000100000000000011001100001000",
			2659 => "0000000011000000001110001100000100",
			2660 => "00000001010001000010101100000111",
			2661 => "11111111010010100010101100000111",
			2662 => "0000000110000000001010011000000100",
			2663 => "00000001100010000010101100000111",
			2664 => "00000000000111100010101100000111",
			2665 => "0000001001000000001011101000010000",
			2666 => "0000001100000000000100010100001000",
			2667 => "0000001100000000000100010100000100",
			2668 => "11111111100011110010101100000111",
			2669 => "00000001011000010010101100000111",
			2670 => "0000001011000000000100000000000100",
			2671 => "11111110100000010010101100000111",
			2672 => "11111111011001110010101100000111",
			2673 => "0000001000000000000111000100001000",
			2674 => "0000000001000000001001111000000100",
			2675 => "00000000010101000010101100000111",
			2676 => "11111111010010010010101100000111",
			2677 => "00000010000110100010101100000111",
			2678 => "0000000111000000000100000001100000",
			2679 => "0000001010000000001100011100110100",
			2680 => "0000000100000000001010110100011100",
			2681 => "0000001100000000000100000000010000",
			2682 => "0000000110000000001101111100001000",
			2683 => "0000000001000000001110100000000100",
			2684 => "00000000000000000010101100000111",
			2685 => "00000010001000000010101100000111",
			2686 => "0000000100000000001011110000000100",
			2687 => "11111110001111010010101100000111",
			2688 => "00000000000000000010101100000111",
			2689 => "0000001101000000001010111000001000",
			2690 => "0000001000000000000110001000000100",
			2691 => "00000010110011000010101100000111",
			2692 => "00000000011010000010101100000111",
			2693 => "11111111000001010010101100000111",
			2694 => "0000001101000000000101101100001100",
			2695 => "0000000111000000000111111000001000",
			2696 => "0000001111000000001110101100000100",
			2697 => "00000001001101010010101100000111",
			2698 => "00000000000000000010101100000111",
			2699 => "11111101100101110010101100000111",
			2700 => "0000001100000000000100000000001000",
			2701 => "0000001101000000000000001100000100",
			2702 => "00000000100110110010101100000111",
			2703 => "00000001011010010010101100000111",
			2704 => "11111111011111010010101100000111",
			2705 => "0000001011000000001001110000100000",
			2706 => "0000000100000000000011010100010000",
			2707 => "0000000101000000000000001100001000",
			2708 => "0000001001000000000111100100000100",
			2709 => "11111110011110100010101100000111",
			2710 => "00000000001111010010101100000111",
			2711 => "0000000110000000001010011000000100",
			2712 => "11111101000000110010101100000111",
			2713 => "11111110011100010010101100000111",
			2714 => "0000000111000000001100001000001000",
			2715 => "0000001110000000001000111000000100",
			2716 => "00000001101011000010101100000111",
			2717 => "11111111010111100010101100000111",
			2718 => "0000001100000000000100010100000100",
			2719 => "00000000000000000010101100000111",
			2720 => "00000001101110000010101100000111",
			2721 => "0000001100000000000000101000000100",
			2722 => "11111110011110100010101100000111",
			2723 => "0000001110000000001100101100000100",
			2724 => "00000000110000110010101100000111",
			2725 => "00000010011010000010101100000111",
			2726 => "0000000111000000001000111000011100",
			2727 => "0000001111000000000000110100000100",
			2728 => "00000001010111100010101100000111",
			2729 => "0000001100000000000100000000001100",
			2730 => "0000000111000000001000111100001000",
			2731 => "0000001001000000001011101000000100",
			2732 => "11111110001000000010101100000111",
			2733 => "11111111110010110010101100000111",
			2734 => "11111101110110010010101100000111",
			2735 => "0000001100000000001000111000001000",
			2736 => "0000000101000000000100001000000100",
			2737 => "00000001110010010010101100000111",
			2738 => "11111111110110000010101100000111",
			2739 => "11111101011101000010101100000111",
			2740 => "0000000011000000000100001000000100",
			2741 => "11111101101010010010101100000111",
			2742 => "0000001001000000000111100100001000",
			2743 => "0000001111000000001110101100000100",
			2744 => "00000001010010110010101100000111",
			2745 => "00000011000000000010101100000111",
			2746 => "0000001100000000000000101000001000",
			2747 => "0000000110000000001010011000000100",
			2748 => "11111111110111110010101100000111",
			2749 => "00000001001000110010101100000111",
			2750 => "0000001100000000000000101000000100",
			2751 => "11111110110010010010101100000111",
			2752 => "00000000000001010010101100000111",
			2753 => "0000000100000000000001001101001000",
			2754 => "0000000100000000000110111100001000",
			2755 => "0000000111000000000100010100000100",
			2756 => "00000000000000000010101111010001",
			2757 => "11111110011100100010101111010001",
			2758 => "0000000011000000000011111100001100",
			2759 => "0000001011000000001010000000000100",
			2760 => "11111111110011110010101111010001",
			2761 => "0000001001000000001100110100000100",
			2762 => "00000001111010010010101111010001",
			2763 => "00000000111011010010101111010001",
			2764 => "0000001001000000001100110100011000",
			2765 => "0000000011000000000000111000001000",
			2766 => "0000001110000000000111000100000100",
			2767 => "11111110011100100010101111010001",
			2768 => "00000001011011100010101111010001",
			2769 => "0000001100000000000000111000001000",
			2770 => "0000001100000000000011111100000100",
			2771 => "11111111101011100010101111010001",
			2772 => "00000001100001110010101111010001",
			2773 => "0000000111000000000111111000000100",
			2774 => "11111101101100010010101111010001",
			2775 => "11111111100011010010101111010001",
			2776 => "0000001110000000001000110000001100",
			2777 => "0000000010000000001111010000001000",
			2778 => "0000000011000000000011010000000100",
			2779 => "11111110100011000010101111010001",
			2780 => "00000001011100010010101111010001",
			2781 => "11111110100011110010101111010001",
			2782 => "0000001111000000000010001000001000",
			2783 => "0000001110000000000111111000000100",
			2784 => "00000000001000000010101111010001",
			2785 => "11111111101010100010101111010001",
			2786 => "0000000011000000001100101100000100",
			2787 => "00000000011101110010101111010001",
			2788 => "00000000000100110010101111010001",
			2789 => "0000000111000000001100001000011100",
			2790 => "0000001100000000000111111000010100",
			2791 => "0000001101000000000100000000000100",
			2792 => "11111110011100110010101111010001",
			2793 => "0000001101000000000011011100001100",
			2794 => "0000000010000000000111111100001000",
			2795 => "0000000010000000001101000100000100",
			2796 => "11111111100011110010101111010001",
			2797 => "00000000110110010010101111010001",
			2798 => "11111111100010100010101111010001",
			2799 => "11111110011000110010101111010001",
			2800 => "0000000010000000001111010000000100",
			2801 => "11111111101001110010101111010001",
			2802 => "00000001001010000010101111010001",
			2803 => "11111110011010110010101111010001",
			2804 => "0000001001000000001001111000111100",
			2805 => "0000000111000000001100001000110100",
			2806 => "0000000111000000001100001000110000",
			2807 => "0000000011000000001100001000011100",
			2808 => "0000000010000000000111111100010000",
			2809 => "0000000100000000000011010100001000",
			2810 => "0000000010000000001111010000000100",
			2811 => "00000000000000000010110011101101",
			2812 => "00000001000110010010110011101101",
			2813 => "0000001110000000000011111100000100",
			2814 => "11111111110010010010110011101101",
			2815 => "11111110011100010010110011101101",
			2816 => "0000001001000000001100110100000100",
			2817 => "11111110101100000010110011101101",
			2818 => "0000000101000000000011011100000100",
			2819 => "00000001111011110010110011101101",
			2820 => "00000000110011000010110011101101",
			2821 => "0000000101000000000110000100010000",
			2822 => "0000000010000000001110101000001000",
			2823 => "0000001000000000001100000100000100",
			2824 => "00000000100011000010110011101101",
			2825 => "11111101001111100010110011101101",
			2826 => "0000001100000000000100010100000100",
			2827 => "11111111011010100010110011101101",
			2828 => "00000000001111010010110011101101",
			2829 => "00000001100010000010110011101101",
			2830 => "11111101101110110010110011101101",
			2831 => "0000000100000000000010010000000100",
			2832 => "00000001110100010010110011101101",
			2833 => "11111110111000010010110011101101",
			2834 => "0000001110000000000011010000010000",
			2835 => "0000000010000000001010010100000100",
			2836 => "11111111010111010010110011101101",
			2837 => "0000001001000000001001111000001000",
			2838 => "0000000100000000001001001100000100",
			2839 => "00000001101011000010110011101101",
			2840 => "00000000000000000010110011101101",
			2841 => "00000001110110010010110011101101",
			2842 => "0000001100000000001010000000010100",
			2843 => "0000001110000000000100000000001100",
			2844 => "0000001010000000000110011000000100",
			2845 => "00000010001010100010110011101101",
			2846 => "0000000100000000000100001100000100",
			2847 => "00000000000000000010110011101101",
			2848 => "00000001110010110010110011101101",
			2849 => "0000000010000000001010001000000100",
			2850 => "11111110100011000010110011101101",
			2851 => "00000001011101100010110011101101",
			2852 => "0000001100000000001110111100010000",
			2853 => "0000000010000000001100010100001100",
			2854 => "0000001101000000000101101100000100",
			2855 => "11111110010101110010110011101101",
			2856 => "0000001000000000001111001000000100",
			2857 => "11111111101001000010110011101101",
			2858 => "00000001010010010010110011101101",
			2859 => "11111110000001100010110011101101",
			2860 => "0000000100000000000100001100010000",
			2861 => "0000000000000000000100010100001000",
			2862 => "0000001000000000000001110100000100",
			2863 => "11111111111111010010110011101101",
			2864 => "11111111010101000010110011101101",
			2865 => "0000001110000000001100110000000100",
			2866 => "00000001111011010010110011101101",
			2867 => "00000000110100110010110011101101",
			2868 => "0000001000000000000111000100001000",
			2869 => "0000000111000000001100001000000100",
			2870 => "00000000000001010010110011101101",
			2871 => "11111101111110000010110011101101",
			2872 => "0000001000000000000010101000000100",
			2873 => "00000000101111010010110011101101",
			2874 => "00000000000001000010110011101101",
			2875 => "0000001100000000001110001101011100",
			2876 => "0000000100000000001011100101010000",
			2877 => "0000000100000000000000010000010000",
			2878 => "0000001110000000001000111000000100",
			2879 => "11111111011111010010111000101001",
			2880 => "0000001011000000001110001100000100",
			2881 => "11111110000100010010111000101001",
			2882 => "0000001011000000001101111000000100",
			2883 => "00000000000000010010111000101001",
			2884 => "11111110011010100010111000101001",
			2885 => "0000001100000000000000101000100000",
			2886 => "0000001110000000000000001100010000",
			2887 => "0000001001000000001101101000001000",
			2888 => "0000001110000000001100001000000100",
			2889 => "00000000011001100010111000101001",
			2890 => "00000000000100000010111000101001",
			2891 => "0000001111000000001001010100000100",
			2892 => "00000000010111010010111000101001",
			2893 => "00000010000010100010111000101001",
			2894 => "0000001100000000000100010100001000",
			2895 => "0000000110000000001101011000000100",
			2896 => "00000000101100110010111000101001",
			2897 => "11111110101011000010111000101001",
			2898 => "0000001011000000000101101100000100",
			2899 => "11111110111110100010111000101001",
			2900 => "00000001011010010010111000101001",
			2901 => "0000001100000000000000101000010000",
			2902 => "0000001010000000000110011000001000",
			2903 => "0000000010000000000111111100000100",
			2904 => "00000001011001100010111000101001",
			2905 => "00000011001110010010111000101001",
			2906 => "0000001000000000001011010100000100",
			2907 => "11111110000100100010111000101001",
			2908 => "00000001000000110010111000101001",
			2909 => "0000001100000000000000101000001000",
			2910 => "0000000010000000000101110000000100",
			2911 => "00000000100010010010111000101001",
			2912 => "11111101101010010010111000101001",
			2913 => "0000001111000000001101000100000100",
			2914 => "00000000101101100010111000101001",
			2915 => "00000000001000110010111000101001",
			2916 => "0000001001000000000110000000000100",
			2917 => "11111110011000110010111000101001",
			2918 => "0000001111000000001001001000000100",
			2919 => "00000001000111010010111000101001",
			2920 => "11111110010000100010111000101001",
			2921 => "0000001000000000001001101000001100",
			2922 => "0000001110000000001010001100001000",
			2923 => "0000000101000000000100000100000100",
			2924 => "11111111111001100010111000101001",
			2925 => "00000010000101100010111000101001",
			2926 => "11111110011010000010111000101001",
			2927 => "0000000100000000000110110000101100",
			2928 => "0000001000000000000110001000010000",
			2929 => "0000000010000000000101000000001100",
			2930 => "0000000101000000001111010000001000",
			2931 => "0000001111000000000110111000000100",
			2932 => "00000001011000110010111000101001",
			2933 => "11111110100000100010111000101001",
			2934 => "00000010010101000010111000101001",
			2935 => "11111110011000110010111000101001",
			2936 => "0000000100000000000011101100010000",
			2937 => "0000000100000000001001001100001000",
			2938 => "0000001010000000001100011100000100",
			2939 => "00000000011110000010111000101001",
			2940 => "11111110101101100010111000101001",
			2941 => "0000001110000000001000001000000100",
			2942 => "00000010011111100010111000101001",
			2943 => "00000000000000000010111000101001",
			2944 => "0000001000000000000001110100000100",
			2945 => "11111110000110100010111000101001",
			2946 => "0000000110000000001001111100000100",
			2947 => "11111111000001010010111000101001",
			2948 => "00000001011110010010111000101001",
			2949 => "0000001100000000000000001100001000",
			2950 => "0000000100000000000011000100000100",
			2951 => "00000001011000010010111000101001",
			2952 => "11111110100001000010111000101001",
			2953 => "11111110011000110010111000101001",
			2954 => "0000000100000000000001001101111000",
			2955 => "0000001000000000001101010001101000",
			2956 => "0000000100000000000011011001000000",
			2957 => "0000001110000000000011010000100000",
			2958 => "0000001111000000000001101000010000",
			2959 => "0000001110000000001000110000001000",
			2960 => "0000000101000000001000111000000100",
			2961 => "11111111110101000010111101000101",
			2962 => "00000001010100110010111101000101",
			2963 => "0000000111000000000000101000000100",
			2964 => "11111110111011010010111101000101",
			2965 => "00000001110100010010111101000101",
			2966 => "0000001001000000000010001100001000",
			2967 => "0000001110000000001111000100000100",
			2968 => "00000001000111000010111101000101",
			2969 => "11111111000000110010111101000101",
			2970 => "0000000111000000000000101000000100",
			2971 => "00000001001011100010111101000101",
			2972 => "11111111011100100010111101000101",
			2973 => "0000000111000000000111111000010000",
			2974 => "0000000111000000001110111100001000",
			2975 => "0000001100000000001010000000000100",
			2976 => "11111101110101100010111101000101",
			2977 => "00000001000101000010111101000101",
			2978 => "0000001100000000000000110000000100",
			2979 => "11111111110101010010111101000101",
			2980 => "11111101001010110010111101000101",
			2981 => "0000001111000000000101100100001000",
			2982 => "0000001011000000000100010100000100",
			2983 => "11111110100100000010111101000101",
			2984 => "11111111110111010010111101000101",
			2985 => "0000000110000000001010011000000100",
			2986 => "00000000001100100010111101000101",
			2987 => "11111111111010010010111101000101",
			2988 => "0000001111000000001001001000001000",
			2989 => "0000001100000000000111111000000100",
			2990 => "11111111011100110010111101000101",
			2991 => "00000001111011010010111101000101",
			2992 => "0000001000000000000111000000010000",
			2993 => "0000001010000000000110011100001000",
			2994 => "0000001000000000000010101000000100",
			2995 => "11111101110010110010111101000101",
			2996 => "00000000110101000010111101000101",
			2997 => "0000000010000000001111010100000100",
			2998 => "11111011001100110010111101000101",
			2999 => "11111110101010110010111101000101",
			3000 => "0000001100000000000100010100001000",
			3001 => "0000000111000000001011000100000100",
			3002 => "11111111100011110010111101000101",
			3003 => "11111101001110010010111101000101",
			3004 => "0000001010000000000001010100000100",
			3005 => "00000001101101000010111101000101",
			3006 => "11111111101001010010111101000101",
			3007 => "0000000110000000001010011000000100",
			3008 => "00000000000101100010111101000101",
			3009 => "0000001010000000001001101000001000",
			3010 => "0000001010000000001100000100000100",
			3011 => "00000001100101100010111101000101",
			3012 => "00000000000000000010111101000101",
			3013 => "00000010010010110010111101000101",
			3014 => "0000000111000000001100001000010100",
			3015 => "0000001100000000000111111000001100",
			3016 => "0000000101000000001001110000000100",
			3017 => "11111110101001110010111101000101",
			3018 => "0000000101000000000011011100000100",
			3019 => "00000000100000010010111101000101",
			3020 => "11111110100000000010111101000101",
			3021 => "0000000100000000000100100000000100",
			3022 => "00000000111111100010111101000101",
			3023 => "11111111111010100010111101000101",
			3024 => "11111110011011110010111101000101",
			3025 => "0000001110000000000011111101010100",
			3026 => "0000000100000000001001000000101000",
			3027 => "0000000010000000001111010000011100",
			3028 => "0000000000000000000000101000010100",
			3029 => "0000000100000000000010100100001100",
			3030 => "0000001000000000000010101000001000",
			3031 => "0000000000000000000100010100000100",
			3032 => "00000000001101100011000011110001",
			3033 => "00000001100101000011000011110001",
			3034 => "11111101111111100011000011110001",
			3035 => "0000001101000000001101100000000100",
			3036 => "11111111110110100011000011110001",
			3037 => "11111100010001010011000011110001",
			3038 => "0000001010000000001100011100000100",
			3039 => "00000000011100100011000011110001",
			3040 => "00000001100111110011000011110001",
			3041 => "0000001001000000001100110100000100",
			3042 => "11111110001100010011000011110001",
			3043 => "0000000000000000000100010100000100",
			3044 => "00000000111010100011000011110001",
			3045 => "00000001111100000011000011110001",
			3046 => "0000001001000000000010001100100100",
			3047 => "0000001101000000001101100000011000",
			3048 => "0000000101000000000011011100010000",
			3049 => "0000000110000000000100110100001000",
			3050 => "0000000111000000000100010100000100",
			3051 => "11111101101011100011000011110001",
			3052 => "00000000100101110011000011110001",
			3053 => "0000000101000000001001110000000100",
			3054 => "11111111111101100011000011110001",
			3055 => "00000001100110100011000011110001",
			3056 => "0000001001000000000000011000000100",
			3057 => "00000000000000000011000011110001",
			3058 => "11111100101100110011000011110001",
			3059 => "0000000100000000000110110000000100",
			3060 => "00000001101101010011000011110001",
			3061 => "0000000111000000000100010100000100",
			3062 => "00000000000000000011000011110001",
			3063 => "11111110101010010011000011110001",
			3064 => "0000000100000000001100111100000100",
			3065 => "00000001110010110011000011110001",
			3066 => "11111111101011000011000011110001",
			3067 => "0000001001000000001001111000111100",
			3068 => "0000001111000000001010001100011000",
			3069 => "0000000100000000001101001000010000",
			3070 => "0000000100000000000110001100001000",
			3071 => "0000001111000000000001101000000100",
			3072 => "11111111011100000011000011110001",
			3073 => "11111101010110000011000011110001",
			3074 => "0000001110000000000011010000000100",
			3075 => "00000010000010100011000011110001",
			3076 => "11111111011000110011000011110001",
			3077 => "0000001010000000001010110000000100",
			3078 => "11111011101110110011000011110001",
			3079 => "11111101101010100011000011110001",
			3080 => "0000000011000000000000101000000100",
			3081 => "00000001101001010011000011110001",
			3082 => "0000001010000000001001000100010000",
			3083 => "0000000011000000000100000000001000",
			3084 => "0000001001000000000010001100000100",
			3085 => "11111110001000110011000011110001",
			3086 => "00000001111110010011000011110001",
			3087 => "0000000000000000000011010000000100",
			3088 => "11111111001110100011000011110001",
			3089 => "00000010011111100011000011110001",
			3090 => "0000001111000000000110110100001000",
			3091 => "0000000011000000001000111100000100",
			3092 => "11111111001101000011000011110001",
			3093 => "11111101001111110011000011110001",
			3094 => "0000000010000000000100101000000100",
			3095 => "00000001011111100011000011110001",
			3096 => "11111111101011100011000011110001",
			3097 => "0000000101000000000011011100010100",
			3098 => "0000000110000000001101111100001100",
			3099 => "0000000000000000000011111100000100",
			3100 => "11111110010100010011000011110001",
			3101 => "0000001111000000000110110100000100",
			3102 => "00000001011011010011000011110001",
			3103 => "11111111010111110011000011110001",
			3104 => "0000001011000000000100010100000100",
			3105 => "11111101101001100011000011110001",
			3106 => "11111111001011000011000011110001",
			3107 => "0000000011000000001100110000010100",
			3108 => "0000001101000000001101111000010000",
			3109 => "0000001111000000001111011100001000",
			3110 => "0000000011000000001000111100000100",
			3111 => "00000000011001110011000011110001",
			3112 => "11111110100101010011000011110001",
			3113 => "0000000111000000000111111000000100",
			3114 => "11111110101111010011000011110001",
			3115 => "00000000011010010011000011110001",
			3116 => "00000010000101000011000011110001",
			3117 => "0000001111000000001010010100010000",
			3118 => "0000001001000000000110101000001000",
			3119 => "0000001111000000000111110000000100",
			3120 => "11111110111101000011000011110001",
			3121 => "00000000011001010011000011110001",
			3122 => "0000001111000000000111110000000100",
			3123 => "11111111111101100011000011110001",
			3124 => "11111111001001100011000011110001",
			3125 => "0000000011000000001101111000001000",
			3126 => "0000000000000000000000110000000100",
			3127 => "00000010000001010011000011110001",
			3128 => "00000000011011000011000011110001",
			3129 => "0000001001000000000111100100000100",
			3130 => "11111111001010000011000011110001",
			3131 => "00000000000101000011000011110001",
			3132 => "0000001000000000000111000001101100",
			3133 => "0000001010000000000110011101001100",
			3134 => "0000000011000000000000110000001100",
			3135 => "0000000110000000001110010100000100",
			3136 => "11111110010101010011001001110101",
			3137 => "0000001011000000001110111100000100",
			3138 => "11111111111000110011001001110101",
			3139 => "00000001101111010011001001110101",
			3140 => "0000001001000000001001111000100000",
			3141 => "0000000011000000001000111100010000",
			3142 => "0000000010000000001111010000001000",
			3143 => "0000000100000000000010111000000100",
			3144 => "00000000010010000011001001110101",
			3145 => "11111111011110100011001001110101",
			3146 => "0000001100000000000111111000000100",
			3147 => "00000000000011000011001001110101",
			3148 => "00000001011100110011001001110101",
			3149 => "0000000101000000001101100000001000",
			3150 => "0000000110000000000100110100000100",
			3151 => "11111111001010000011001001110101",
			3152 => "00000001011101000011001001110101",
			3153 => "0000001110000000001110111100000100",
			3154 => "11111111010010110011001001110101",
			3155 => "11111101100111010011001001110101",
			3156 => "0000000001000000001110100000010000",
			3157 => "0000000101000000001100110000001000",
			3158 => "0000000101000000000011011100000100",
			3159 => "11111111110111100011001001110101",
			3160 => "00000000111111110011001001110101",
			3161 => "0000000111000000000100010100000100",
			3162 => "11111110000000000011001001110101",
			3163 => "00000000001000100011001001110101",
			3164 => "0000001001000000000110101000001000",
			3165 => "0000000111000000000100010100000100",
			3166 => "00000000001100110011001001110101",
			3167 => "11111111011010100011001001110101",
			3168 => "0000001110000000000000101000000100",
			3169 => "00000000010101010011001001110101",
			3170 => "00000000000000000011001001110101",
			3171 => "0000001001000000000110101000000100",
			3172 => "11111100110111010011001001110101",
			3173 => "0000001011000000001000111100001000",
			3174 => "0000000100000000001111100000000100",
			3175 => "11111110111101000011001001110101",
			3176 => "00000001101001000011001001110101",
			3177 => "0000001001000000001011101000001000",
			3178 => "0000001110000000001101100000000100",
			3179 => "00000000000000000011001001110101",
			3180 => "11111101001101010011001001110101",
			3181 => "0000001110000000001010111000000100",
			3182 => "00000001011011010011001001110101",
			3183 => "0000000001000000001001111000000100",
			3184 => "11111110000100100011001001110101",
			3185 => "11111111111101110011001001110101",
			3186 => "0000000100000000000011011000010100",
			3187 => "0000000100000000001001000000010000",
			3188 => "0000001011000000001011000100000100",
			3189 => "00000001100101000011001001110101",
			3190 => "0000001011000000001100001000000100",
			3191 => "11111110001011110011001001110101",
			3192 => "0000000110000000001011001100000100",
			3193 => "00000001101001000011001001110101",
			3194 => "11111111000100100011001001110101",
			3195 => "00000001101111110011001001110101",
			3196 => "0000001100000000000111111000011000",
			3197 => "0000001011000000000100010100010000",
			3198 => "0000000111000000000111111000000100",
			3199 => "11111110100010010011001001110101",
			3200 => "0000000100000000000110110000000100",
			3201 => "00000001010100000011001001110101",
			3202 => "0000001010000000000110001000000100",
			3203 => "11111110110101110011001001110101",
			3204 => "00000000000000000011001001110101",
			3205 => "0000000011000000001000101100000100",
			3206 => "00000000110001100011001001110101",
			3207 => "11111100100010110011001001110101",
			3208 => "0000000111000000001011000100010100",
			3209 => "0000000100000000000010010000001000",
			3210 => "0000000101000000001101100000000100",
			3211 => "00000010000110000011001001110101",
			3212 => "00000000111111100011001001110101",
			3213 => "0000000110000000000100110100001000",
			3214 => "0000001010000000001100000100000100",
			3215 => "11111110101100000011001001110101",
			3216 => "00000000000000000011001001110101",
			3217 => "00000000111110000011001001110101",
			3218 => "0000001100000000000100010100001000",
			3219 => "0000000111000000001100001000000100",
			3220 => "11111110000011100011001001110101",
			3221 => "00000000010000000011001001110101",
			3222 => "0000000000000000001100101100001000",
			3223 => "0000001001000000000110101000000100",
			3224 => "00000001101100010011001001110101",
			3225 => "00000000011010110011001001110101",
			3226 => "0000000010000000001110110100000100",
			3227 => "00000000000000000011001001110101",
			3228 => "11111110101101100011001001110101",
			3229 => "0000000111000000001100101001100100",
			3230 => "0000000100000000000110110001000100",
			3231 => "0000000110000000000001000100000100",
			3232 => "11111110010111100011001111011001",
			3233 => "0000001110000000000100010100100000",
			3234 => "0000000101000000000110000100010000",
			3235 => "0000000011000000000111111000001000",
			3236 => "0000001001000000001100110100000100",
			3237 => "00000000101100010011001111011001",
			3238 => "00000001100001000011001111011001",
			3239 => "0000001001000000001100110100000100",
			3240 => "11111110000100000011001111011001",
			3241 => "00000000101001100011001111011001",
			3242 => "0000001011000000000100000000001000",
			3243 => "0000001111000000001000011000000100",
			3244 => "00000000010010000011001111011001",
			3245 => "00000001111101100011001111011001",
			3246 => "0000000111000000001100001000000100",
			3247 => "00000000001011110011001111011001",
			3248 => "00000001101011110011001111011001",
			3249 => "0000000010000000001010001000010000",
			3250 => "0000000110000000000001111000001000",
			3251 => "0000000101000000001110001100000100",
			3252 => "00000000001110000011001111011001",
			3253 => "00000001111011100011001111011001",
			3254 => "0000000010000000001110000100000100",
			3255 => "11111111001111010011001111011001",
			3256 => "00000000001111010011001111011001",
			3257 => "0000000110000000001100011000001000",
			3258 => "0000001101000000000101101100000100",
			3259 => "11111111100110110011001111011001",
			3260 => "00000001010010000011001111011001",
			3261 => "0000000100000000000100001100000100",
			3262 => "00000000010000000011001111011001",
			3263 => "00000000111100110011001111011001",
			3264 => "0000000010000000000010010100011100",
			3265 => "0000000001000000001110100000010100",
			3266 => "0000001110000000001000101100001100",
			3267 => "0000000001000000001100100000000100",
			3268 => "11111110010111010011001111011001",
			3269 => "0000000100000000000011111000000100",
			3270 => "11111110010010000011001111011001",
			3271 => "00000000101000000011001111011001",
			3272 => "0000000001000000000000011000000100",
			3273 => "11111110101001100011001111011001",
			3274 => "11111100110010010011001111011001",
			3275 => "0000001110000000000100000000000100",
			3276 => "00000000111101010011001111011001",
			3277 => "11111110011001110011001111011001",
			3278 => "00000000000000000011001111011001",
			3279 => "0000001000000000001001101000010100",
			3280 => "0000001100000000000110000100001000",
			3281 => "0000001100000000000110000100000100",
			3282 => "11111110110001000011001111011001",
			3283 => "00000010001000000011001111011001",
			3284 => "0000001110000000001010001100001000",
			3285 => "0000000101000000000100000100000100",
			3286 => "11111110110010000011001111011001",
			3287 => "00000010111110010011001111011001",
			3288 => "11111110010110110011001111011001",
			3289 => "0000000100000000000010010000100100",
			3290 => "0000001000000000000111000000100000",
			3291 => "0000001111000000001011110000010000",
			3292 => "0000000100000000000011110100001000",
			3293 => "0000001100000000000100001000000100",
			3294 => "00000000000000000011001111011001",
			3295 => "00000010100011010011001111011001",
			3296 => "0000001001000000001101011000000100",
			3297 => "00000000111100100011001111011001",
			3298 => "11111110011010000011001111011001",
			3299 => "0000001100000000000111010000001000",
			3300 => "0000001000000000000111000100000100",
			3301 => "11111110010111010011001111011001",
			3302 => "00000000000100110011001111011001",
			3303 => "0000001111000000000010111000000100",
			3304 => "00000011101011110011001111011001",
			3305 => "11111111100000010011001111011001",
			3306 => "00000010001100010011001111011001",
			3307 => "0000000100000000000000000000010100",
			3308 => "0000001000000000000000110000001100",
			3309 => "0000000100000000000011111000001000",
			3310 => "0000000100000000001011100100000100",
			3311 => "11111110011101110011001111011001",
			3312 => "00000000001110100011001111011001",
			3313 => "11111110011011100011001111011001",
			3314 => "0000001000000000001010000000000100",
			3315 => "00000001001000010011001111011001",
			3316 => "11111110101110010011001111011001",
			3317 => "11111110010111010011001111011001",
			3318 => "0000000111000000001110001110000000",
			3319 => "0000000001000000000000011000010000",
			3320 => "0000000001000000001100100000000100",
			3321 => "11111110001110110011010101001101",
			3322 => "0000000011000000001000110000000100",
			3323 => "00000010100100000011010101001101",
			3324 => "0000000111000000000111111000000100",
			3325 => "11111110001110010011010101001101",
			3326 => "00000000011111100011010101001101",
			3327 => "0000001110000000001101100000111100",
			3328 => "0000000000000000000100010100100000",
			3329 => "0000000011000000000100000000010000",
			3330 => "0000001001000000001100110100001000",
			3331 => "0000000011000000000000111000000100",
			3332 => "00000011000111000011010101001101",
			3333 => "11111101101001010011010101001101",
			3334 => "0000000100000000000011010100000100",
			3335 => "00000010010010010011010101001101",
			3336 => "00000000011110000011010101001101",
			3337 => "0000001001000000000010001100001000",
			3338 => "0000001100000000000111111000000100",
			3339 => "11111101111100100011010101001101",
			3340 => "11111110110100010011010101001101",
			3341 => "0000000010000000001010001000000100",
			3342 => "00000001010101100011010101001101",
			3343 => "00000010010100010011010101001101",
			3344 => "0000000100000000000110110000010000",
			3345 => "0000000111000000000111111000001000",
			3346 => "0000000010000000001110000100000100",
			3347 => "00000010101100110011010101001101",
			3348 => "00000000111000100011010101001101",
			3349 => "0000001000000000000111000000000100",
			3350 => "00000010011000100011010101001101",
			3351 => "00000010110111010011010101001101",
			3352 => "0000000000000000001101111000000100",
			3353 => "11111110100010110011010101001101",
			3354 => "0000001111000000001110101100000100",
			3355 => "00000010010011110011010101001101",
			3356 => "11111110100001010011010101001101",
			3357 => "0000000100000000001101001000011000",
			3358 => "0000000100000000000000010000001000",
			3359 => "0000001100000000000100000000000100",
			3360 => "11111111000110110011010101001101",
			3361 => "11111110010001010011010101001101",
			3362 => "0000001100000000001000111000001000",
			3363 => "0000001010000000000111110100000100",
			3364 => "00000010001000100011010101001101",
			3365 => "11111111111101000011010101001101",
			3366 => "0000000111000000001001110000000100",
			3367 => "00000000100000100011010101001101",
			3368 => "00000010011101010011010101001101",
			3369 => "0000001101000000001000000000010000",
			3370 => "0000000111000000001100001000001000",
			3371 => "0000001111000000000010110100000100",
			3372 => "11111110110001000011010101001101",
			3373 => "00000001010001110011010101001101",
			3374 => "0000000111000000001001110000000100",
			3375 => "00000001110000110011010101001101",
			3376 => "00000010110010010011010101001101",
			3377 => "0000000000000000000011010000000100",
			3378 => "00000010110000000011010101001101",
			3379 => "0000000001000000001001111000000100",
			3380 => "00000001001101100011010101001101",
			3381 => "11111111000111100011010101001101",
			3382 => "0000000111000000001100101000011000",
			3383 => "0000000100000000000111011100001100",
			3384 => "0000001010000000001001000100000100",
			3385 => "11111110010011010011010101001101",
			3386 => "0000001100000000000110000100000100",
			3387 => "00000000111010000011010101001101",
			3388 => "00000011011001000011010101001101",
			3389 => "0000000111000000001101111000001000",
			3390 => "0000001110000000001000000000000100",
			3391 => "11111110100100000011010101001101",
			3392 => "00000001100100100011010101001101",
			3393 => "11111110010001100011010101001101",
			3394 => "0000001000000000001001101000000100",
			3395 => "11111110001110110011010101001101",
			3396 => "0000000100000000000110110000011100",
			3397 => "0000001000000000001111001000001100",
			3398 => "0000001001000000001101011000000100",
			3399 => "00000010101100110011010101001101",
			3400 => "0000001100000000001011011100000100",
			3401 => "11111110011101110011010101001101",
			3402 => "00000000110111000011010101001101",
			3403 => "0000000010000000001110111000001000",
			3404 => "0000000100000000001001001100000100",
			3405 => "11111110111110110011010101001101",
			3406 => "00000010100100110011010101001101",
			3407 => "0000000101000000000110111100000100",
			3408 => "11111110100000110011010101001101",
			3409 => "00000001101010000011010101001101",
			3410 => "11111110001110100011010101001101",
			3411 => "0000000111000000001101111010001000",
			3412 => "0000000001000000000000011000011000",
			3413 => "0000000010000000001010010100001000",
			3414 => "0000000101000000001000111100000100",
			3415 => "11111110101011110011011011101001",
			3416 => "00000001001101000011011011101001",
			3417 => "0000000110000000001100011000001000",
			3418 => "0000000010000000000001001000000100",
			3419 => "11111111010101110011011011101001",
			3420 => "11111110010101110011011011101001",
			3421 => "0000001010000000001000101100000100",
			3422 => "00000000011001110011011011101001",
			3423 => "11111110100000100011011011101001",
			3424 => "0000001110000000001101111001000000",
			3425 => "0000000111000000001100001000100000",
			3426 => "0000000011000000001101100000010000",
			3427 => "0000000111000000000111111000001000",
			3428 => "0000000010000000000001000000000100",
			3429 => "00000000011100110011011011101001",
			3430 => "11111110100110000011011011101001",
			3431 => "0000000011000000001011000100000100",
			3432 => "00000001010100010011011011101001",
			3433 => "00000000110101010011011011101001",
			3434 => "0000000010000000000100101000001000",
			3435 => "0000001001000000000110101000000100",
			3436 => "11111110110100000011011011101001",
			3437 => "11111111111110000011011011101001",
			3438 => "0000001001000000001001111000000100",
			3439 => "11111111010100000011011011101001",
			3440 => "00000000101100010011011011101001",
			3441 => "0000001101000000001110110000010000",
			3442 => "0000000010000000001100010100001000",
			3443 => "0000000110000000000001111000000100",
			3444 => "00000010000000100011011011101001",
			3445 => "00000000111000010011011011101001",
			3446 => "0000001000000000000111000100000100",
			3447 => "00000010111100010011011011101001",
			3448 => "00000001011010000011011011101001",
			3449 => "0000000110000000001010011000001000",
			3450 => "0000000010000000000001001000000100",
			3451 => "11111110100110110011011011101001",
			3452 => "11111101000111000011011011101001",
			3453 => "0000000010000000000111011000000100",
			3454 => "00000001111101010011011011101001",
			3455 => "11111110100001110011011011101001",
			3456 => "0000000010000000000011001000010100",
			3457 => "0000000101000000001000000000010000",
			3458 => "0000000111000000001000111000001000",
			3459 => "0000000001000000001001111000000100",
			3460 => "11111111001010000011011011101001",
			3461 => "00000001001101110011011011101001",
			3462 => "0000000110000000001100011000000100",
			3463 => "00000000001111110011011011101001",
			3464 => "00000001111101100011011011101001",
			3465 => "11111110001100000011011011101001",
			3466 => "0000000110000000001100011000001100",
			3467 => "0000000110000000001101111100000100",
			3468 => "11111111100100010011011011101001",
			3469 => "0000001000000000001001101000000100",
			3470 => "00000000110111110011011011101001",
			3471 => "00000011101111100011011011101001",
			3472 => "0000000111000000001001110000001000",
			3473 => "0000000100000000000000010100000100",
			3474 => "11111111101001010011011011101001",
			3475 => "00000000101010000011011011101001",
			3476 => "0000001101000000001000000000000100",
			3477 => "00000001011011110011011011101001",
			3478 => "00000000010001100011011011101001",
			3479 => "0000001000000000001001101000001100",
			3480 => "0000000001000000001011101000001000",
			3481 => "0000000001000000001011101000000100",
			3482 => "11111110011100100011011011101001",
			3483 => "00000010101101010011011011101001",
			3484 => "11111110010110010011011011101001",
			3485 => "0000000100000000000010010000101100",
			3486 => "0000001000000000000001110100011000",
			3487 => "0000001110000000001011110000001100",
			3488 => "0000000100000000001011100000001000",
			3489 => "0000000100000000000010111000000100",
			3490 => "11111111100001000011011011101001",
			3491 => "00000010010010010011011011101001",
			3492 => "11111110001000110011011011101001",
			3493 => "0000000110000000001001111100000100",
			3494 => "11111110010100000011011011101001",
			3495 => "0000000110000000000100101100000100",
			3496 => "00000000100100100011011011101001",
			3497 => "11111110010100100011011011101001",
			3498 => "0000000100000000001101110100001100",
			3499 => "0000000010000000001101001000001000",
			3500 => "0000000010000000001100001100000100",
			3501 => "00000001110101110011011011101001",
			3502 => "00000000101101110011011011101001",
			3503 => "00000010101111110011011011101001",
			3504 => "0000001000000000001010101100000100",
			3505 => "11111110000011000011011011101001",
			3506 => "00000010000010000011011011101001",
			3507 => "0000000100000000000000000000001100",
			3508 => "0000001000000000000000110000000100",
			3509 => "11111110100001110011011011101001",
			3510 => "0000001000000000001010000000000100",
			3511 => "00000001000000000011011011101001",
			3512 => "11111110100111110011011011101001",
			3513 => "11111110010110000011011011101001",
			3514 => "0000000000000000000010101000110000",
			3515 => "0000000110000000000111101000010000",
			3516 => "0000001111000000001000000000000100",
			3517 => "11111110000101110011100010011101",
			3518 => "0000001000000000001000010100000100",
			3519 => "11111111001100110011100010011101",
			3520 => "0000000001000000001110100000000100",
			3521 => "00000000000000000011100010011101",
			3522 => "00000001101010100011100010011101",
			3523 => "0000001000000000000110011100011000",
			3524 => "0000000110000000000111101000001000",
			3525 => "0000001000000000000011101000000100",
			3526 => "00000000000000000011100010011101",
			3527 => "11111100010111110011100010011101",
			3528 => "0000000110000000000001111000001100",
			3529 => "0000000110000000000001111000000100",
			3530 => "11111110100111100011100010011101",
			3531 => "0000000110000000000001111000000100",
			3532 => "00000000000011000011100010011101",
			3533 => "11111111111110100011100010011101",
			3534 => "11111110010000110011100010011101",
			3535 => "0000000110000000001011001100000100",
			3536 => "00000001010011100011100010011101",
			3537 => "11111110111000110011100010011101",
			3538 => "0000001001000000001111001101100000",
			3539 => "0000000111000000000100000000101000",
			3540 => "0000000111000000000100000000011100",
			3541 => "0000000111000000000100000000010000",
			3542 => "0000000111000000001100001000001000",
			3543 => "0000000111000000001100001000000100",
			3544 => "00000000000001010011100010011101",
			3545 => "00000000111000110011100010011101",
			3546 => "0000001011000000000100000000000100",
			3547 => "11111110111010010011100010011101",
			3548 => "11111111110110010011100010011101",
			3549 => "0000001100000000000100010100000100",
			3550 => "11111110100010010011100010011101",
			3551 => "0000001101000000001101111000000100",
			3552 => "00000010100010000011100010011101",
			3553 => "00000000011111000011100010011101",
			3554 => "0000001110000000001110001100001000",
			3555 => "0000000110000000001100011000000100",
			3556 => "00000001101100110011100010011101",
			3557 => "00000010011110110011100010011101",
			3558 => "00000000011011100011100010011101",
			3559 => "0000000111000000001000111000011100",
			3560 => "0000001000000000000110001000001100",
			3561 => "0000000100000000000010111000001000",
			3562 => "0000000000000000000011111100000100",
			3563 => "00000000001011110011100010011101",
			3564 => "11111110000111000011100010011101",
			3565 => "00000001101101000011100010011101",
			3566 => "0000000011000000000000001100001000",
			3567 => "0000000011000000001101111000000100",
			3568 => "11111111000110000011100010011101",
			3569 => "00000001111000000011100010011101",
			3570 => "0000000001000000000010001100000100",
			3571 => "11111101101001110011100010011101",
			3572 => "11111111100011000011100010011101",
			3573 => "0000001111000000001001010000010000",
			3574 => "0000001001000000000111100100001000",
			3575 => "0000001011000000001101100000000100",
			3576 => "11111111010100100011100010011101",
			3577 => "11111100100011110011100010011101",
			3578 => "0000001001000000000111100100000100",
			3579 => "00000010000001100011100010011101",
			3580 => "00000000000000000011100010011101",
			3581 => "0000000001000000001001111000001000",
			3582 => "0000000111000000001001110000000100",
			3583 => "11111101100111010011100010011101",
			3584 => "11111111100101000011100010011101",
			3585 => "00000000000000000011100010011101",
			3586 => "0000001100000000000000101000001100",
			3587 => "0000001100000000000000101000001000",
			3588 => "0000001011000000001101100000000100",
			3589 => "00000010000101100011100010011101",
			3590 => "11111110010000000011100010011101",
			3591 => "00000010111101000011100010011101",
			3592 => "0000001110000000001010111000100000",
			3593 => "0000000010000000000110010000010000",
			3594 => "0000001110000000001101010100001000",
			3595 => "0000001000000000000110001000000100",
			3596 => "11111111011100110011100010011101",
			3597 => "00000001110010100011100010011101",
			3598 => "0000000011000000001001001000000100",
			3599 => "00000011000100000011100010011101",
			3600 => "00000001011011010011100010011101",
			3601 => "0000001110000000001101010100001000",
			3602 => "0000001101000000001001001000000100",
			3603 => "00000001110110100011100010011101",
			3604 => "00000000000000000011100010011101",
			3605 => "0000000110000000001011001100000100",
			3606 => "11111101100010010011100010011101",
			3607 => "00000001000101100011100010011101",
			3608 => "0000001111000000001110101000010000",
			3609 => "0000000100000000000110111000001000",
			3610 => "0000001000000000000001110000000100",
			3611 => "11111111001010100011100010011101",
			3612 => "00000001010110000011100010011101",
			3613 => "0000000111000000001001110000000100",
			3614 => "11111110010011100011100010011101",
			3615 => "11111101000110110011100010011101",
			3616 => "0000000111000000001000111000001000",
			3617 => "0000000010000000001100010000000100",
			3618 => "11111101110010000011100010011101",
			3619 => "00000000011100000011100010011101",
			3620 => "0000000011000000001111011100000100",
			3621 => "00000001000101000011100010011101",
			3622 => "00000000000010110011100010011101",
			3623 => "0000000101000000000100011001111000",
			3624 => "0000000001000000000000011000011100",
			3625 => "0000000110000000001101111100010000",
			3626 => "0000000110000000001101111100001000",
			3627 => "0000000010000000000101110100000100",
			3628 => "11100101110111110011101010010001",
			3629 => "11100100110111110011101010010001",
			3630 => "0000000101000000001000111100000100",
			3631 => "11100101000000110011101010010001",
			3632 => "11100110111001010011101010010001",
			3633 => "0000000011000000001000110000000100",
			3634 => "11101101010100010011101010010001",
			3635 => "0000000010000000000001000000000100",
			3636 => "11101001100100110011101010010001",
			3637 => "11100101000000110011101010010001",
			3638 => "0000000011000000001101100000101000",
			3639 => "0000000110000000000001000100001000",
			3640 => "0000000101000000001001110000000100",
			3641 => "11100100111110000011101010010001",
			3642 => "11100101111110000011101010010001",
			3643 => "0000000011000000001001110000010000",
			3644 => "0000000111000000000111111000001000",
			3645 => "0000001100000000000000110000000100",
			3646 => "11100111101110010011101010010001",
			3647 => "11101011101001000011101010010001",
			3648 => "0000000011000000000100010100000100",
			3649 => "11101101101101000011101010010001",
			3650 => "11101100100001110011101010010001",
			3651 => "0000001101000000001100101100001000",
			3652 => "0000000111000000000000101000000100",
			3653 => "11101000111110010011101010010001",
			3654 => "11101011111000100011101010010001",
			3655 => "0000001001000000000110101000000100",
			3656 => "11101010110110010011101010010001",
			3657 => "11101101001101110011101010010001",
			3658 => "0000000000000000000000110000011000",
			3659 => "0000000110000000001011111100001000",
			3660 => "0000000110000000000001000100000100",
			3661 => "11100100111000110011101010010001",
			3662 => "11100101101010010011101010010001",
			3663 => "0000000110000000001101111100001000",
			3664 => "0000000111000000001011000100000100",
			3665 => "11101000011010110011101010010001",
			3666 => "11101011000011110011101010010001",
			3667 => "0000000000000000000011111100000100",
			3668 => "11100111010100000011101010010001",
			3669 => "11101000110011100011101010010001",
			3670 => "0000000110000000001011001100010000",
			3671 => "0000000000000000000111111000001000",
			3672 => "0000000111000000000000101000000100",
			3673 => "11101000111101110011101010010001",
			3674 => "11101011010110000011101010010001",
			3675 => "0000001001000000001001111000000100",
			3676 => "11101001011100000011101010010001",
			3677 => "11101100111011000011101010010001",
			3678 => "0000000111000000001101100000001000",
			3679 => "0000000011000000001010111100000100",
			3680 => "11101010011111010011101010010001",
			3681 => "11100101010010100011101010010001",
			3682 => "11101001111011000011101010010001",
			3683 => "0000000111000000001110001101001000",
			3684 => "0000000011000000000001101000010100",
			3685 => "0000001100000000000110000100010000",
			3686 => "0000001101000000001001001000001000",
			3687 => "0000000011000000001001110100000100",
			3688 => "11100100111010010011101010010001",
			3689 => "11101001111111100011101010010001",
			3690 => "0000001100000000001100110000000100",
			3691 => "11100100111010000011101010010001",
			3692 => "11100101111110000011101010010001",
			3693 => "11101000100110110011101010010001",
			3694 => "0000000110000000001001100100011000",
			3695 => "0000000000000000000001110100001000",
			3696 => "0000000111000000000101101100000100",
			3697 => "11100101111110000011101010010001",
			3698 => "11100100111010000011101010010001",
			3699 => "0000001000000000000010101000001000",
			3700 => "0000000111000000001001110000000100",
			3701 => "11100110001100000011101010010001",
			3702 => "11101011101111110011101010010001",
			3703 => "0000000000000000001100110000000100",
			3704 => "11100101111110000011101010010001",
			3705 => "11100101000001110011101010010001",
			3706 => "0000000111000000000110000100010000",
			3707 => "0000000001000000000111100100001000",
			3708 => "0000000000000000000011010000000100",
			3709 => "11101000100110110011101010010001",
			3710 => "11100101001100110011101010010001",
			3711 => "0000001000000000000111000100000100",
			3712 => "11100100111000100011101010010001",
			3713 => "11100101100010110011101010010001",
			3714 => "0000000010000000001000100000000100",
			3715 => "11101110010000100011101010010001",
			3716 => "0000000011000000001101000100000100",
			3717 => "11100100111101010011101010010001",
			3718 => "11101000010001100011101010010001",
			3719 => "0000001001000000001000010100110100",
			3720 => "0000000111000000001101111000011000",
			3721 => "0000001111000000000110010000010000",
			3722 => "0000001101000000001000011000001000",
			3723 => "0000001111000000001110101100000100",
			3724 => "11100100111001110011101010010001",
			3725 => "11101010011111010011101010010001",
			3726 => "0000000011000000000000110100000100",
			3727 => "11100100111011010011101010010001",
			3728 => "11100101110100000011101010010001",
			3729 => "0000001100000000001100110000000100",
			3730 => "11100100111101110011101010010001",
			3731 => "11101100001001000011101010010001",
			3732 => "0000001000000000001001101000001100",
			3733 => "0000001100000000000110000100001000",
			3734 => "0000001100000000000110000100000100",
			3735 => "11100100111100100011101010010001",
			3736 => "11100110001010010011101010010001",
			3737 => "11100100110111110011101010010001",
			3738 => "0000000000000000001000111100001000",
			3739 => "0000000001000000001101101000000100",
			3740 => "11101101100110010011101010010001",
			3741 => "11100101011001110011101010010001",
			3742 => "0000001010000000000001010100000100",
			3743 => "11100101110010100011101010010001",
			3744 => "11100100111000000011101010010001",
			3745 => "0000000000000000000011010000000100",
			3746 => "11100100111111000011101010010001",
			3747 => "11101001100011000011101010010001",
			3748 => "0000000100000000000110110010101000",
			3749 => "0000000001000000001011101001110100",
			3750 => "0000000001000000001001111001000000",
			3751 => "0000001110000000001101111000100000",
			3752 => "0000001001000000000111100100010000",
			3753 => "0000000011000000001101111000001000",
			3754 => "0000001001000000000110101000000100",
			3755 => "11111111111111010011110000010101",
			3756 => "00000000010011010011110000010101",
			3757 => "0000000010000000000110010000000100",
			3758 => "11111111000101010011110000010101",
			3759 => "00000000100110100011110000010101",
			3760 => "0000000010000000001110101000001000",
			3761 => "0000001000000000000101000100000100",
			3762 => "00000000100100100011110000010101",
			3763 => "11111110000111010011110000010101",
			3764 => "0000001010000000001000100100000100",
			3765 => "00000001100011110011110000010101",
			3766 => "00000000011011110011110000010101",
			3767 => "0000001011000000001100001000010000",
			3768 => "0000000111000000001011000100001000",
			3769 => "0000001101000000001100101100000100",
			3770 => "00000001000011100011110000010101",
			3771 => "11111110001100110011110000010101",
			3772 => "0000000110000000001100011000000100",
			3773 => "00000011101101110011110000010101",
			3774 => "00000000100101010011110000010101",
			3775 => "0000000001000000001100110100001000",
			3776 => "0000001111000000000001000000000100",
			3777 => "11111101011011000011110000010101",
			3778 => "00000000110110100011110000010101",
			3779 => "0000000010000000000010000000000100",
			3780 => "11111111100010100011110000010101",
			3781 => "00000000000011010011110000010101",
			3782 => "0000001110000000001010111000011000",
			3783 => "0000001000000000001011010100001100",
			3784 => "0000000111000000001000111000000100",
			3785 => "00000001110001000011110000010101",
			3786 => "0000001110000000000000001100000100",
			3787 => "00000000111111100011110000010101",
			3788 => "11111110011100110011110000010101",
			3789 => "0000001011000000001101100000000100",
			3790 => "00000000001010000011110000010101",
			3791 => "0000000110000000001010011000000100",
			3792 => "00000010100110010011110000010101",
			3793 => "00000001101011000011110000010101",
			3794 => "0000000111000000001101100000010000",
			3795 => "0000000001000000000110101000001000",
			3796 => "0000001100000000000000101000000100",
			3797 => "00000001111110010011110000010101",
			3798 => "11111111110011010011110000010101",
			3799 => "0000000100000000001110000000000100",
			3800 => "11111111110110100011110000010101",
			3801 => "11111110000110110011110000010101",
			3802 => "0000001000000000001010110000000100",
			3803 => "11111110100000000011110000010101",
			3804 => "0000001101000000000000011100000100",
			3805 => "00000000100001010011110000010101",
			3806 => "00000001111010010011110000010101",
			3807 => "0000001000000000000110001000010100",
			3808 => "0000001100000000001011011100010000",
			3809 => "0000000100000000001000001000000100",
			3810 => "11111110011000010011110000010101",
			3811 => "0000000100000000001000001000001000",
			3812 => "0000001000000000001100000100000100",
			3813 => "00000000000000000011110000010101",
			3814 => "00000000111101000011110000010101",
			3815 => "11111110101110000011110000010101",
			3816 => "00000000011111000011110000010101",
			3817 => "0000001011000000001000000000000100",
			3818 => "11111110011010100011110000010101",
			3819 => "0000000110000000001001111100010000",
			3820 => "0000000100000000001011100000001000",
			3821 => "0000001010000000001100011100000100",
			3822 => "00000001011011010011110000010101",
			3823 => "11111111101110110011110000010101",
			3824 => "0000001010000000000001010100000100",
			3825 => "11111110100001110011110000010101",
			3826 => "00000001000100100011110000010101",
			3827 => "0000001110000000000011010100001000",
			3828 => "0000000100000000001110111000000100",
			3829 => "11111111011100000011110000010101",
			3830 => "00000001010011010011110000010101",
			3831 => "11111111111011110011110000010101",
			3832 => "0000000110000000001011001100000100",
			3833 => "11111110010111100011110000010101",
			3834 => "0000000010000000000010000100001000",
			3835 => "0000000001000000001110011100000100",
			3836 => "11111111111001110011110000010101",
			3837 => "00000001011111110011110000010101",
			3838 => "0000001010000000001100000100001100",
			3839 => "0000001000000000001111000100000100",
			3840 => "11111110110010000011110000010101",
			3841 => "0000000100000000000101100000000100",
			3842 => "00000001110001100011110000010101",
			3843 => "00000000000000000011110000010101",
			3844 => "11111110100110010011110000010101",
			3845 => "0000001100000000000000001110010000",
			3846 => "0000000100000000000110110001111000",
			3847 => "0000001110000000001000111100111100",
			3848 => "0000001001000000000110101000011100",
			3849 => "0000001011000000000100000000010000",
			3850 => "0000001101000000001100101100001000",
			3851 => "0000000011000000001001110000000100",
			3852 => "00000000010011010011110110011001",
			3853 => "11111111100000100011110110011001",
			3854 => "0000000010000000000111111100000100",
			3855 => "00000000010010010011110110011001",
			3856 => "00000001011000100011110110011001",
			3857 => "0000001010000000001100011100001000",
			3858 => "0000000010000000000101110000000100",
			3859 => "11111111000001100011110110011001",
			3860 => "11111100111000000011110110011001",
			3861 => "00000001101010100011110110011001",
			3862 => "0000000001000000001100110100010000",
			3863 => "0000001110000000001100001000001000",
			3864 => "0000000101000000000110000100000100",
			3865 => "00000000011010010011110110011001",
			3866 => "00000010100000010011110110011001",
			3867 => "0000001111000000001011110100000100",
			3868 => "11111111111111000011110110011001",
			3869 => "00000010101001010011110110011001",
			3870 => "0000001001000000000111100100001000",
			3871 => "0000001011000000001100001000000100",
			3872 => "11111111000000010011110110011001",
			3873 => "00000000011101010011110110011001",
			3874 => "0000001111000000000101100100000100",
			3875 => "00000000001001010011110110011001",
			3876 => "00000001000111110011110110011001",
			3877 => "0000001111000000000010001000011100",
			3878 => "0000001001000000001101101000010000",
			3879 => "0000001011000000000000101000001000",
			3880 => "0000001100000000000111111000000100",
			3881 => "00000011010010110011110110011001",
			3882 => "11111111110100100011110110011001",
			3883 => "0000001000000000000001010100000100",
			3884 => "11111110110001100011110110011001",
			3885 => "11111101101010100011110110011001",
			3886 => "0000000101000000001101111000000100",
			3887 => "11111101110001000011110110011001",
			3888 => "0000001110000000000101101100000100",
			3889 => "00000000110101100011110110011001",
			3890 => "11111110101101110011110110011001",
			3891 => "0000001001000000001101101000010000",
			3892 => "0000000010000000000010000000001000",
			3893 => "0000001110000000000101101100000100",
			3894 => "11111111111001110011110110011001",
			3895 => "11111110111000110011110110011001",
			3896 => "0000000101000000001010111100000100",
			3897 => "00000000110000010011110110011001",
			3898 => "11111110000010100011110110011001",
			3899 => "0000001110000000001101111000001000",
			3900 => "0000001101000000001101111000000100",
			3901 => "11111110010010110011110110011001",
			3902 => "00000000110110000011110110011001",
			3903 => "0000001001000000001111001100000100",
			3904 => "11111111101101110011110110011001",
			3905 => "00000000010101100011110110011001",
			3906 => "0000001011000000000100011000010100",
			3907 => "0000000001000000001100100000000100",
			3908 => "11111110011010000011110110011001",
			3909 => "0000001111000000001001001000000100",
			3910 => "00000000001101100011110110011001",
			3911 => "0000000010000000001010001000000100",
			3912 => "11111101011101000011110110011001",
			3913 => "0000000010000000001001100000000100",
			3914 => "00000001000101010011110110011001",
			3915 => "11111110001010000011110110011001",
			3916 => "00000001101110000011110110011001",
			3917 => "0000001000000000001001101000001000",
			3918 => "0000001110000000001010001100000100",
			3919 => "00000001011001110011110110011001",
			3920 => "11111110011000110011110110011001",
			3921 => "0000000100000000000011111000101000",
			3922 => "0000001110000000001100111000010100",
			3923 => "0000000010000000001011110000001100",
			3924 => "0000001001000000001011001100001000",
			3925 => "0000000100000000001101110100000100",
			3926 => "00000001101010000011110110011001",
			3927 => "00000000000000000011110110011001",
			3928 => "11111110101101000011110110011001",
			3929 => "0000000010000000000101000000000100",
			3930 => "00000010011111100011110110011001",
			3931 => "00000000100101010011110110011001",
			3932 => "0000001100000000001011011100001100",
			3933 => "0000001000000000000110001000000100",
			3934 => "11111110011011010011110110011001",
			3935 => "0000000000000000000000111000000100",
			3936 => "00000001000001110011110110011001",
			3937 => "11111110111100110011110110011001",
			3938 => "0000000001000000001100011000000100",
			3939 => "11111110101001010011110110011001",
			3940 => "00000010010000000011110110011001",
			3941 => "11111110011001100011110110011001",
			3942 => "0000000101000000000100011010101100",
			3943 => "0000001010000000001001000101011100",
			3944 => "0000001011000000000100010100011100",
			3945 => "0000000000000000001111000100001000",
			3946 => "0000001110000000001010000000000100",
			3947 => "11111100101010010011111101111101",
			3948 => "11111110101011010011111101111101",
			3949 => "0000000100000000001100001100000100",
			3950 => "00000001010101110011111101111101",
			3951 => "0000001110000000000011010000001000",
			3952 => "0000001010000000001000010100000100",
			3953 => "11111101000111000011111101111101",
			3954 => "00000000011100100011111101111101",
			3955 => "0000001000000000001001101000000100",
			3956 => "11111010110001110011111101111101",
			3957 => "11111110000110100011111101111101",
			3958 => "0000000010000000000100101000100000",
			3959 => "0000000100000000001100001100010000",
			3960 => "0000001110000000000000110000001000",
			3961 => "0000000100000000000101000000000100",
			3962 => "00000001101100000011111101111101",
			3963 => "11111111100110010011111101111101",
			3964 => "0000001001000000001001111000000100",
			3965 => "11111101110111000011111101111101",
			3966 => "00000000001010100011111101111101",
			3967 => "0000001111000000001011011100001000",
			3968 => "0000000010000000001001010000000100",
			3969 => "00000000011111110011111101111101",
			3970 => "11111101011100000011111101111101",
			3971 => "0000000010000000001111010000000100",
			3972 => "00000000011011110011111101111101",
			3973 => "00000001101010100011111101111101",
			3974 => "0000001000000000001001101000010000",
			3975 => "0000001010000000001000010100001000",
			3976 => "0000000100000000001110000000000100",
			3977 => "11111111110110100011111101111101",
			3978 => "00000001111010110011111101111101",
			3979 => "0000000010000000000011001000000100",
			3980 => "11111110111000100011111101111101",
			3981 => "00000010000001110011111101111101",
			3982 => "0000000110000000001101111100001000",
			3983 => "0000000101000000000110000100000100",
			3984 => "00000010101001110011111101111101",
			3985 => "11111111101001100011111101111101",
			3986 => "0000000111000000001100001000000100",
			3987 => "00000100000100110011111101111101",
			3988 => "00000001001111000011111101111101",
			3989 => "0000000100000000000011001100011000",
			3990 => "0000000000000000000000110000010000",
			3991 => "0000000000000000001111000100000100",
			3992 => "00000010111111110011111101111101",
			3993 => "0000000001000000000110000000000100",
			3994 => "00000001111110010011111101111101",
			3995 => "0000000101000000001101010100000100",
			3996 => "11111111011000110011111101111101",
			3997 => "00000000011000010011111101111101",
			3998 => "0000000010000000001001011100000100",
			3999 => "00000011111101010011111101111101",
			4000 => "00000001011111010011111101111101",
			4001 => "0000000110000000000001111000011000",
			4002 => "0000000111000000001011000100010000",
			4003 => "0000000111000000000100010100001000",
			4004 => "0000001000000000000110001000000100",
			4005 => "00000001100010110011111101111101",
			4006 => "11111110011101010011111101111101",
			4007 => "0000001111000000001001110100000100",
			4008 => "00000000000000010011111101111101",
			4009 => "11111011110011010011111101111101",
			4010 => "0000000101000000000011011100000100",
			4011 => "11111101001110110011111101111101",
			4012 => "00000001110010110011111101111101",
			4013 => "0000001010000000000001010000010000",
			4014 => "0000001001000000000111100100001000",
			4015 => "0000001110000000001100001000000100",
			4016 => "00000000100101110011111101111101",
			4017 => "11111111111001100011111101111101",
			4018 => "0000001100000000001000111000000100",
			4019 => "00000001010100010011111101111101",
			4020 => "11111110111101100011111101111101",
			4021 => "0000000100000000001001001100001000",
			4022 => "0000001001000000001011101000000100",
			4023 => "11111111001111010011111101111101",
			4024 => "00000000110101110011111101111101",
			4025 => "0000001100000000001110111100000100",
			4026 => "11111111100111100011111101111101",
			4027 => "00000000010100000011111101111101",
			4028 => "0000001000000000000001010100011000",
			4029 => "0000000101000000001000000000010100",
			4030 => "0000000111000000001101100000001100",
			4031 => "0000000110000000001101111100001000",
			4032 => "0000001100000000001000111000000100",
			4033 => "00000000111001000011111101111101",
			4034 => "00000000000000000011111101111101",
			4035 => "11111110000010110011111101111101",
			4036 => "0000001111000000001010111000000100",
			4037 => "11111111010110010011111101111101",
			4038 => "00000010010101000011111101111101",
			4039 => "11111110011000010011111101111101",
			4040 => "0000000100000000000000000000101100",
			4041 => "0000001011000000000110000100010000",
			4042 => "0000000000000000000010111100000100",
			4043 => "00000001000100100011111101111101",
			4044 => "0000001001000000001111001100000100",
			4045 => "11111100101111100011111101111101",
			4046 => "0000000010000000001100000000000100",
			4047 => "11111111001110110011111101111101",
			4048 => "11111101111010110011111101111101",
			4049 => "0000001110000000000001011100001100",
			4050 => "0000001000000000000001010100000100",
			4051 => "00000011100010100011111101111101",
			4052 => "0000001010000000001100000100000100",
			4053 => "11111111111010010011111101111101",
			4054 => "00000001111101000011111101111101",
			4055 => "0000000110000000001001111100001000",
			4056 => "0000001100000000001011011100000100",
			4057 => "11111110011001110011111101111101",
			4058 => "00000000100111010011111101111101",
			4059 => "0000001111000000000000010100000100",
			4060 => "00000000110011110011111101111101",
			4061 => "11111111001110010011111101111101",
			4062 => "11111110011010010011111101111101",
			4063 => "0000001001000000001001111010001000",
			4064 => "0000000101000000001101100001000100",
			4065 => "0000000101000000000011011100111100",
			4066 => "0000000010000000001001010000011100",
			4067 => "0000000011000000001100001000010000",
			4068 => "0000000100000000000000010100001000",
			4069 => "0000001000000000001100000100000100",
			4070 => "11111110000010010100000110101001",
			4071 => "00000000010111010100000110101001",
			4072 => "0000001010000000001010110000000100",
			4073 => "11111110001110010100000110101001",
			4074 => "11111111101111000100000110101001",
			4075 => "0000001000000000001011010100001000",
			4076 => "0000000011000000000100000000000100",
			4077 => "00000001000010010100000110101001",
			4078 => "11111101111110110100000110101001",
			4079 => "11111101110101110100000110101001",
			4080 => "0000001010000000001010110000010000",
			4081 => "0000001010000000001010110000001000",
			4082 => "0000001101000000001001110000000100",
			4083 => "11111110010011000100000110101001",
			4084 => "00000000101100010100000110101001",
			4085 => "0000000111000000001110111100000100",
			4086 => "11111111110111110100000110101001",
			4087 => "00000010000101110100000110101001",
			4088 => "0000000110000000001101111100001000",
			4089 => "0000000010000000001110010000000100",
			4090 => "11111111101011100100000110101001",
			4091 => "11111101101110110100000110101001",
			4092 => "0000000010000000001110010000000100",
			4093 => "00000000001101000100000110101001",
			4094 => "00000001101000010100000110101001",
			4095 => "0000000100000000001011100000000100",
			4096 => "00000001110010010100000110101001",
			4097 => "11111111110111010100000110101001",
			4098 => "0000000110000000001101111100100100",
			4099 => "0000001101000000001101100000001100",
			4100 => "0000001100000000000100010100001000",
			4101 => "0000000100000000000101010100000100",
			4102 => "11111110100110010100000110101001",
			4103 => "00000001100011110100000110101001",
			4104 => "11111101001110010100000110101001",
			4105 => "0000000000000000000011010000001100",
			4106 => "0000000011000000001100001000000100",
			4107 => "00000001100001100100000110101001",
			4108 => "0000000010000000001110101000000100",
			4109 => "11111101111100000100000110101001",
			4110 => "00000000000000000100000110101001",
			4111 => "0000000010000000001100010100001000",
			4112 => "0000001001000000001100110100000100",
			4113 => "00000000000000000100000110101001",
			4114 => "00000001110101000100000110101001",
			4115 => "11111111110001110100000110101001",
			4116 => "0000001110000000000000111000010100",
			4117 => "0000001110000000000011111100010000",
			4118 => "0000001011000000000100010100001000",
			4119 => "0000000011000000000100010100000100",
			4120 => "11111111111010100100000110101001",
			4121 => "11111101100010110100000110101001",
			4122 => "0000000110000000001101111100000100",
			4123 => "00000001011110010100000110101001",
			4124 => "11111111011010000100000110101001",
			4125 => "00000000111010000100000110101001",
			4126 => "0000001110000000000111111000001000",
			4127 => "0000000010000000001010001000000100",
			4128 => "11111110011100010100000110101001",
			4129 => "11111101000101110100000110101001",
			4130 => "11111111111101110100000110101001",
			4131 => "0000000011000000000101101101001100",
			4132 => "0000000011000000000101101100110100",
			4133 => "0000000011000000001100110000100000",
			4134 => "0000000011000000001100110000010000",
			4135 => "0000000011000000001100110000001000",
			4136 => "0000001101000000001101111000000100",
			4137 => "00000000001000000100000110101001",
			4138 => "00000001111000100100000110101001",
			4139 => "0000001100000000000111111000000100",
			4140 => "00000001011110000100000110101001",
			4141 => "11111110110001110100000110101001",
			4142 => "0000001010000000001100011100001000",
			4143 => "0000000101000000000110000100000100",
			4144 => "00000000100011100100000110101001",
			4145 => "00000010001001100100000110101001",
			4146 => "0000001000000000000010101000000100",
			4147 => "11111101101111010100000110101001",
			4148 => "00000001100001110100000110101001",
			4149 => "0000001010000000001001000100001000",
			4150 => "0000001101000000001100101100000100",
			4151 => "00000001011010110100000110101001",
			4152 => "11111111000111000100000110101001",
			4153 => "0000000010000000001110010000001000",
			4154 => "0000001101000000001110001100000100",
			4155 => "11111110000010100100000110101001",
			4156 => "11111111010001010100000110101001",
			4157 => "11111111111001010100000110101001",
			4158 => "0000001011000000001100001000001100",
			4159 => "0000000111000000001011000100000100",
			4160 => "00000000111010110100000110101001",
			4161 => "0000001110000000001011000100000100",
			4162 => "00000001000110100100000110101001",
			4163 => "00000010011000100100000110101001",
			4164 => "0000001001000000000111100100000100",
			4165 => "11111111101010000100000110101001",
			4166 => "0000000111000000001100001000000100",
			4167 => "00000000011000010100000110101001",
			4168 => "00000001110000000100000110101001",
			4169 => "0000001101000000000101101100001100",
			4170 => "0000001110000000001001110000001000",
			4171 => "0000000010000000001110010000000100",
			4172 => "11111111010110100100000110101001",
			4173 => "11111101011010100100000110101001",
			4174 => "00000000101110100100000110101001",
			4175 => "0000000011000000000110000100011100",
			4176 => "0000000011000000000101101100010000",
			4177 => "0000001010000000001001000100001000",
			4178 => "0000001011000000001100001000000100",
			4179 => "11111110110011000100000110101001",
			4180 => "00000001101100010100000110101001",
			4181 => "0000000000000000000000110000000100",
			4182 => "11111110100001000100000110101001",
			4183 => "00000000001001000100000110101001",
			4184 => "0000001101000000001101111000001000",
			4185 => "0000000010000000000100101000000100",
			4186 => "11111110110001110100000110101001",
			4187 => "11111101110011100100000110101001",
			4188 => "00000000101100110100000110101001",
			4189 => "0000000011000000000110000100001100",
			4190 => "0000001010000000001100011100001000",
			4191 => "0000000010000000001001010000000100",
			4192 => "00000000101111110100000110101001",
			4193 => "00000010010000110100000110101001",
			4194 => "11111110100110110100000110101001",
			4195 => "0000001100000000000000101000001000",
			4196 => "0000001100000000000000101000000100",
			4197 => "11111111111010100100000110101001",
			4198 => "11111111010100100100000110101001",
			4199 => "0000000111000000001100001000000100",
			4200 => "00000000010111110100000110101001",
			4201 => "11111111111110110100000110101001",
			4202 => "0000000011000000000100000010001100",
			4203 => "0000000100000000000011010101000100",
			4204 => "0000000000000000000100010100110100",
			4205 => "0000000011000000000100000000100000",
			4206 => "0000000011000000001100001000010000",
			4207 => "0000000110000000000100110100001000",
			4208 => "0000001110000000000011111100000100",
			4209 => "00000000000110110100001111001101",
			4210 => "00000000110110010100001111001101",
			4211 => "0000001001000000001001111000000100",
			4212 => "11111110010100000100001111001101",
			4213 => "11111111111011000100001111001101",
			4214 => "0000000100000000001010110100001000",
			4215 => "0000000111000000001011000100000100",
			4216 => "11111101010001010100001111001101",
			4217 => "00000000100001010100001111001101",
			4218 => "0000001110000000000011010000000100",
			4219 => "00000000000110110100001111001101",
			4220 => "00000001110010010100001111001101",
			4221 => "0000001011000000000100010100001100",
			4222 => "0000000100000000001010110100000100",
			4223 => "00000001101011010100001111001101",
			4224 => "0000000100000000000000010100000100",
			4225 => "11111110110000000100001111001101",
			4226 => "00000000001110000100001111001101",
			4227 => "0000001001000000000110101000000100",
			4228 => "00000001111010110100001111001101",
			4229 => "00000000000000000100001111001101",
			4230 => "0000000110000000000100110100000100",
			4231 => "00000001110010000100001111001101",
			4232 => "0000001101000000001101100000000100",
			4233 => "11111110110000100100001111001101",
			4234 => "0000001101000000001100101100000100",
			4235 => "00000001011100110100001111001101",
			4236 => "00000000000000000100001111001101",
			4237 => "0000000100000000000011110100011000",
			4238 => "0000000001000000001110100000010100",
			4239 => "0000000110000000001101111100000100",
			4240 => "11111101011000000100001111001101",
			4241 => "0000000011000000001100001000001000",
			4242 => "0000001011000000000100010100000100",
			4243 => "11111111001000110100001111001101",
			4244 => "00000000110100000100001111001101",
			4245 => "0000000110000000000100110100000100",
			4246 => "11111111100110010100001111001101",
			4247 => "11111100111110010100001111001101",
			4248 => "00000001011101110100001111001101",
			4249 => "0000000001000000000110000000011100",
			4250 => "0000001111000000001110110000001100",
			4251 => "0000000100000000000110110000000100",
			4252 => "00000001011010000100001111001101",
			4253 => "0000000110000000001011001100000100",
			4254 => "11111111000011010100001111001101",
			4255 => "00000000000000000100001111001101",
			4256 => "0000001011000000001110111100001000",
			4257 => "0000000101000000001000111000000100",
			4258 => "11111111010001010100001111001101",
			4259 => "00000001010111000100001111001101",
			4260 => "0000001100000000000100010100000100",
			4261 => "11111110000010010100001111001101",
			4262 => "00000000110010110100001111001101",
			4263 => "0000000001000000000110000000001000",
			4264 => "0000000000000000001000111000000100",
			4265 => "00000001110000100100001111001101",
			4266 => "11111111010110000100001111001101",
			4267 => "0000001011000000000111111000000100",
			4268 => "11111101111110100100001111001101",
			4269 => "0000001111000000000101100100000100",
			4270 => "11111111111010000100001111001101",
			4271 => "00000001011110100100001111001101",
			4272 => "0000001001000000000010001100011100",
			4273 => "0000000110000000000001111000001100",
			4274 => "0000001110000000000000110000001000",
			4275 => "0000000100000000001101110100000100",
			4276 => "00000001110100000100001111001101",
			4277 => "00000000000000000100001111001101",
			4278 => "00000000000000000100001111001101",
			4279 => "0000000110000000001101111100000100",
			4280 => "11111101100001110100001111001101",
			4281 => "0000001110000000001010000000001000",
			4282 => "0000001111000000000110110100000100",
			4283 => "00000010001110000100001111001101",
			4284 => "11111111101100100100001111001101",
			4285 => "11111110100100010100001111001101",
			4286 => "0000001111000000000001011000110000",
			4287 => "0000001001000000000110101000010100",
			4288 => "0000000001000000001110100000010000",
			4289 => "0000001110000000000000110000001000",
			4290 => "0000000111000000000100010100000100",
			4291 => "00000000000100110100001111001101",
			4292 => "00000001110011110100001111001101",
			4293 => "0000000101000000000101101100000100",
			4294 => "11111110011101010100001111001101",
			4295 => "00000000100111000100001111001101",
			4296 => "11111101011000000100001111001101",
			4297 => "0000001101000000001110001100010000",
			4298 => "0000001111000000000000011100001000",
			4299 => "0000001000000000001001101000000100",
			4300 => "00000001011000100100001111001101",
			4301 => "00000000000001000100001111001101",
			4302 => "0000000011000000000011011100000100",
			4303 => "11111110001100000100001111001101",
			4304 => "11111111101011110100001111001101",
			4305 => "0000001110000000000000110000000100",
			4306 => "11111101101010000100001111001101",
			4307 => "0000000100000000001010110100000100",
			4308 => "11111111000111110100001111001101",
			4309 => "00000001001001110100001111001101",
			4310 => "0000001000000000000110001000100000",
			4311 => "0000000100000000000011001100010000",
			4312 => "0000001110000000000111111000001000",
			4313 => "0000001101000000000110000100000100",
			4314 => "11111101111110100100001111001101",
			4315 => "00000000101110110100001111001101",
			4316 => "0000000101000000001101111000000100",
			4317 => "00000000010000110100001111001101",
			4318 => "11111111110111110100001111001101",
			4319 => "0000001111000000001010010100001000",
			4320 => "0000001000000000001001101000000100",
			4321 => "00000010000101010100001111001101",
			4322 => "00000000000011000100001111001101",
			4323 => "0000001101000000001100101000000100",
			4324 => "00000010000011000100001111001101",
			4325 => "00000000100101000100001111001101",
			4326 => "0000000111000000000111111000001100",
			4327 => "0000000101000000001100110000001000",
			4328 => "0000000101000000001101100000000100",
			4329 => "00000000011100100100001111001101",
			4330 => "00000010010111100100001111001101",
			4331 => "11111111001000000100001111001101",
			4332 => "0000000000000000000100010100001000",
			4333 => "0000001000000000000111000100000100",
			4334 => "11111111111011100100001111001101",
			4335 => "11111111100101010100001111001101",
			4336 => "0000000100000000000000010100000100",
			4337 => "00000001110101100100001111001101",
			4338 => "00000000000011000100001111001101",
			4339 => "0000000010000000000010110101110000",
			4340 => "0000000010000000000001001000100100",
			4341 => "0000000000000000001000110000010000",
			4342 => "0000001011000000001011000100000100",
			4343 => "11111101110110110100011000100001",
			4344 => "0000001100000000000100010100001000",
			4345 => "0000000000000000000110001000000100",
			4346 => "11111111110101110100011000100001",
			4347 => "00000001010010000100011000100001",
			4348 => "11111110011100010100011000100001",
			4349 => "0000001100000000001010000000010000",
			4350 => "0000000111000000000111111000001000",
			4351 => "0000000111000000001010000000000100",
			4352 => "00000000000111100100011000100001",
			4353 => "11111110110011000100011000100001",
			4354 => "0000000001000000001100100000000100",
			4355 => "00000000000000000100011000100001",
			4356 => "00000001000011100100011000100001",
			4357 => "00000001101101100100011000100001",
			4358 => "0000001011000000000100010100101000",
			4359 => "0000000111000000000111111000011100",
			4360 => "0000000111000000001110111100001100",
			4361 => "0000000110000000000001111000000100",
			4362 => "00000000000000000100011000100001",
			4363 => "0000001010000000001100000100000100",
			4364 => "00000001010101010100011000100001",
			4365 => "00000000000000000100011000100001",
			4366 => "0000001100000000001010000000001000",
			4367 => "0000000010000000001110101100000100",
			4368 => "00000000000000000100011000100001",
			4369 => "00000000001000100100011000100001",
			4370 => "0000000110000000000001111000000100",
			4371 => "00000000000000000100011000100001",
			4372 => "11111101001100110100011000100001",
			4373 => "0000001111000000000110100100001000",
			4374 => "0000000001000000000000011000000100",
			4375 => "00000000000000000100011000100001",
			4376 => "00000001101001110100011000100001",
			4377 => "11111111110110010100011000100001",
			4378 => "0000000101000000001100110000010000",
			4379 => "0000000010000000000000110100000100",
			4380 => "00000000000111110100011000100001",
			4381 => "0000001100000000000100010100001000",
			4382 => "0000000000000000001110111100000100",
			4383 => "11111101111010110100011000100001",
			4384 => "11111100011100000100011000100001",
			4385 => "11111111000001100100011000100001",
			4386 => "0000000000000000000000111000010000",
			4387 => "0000000110000000000111101000001000",
			4388 => "0000001111000000001111011100000100",
			4389 => "00000001011110010100011000100001",
			4390 => "11111111101001100100011000100001",
			4391 => "0000001001000000000110101000000100",
			4392 => "11111101001101110100011000100001",
			4393 => "11111111010011100100011000100001",
			4394 => "00000001101000010100011000100001",
			4395 => "0000000000000000000010111101011000",
			4396 => "0000000100000000000110001100110100",
			4397 => "0000001010000000000110011000100000",
			4398 => "0000001010000000001000010100010000",
			4399 => "0000001000000000001001101000001000",
			4400 => "0000000100000000001100001100000100",
			4401 => "00000000001101010100011000100001",
			4402 => "11111110001011010100011000100001",
			4403 => "0000001011000000001100001000000100",
			4404 => "00000010011101110100011000100001",
			4405 => "00000000011011110100011000100001",
			4406 => "0000000100000000001000110100001000",
			4407 => "0000000001000000000010001100000100",
			4408 => "00000010101000010100011000100001",
			4409 => "00000000000010000100011000100001",
			4410 => "0000001100000000000100000000000100",
			4411 => "11111110011011100100011000100001",
			4412 => "00000000000000000100011000100001",
			4413 => "0000000101000000000100011000001000",
			4414 => "0000000001000000001001111000000100",
			4415 => "00000000101111100100011000100001",
			4416 => "00000010011011100100011000100001",
			4417 => "0000000111000000001101100000000100",
			4418 => "11111110011110000100011000100001",
			4419 => "0000001000000000001011010100000100",
			4420 => "11111110111010010100011000100001",
			4421 => "00000001011011100100011000100001",
			4422 => "0000000001000000000110000000000100",
			4423 => "11111101011010110100011000100001",
			4424 => "0000000000000000000010011000010000",
			4425 => "0000001000000000001001101000001000",
			4426 => "0000000000000000001111000100000100",
			4427 => "11111111110001000100011000100001",
			4428 => "11111011110111010100011000100001",
			4429 => "0000001100000000001001110100000100",
			4430 => "00000000000000000100011000100001",
			4431 => "00000001100010010100011000100001",
			4432 => "0000001100000000000100000000001000",
			4433 => "0000001011000000001000111100000100",
			4434 => "00000000111100110100011000100001",
			4435 => "00000010101000100100011000100001",
			4436 => "0000001000000000001001101000000100",
			4437 => "00000001001111000100011000100001",
			4438 => "11111110110110000100011000100001",
			4439 => "0000000011000000001100001000111000",
			4440 => "0000000100000000001110111000011000",
			4441 => "0000001011000000001011000100010000",
			4442 => "0000000111000000000100010100001000",
			4443 => "0000000110000000000001111000000100",
			4444 => "11111111100011010100011000100001",
			4445 => "00000001010110010100011000100001",
			4446 => "0000000100000000001101001000000100",
			4447 => "00000001110001100100011000100001",
			4448 => "11111111001010000100011000100001",
			4449 => "0000001011000000000000101000000100",
			4450 => "00000001110111100100011000100001",
			4451 => "00000000010011110100011000100001",
			4452 => "0000000000000000000111111000010000",
			4453 => "0000001100000000001010000000001000",
			4454 => "0000001011000000000111111000000100",
			4455 => "11111110100001010100011000100001",
			4456 => "00000001101111100100011000100001",
			4457 => "0000000110000000000001111000000100",
			4458 => "11111111111111000100011000100001",
			4459 => "11111110001011000100011000100001",
			4460 => "0000001100000000000111111000001000",
			4461 => "0000001100000000000111111000000100",
			4462 => "00000000011101010100011000100001",
			4463 => "11111110100011100100011000100001",
			4464 => "0000001100000000000111111000000100",
			4465 => "00000001100001010100011000100001",
			4466 => "00000000001011110100011000100001",
			4467 => "0000001000000000001001101000011000",
			4468 => "0000000011000000001101111000001100",
			4469 => "0000001100000000000000101000001000",
			4470 => "0000001011000000001011000100000100",
			4471 => "00000000101100010100011000100001",
			4472 => "11111110111001000100011000100001",
			4473 => "00000001111110100100011000100001",
			4474 => "0000000011000000000100011000001000",
			4475 => "0000000000000000000010111100000100",
			4476 => "11111110100110100100011000100001",
			4477 => "11111101011101010100011000100001",
			4478 => "00000000101001110100011000100001",
			4479 => "0000001000000000001001101000000100",
			4480 => "00000001101011010100011000100001",
			4481 => "0000001100000000000111111000001000",
			4482 => "0000001100000000001010000000000100",
			4483 => "11111111111011010100011000100001",
			4484 => "11111111000111010100011000100001",
			4485 => "0000001100000000000111111000000100",
			4486 => "00000000100111000100011000100001",
			4487 => "11111111111111110100011000100001",
			4488 => "0000000111000000000100010110010000",
			4489 => "0000000011000000000000101000111000",
			4490 => "0000001000000000001100000100010000",
			4491 => "0000000010000000000010110100001000",
			4492 => "0000001100000000000111111000000100",
			4493 => "11111110000000010100100010101101",
			4494 => "00000001011111010100100010101101",
			4495 => "0000001110000000001101010000000100",
			4496 => "00000000000000000100100010101101",
			4497 => "11111011011010110100100010101101",
			4498 => "0000000100000000000000010100010000",
			4499 => "0000000110000000001101111100001100",
			4500 => "0000001100000000000000110000000100",
			4501 => "00000000101001110100100010101101",
			4502 => "0000000001000000000110000000000100",
			4503 => "00000000111001100100100010101101",
			4504 => "00000001110101100100100010101101",
			4505 => "00000000011001100100100010101101",
			4506 => "0000000000000000001110111100001000",
			4507 => "0000000011000000001110111100000100",
			4508 => "00000000000000000100100010101101",
			4509 => "11111100110110010100100010101101",
			4510 => "0000001001000000000010001100001000",
			4511 => "0000000010000000001101000100000100",
			4512 => "00000001001110100100100010101101",
			4513 => "11111111100110100100100010101101",
			4514 => "0000001110000000001101010000000100",
			4515 => "11111111001001110100100010101101",
			4516 => "00000001101000100100100010101101",
			4517 => "0000001100000000000111111000101000",
			4518 => "0000001100000000000000110000010000",
			4519 => "0000000100000000000011010100001100",
			4520 => "0000000011000000001101100000001000",
			4521 => "0000000111000000000111111000000100",
			4522 => "00000000110011110100100010101101",
			4523 => "00000010100101010100100010101101",
			4524 => "11111110010111100100100010101101",
			4525 => "11111101101010100100100010101101",
			4526 => "0000000010000000001110101000001000",
			4527 => "0000001000000000001001101000000100",
			4528 => "11111111001001010100100010101101",
			4529 => "11111100010111110100100010101101",
			4530 => "0000001010000000000110011000001000",
			4531 => "0000000000000000000010111100000100",
			4532 => "11111101111011000100100010101101",
			4533 => "00000000000101110100100010101101",
			4534 => "0000001000000000000111000100000100",
			4535 => "11111101101010100100100010101101",
			4536 => "11111111001010010100100010101101",
			4537 => "0000000111000000000111111000011000",
			4538 => "0000000011000000001100001000001000",
			4539 => "0000000010000000001001010000000100",
			4540 => "00000001110111110100100010101101",
			4541 => "11111111110110010100100010101101",
			4542 => "0000001111000000000111110000001000",
			4543 => "0000001100000000000100010100000100",
			4544 => "11111100101111100100100010101101",
			4545 => "11111110111111110100100010101101",
			4546 => "0000000010000000001100010100000100",
			4547 => "00000010010000110100100010101101",
			4548 => "11111111101000100100100010101101",
			4549 => "0000001110000000001110111100001100",
			4550 => "0000001111000000000000011100000100",
			4551 => "00000000001001010100100010101101",
			4552 => "0000000011000000000100000000000100",
			4553 => "00000001001111000100100010101101",
			4554 => "00000010011001010100100010101101",
			4555 => "0000000111000000000111111000000100",
			4556 => "00000001011111000100100010101101",
			4557 => "0000001101000000001110001100000100",
			4558 => "11111111000000000100100010101101",
			4559 => "00000000110111010100100010101101",
			4560 => "0000000111000000000000101001001100",
			4561 => "0000000111000000000000101000111000",
			4562 => "0000001111000000000001101000011100",
			4563 => "0000001010000000001000100100001100",
			4564 => "0000000110000000001011111100000100",
			4565 => "11111110000101000100100010101101",
			4566 => "0000001100000000000100010100000100",
			4567 => "00000001111011010100100010101101",
			4568 => "00000000000000000100100010101101",
			4569 => "0000001110000000000010011000001000",
			4570 => "0000001101000000001100110000000100",
			4571 => "11111111010110100100100010101101",
			4572 => "00000001001100110100100010101101",
			4573 => "0000001111000000000110100100000100",
			4574 => "11111011111001010100100010101101",
			4575 => "11111110100111100100100010101101",
			4576 => "0000001100000000000000101000010000",
			4577 => "0000000111000000001011000100001000",
			4578 => "0000000111000000000100010100000100",
			4579 => "00000000011010110100100010101101",
			4580 => "11111111101010000100100010101101",
			4581 => "0000001010000000000110011100000100",
			4582 => "00000000101001000100100010101101",
			4583 => "11111110100110110100100010101101",
			4584 => "0000000001000000001100110100000100",
			4585 => "00000000000000010100100010101101",
			4586 => "0000001001000000000111100100000100",
			4587 => "11111101010100110100100010101101",
			4588 => "11111111000001010100100010101101",
			4589 => "0000001001000000000111100100010000",
			4590 => "0000001101000000001100101100001000",
			4591 => "0000001100000000000100010100000100",
			4592 => "00000010001011000100100010101101",
			4593 => "00000000010100000100100010101101",
			4594 => "0000000011000000001100110000000100",
			4595 => "11111111101100010100100010101101",
			4596 => "00000001001000100100100010101101",
			4597 => "00000010110100100100100010101101",
			4598 => "0000000111000000001100001000110000",
			4599 => "0000001010000000001100011100011100",
			4600 => "0000000000000000001110111100010000",
			4601 => "0000001001000000000110101000001000",
			4602 => "0000000001000000001110100000000100",
			4603 => "11111111100110000100100010101101",
			4604 => "11111101000101010100100010101101",
			4605 => "0000001010000000000001010000000100",
			4606 => "11111111101111000100100010101101",
			4607 => "11111110100101000100100010101101",
			4608 => "0000001101000000001101111000001000",
			4609 => "0000001101000000000110000100000100",
			4610 => "11111111100000100100100010101101",
			4611 => "00000001100001000100100010101101",
			4612 => "11111111001001100100100010101101",
			4613 => "0000001010000000000110011100001000",
			4614 => "0000001000000000000010101000000100",
			4615 => "11111100000010000100100010101101",
			4616 => "11111110100101100100100010101101",
			4617 => "0000001100000000000100010100001000",
			4618 => "0000001100000000000100010100000100",
			4619 => "00000000001001000100100010101101",
			4620 => "11111101100000100100100010101101",
			4621 => "00000000110010010100100010101101",
			4622 => "0000000111000000001100001000100000",
			4623 => "0000000111000000001100001000010000",
			4624 => "0000000010000000001100010100001000",
			4625 => "0000000111000000001100001000000100",
			4626 => "00000000110100000100100010101101",
			4627 => "11111111100011110100100010101101",
			4628 => "0000000110000000001010011000000100",
			4629 => "00000010000001100100100010101101",
			4630 => "00000000001111110100100010101101",
			4631 => "0000000100000000001100001100001000",
			4632 => "0000001000000000001001101000000100",
			4633 => "00000001100000100100100010101101",
			4634 => "00000100000011110100100010101101",
			4635 => "0000000000000000000011010000000100",
			4636 => "11111111111000100100100010101101",
			4637 => "00000001000101010100100010101101",
			4638 => "0000000111000000000100000000001100",
			4639 => "0000000100000000000010100100001000",
			4640 => "0000001010000000000110011100000100",
			4641 => "11111111001010110100100010101101",
			4642 => "11111100011001100100100010101101",
			4643 => "00000001100000010100100010101101",
			4644 => "0000001001000000001101101000001000",
			4645 => "0000001110000000001100101100000100",
			4646 => "11111111111110000100100010101101",
			4647 => "11111111000000110100100010101101",
			4648 => "0000000111000000000100000000000100",
			4649 => "00000001000011000100100010101101",
			4650 => "00000000000101010100100010101101",
			4651 => "0000000100000000000110111100000100",
			4652 => "11111110001100010100101000010001",
			4653 => "0000000111000000000000101001011000",
			4654 => "0000000111000000000100010100110000",
			4655 => "0000000111000000000100010100010000",
			4656 => "0000000001000000001100110100001100",
			4657 => "0000001001000000000111100100001000",
			4658 => "0000000101000000001100101100000100",
			4659 => "11111111111001000100101000010001",
			4660 => "00000010101010100100101000010001",
			4661 => "00000010011001110100101000010001",
			4662 => "11111110001010010100101000010001",
			4663 => "0000001011000000000100010100010000",
			4664 => "0000001111000000001010111000001000",
			4665 => "0000001100000000000111111000000100",
			4666 => "00000000000000000100101000010001",
			4667 => "11111100111001100100101000010001",
			4668 => "0000001011000000000100010100000100",
			4669 => "00000000101000000100101000010001",
			4670 => "00000001110111110100101000010001",
			4671 => "0000001011000000001011000100001000",
			4672 => "0000001100000000000111111000000100",
			4673 => "11111101011100100100101000010001",
			4674 => "11111111100011100100101000010001",
			4675 => "0000001111000000001011110100000100",
			4676 => "00000000001101110100101000010001",
			4677 => "00000001101010010100101000010001",
			4678 => "0000000101000000000011011100010100",
			4679 => "0000000100000000001001001100001000",
			4680 => "0000000111000000001011000100000100",
			4681 => "11111110100001000100101000010001",
			4682 => "00000001101011010100101000010001",
			4683 => "0000000010000000000010011100001000",
			4684 => "0000000011000000001011000100000100",
			4685 => "11111110010001110100101000010001",
			4686 => "11111011111011010100101000010001",
			4687 => "00000000010001010100101000010001",
			4688 => "0000000010000000000010000100010000",
			4689 => "0000000100000000001111100000001000",
			4690 => "0000000001000000000010001100000100",
			4691 => "11111111101000110100101000010001",
			4692 => "00000001001101100100101000010001",
			4693 => "0000001101000000000110000100000100",
			4694 => "11111111111111000100101000010001",
			4695 => "00000001001101100100101000010001",
			4696 => "11111101000110000100101000010001",
			4697 => "0000000111000000000000101000011000",
			4698 => "0000000110000000000111101000000100",
			4699 => "11111110100001000100101000010001",
			4700 => "0000000101000000001110001100010000",
			4701 => "0000000101000000000110000100001000",
			4702 => "0000001100000000000100010100000100",
			4703 => "00000001010000110100101000010001",
			4704 => "11111111010010010100101000010001",
			4705 => "0000000110000000001101111100000100",
			4706 => "00000000110001000100101000010001",
			4707 => "00000010011000100100101000010001",
			4708 => "00000000000101110100101000010001",
			4709 => "0000001010000000000111110100100000",
			4710 => "0000001100000000000100000000010000",
			4711 => "0000000011000000001010111100001000",
			4712 => "0000000011000000000000001100000100",
			4713 => "00000001000011000100101000010001",
			4714 => "11111110101110000100101000010001",
			4715 => "0000000110000000001101111100000100",
			4716 => "00000001111001000100101000010001",
			4717 => "00000000000000000100101000010001",
			4718 => "0000000100000000001111101000001000",
			4719 => "0000000100000000001011101100000100",
			4720 => "11111111010001010100101000010001",
			4721 => "11111110001100010100101000010001",
			4722 => "0000000010000000000111011000000100",
			4723 => "00000001100101010100101000010001",
			4724 => "11111111101010110100101000010001",
			4725 => "0000000100000000000100001100010000",
			4726 => "0000001100000000000111111000001000",
			4727 => "0000000100000000001000001000000100",
			4728 => "00000000010111110100101000010001",
			4729 => "00000010010010000100101000010001",
			4730 => "0000001001000000001011101000000100",
			4731 => "11111111110110000100101000010001",
			4732 => "00000000000110010100101000010001",
			4733 => "0000001000000000001111001000001000",
			4734 => "0000000100000000001111100000000100",
			4735 => "11111011111000010100101000010001",
			4736 => "11111111000110000100101000010001",
			4737 => "0000001000000000000010101000000100",
			4738 => "00000000110111100100101000010001",
			4739 => "11111111111100000100101000010001",
			4740 => "0000001001000000000110101010110000",
			4741 => "0000000011000000000011011101001100",
			4742 => "0000001111000000000110110100100100",
			4743 => "0000000011000000001001110000100000",
			4744 => "0000001110000000000011010000010000",
			4745 => "0000001100000000000100010100001000",
			4746 => "0000001100000000001010000000000100",
			4747 => "00000000100101100100110010100101",
			4748 => "11111111110110000100110010100101",
			4749 => "0000000011000000000100010100000100",
			4750 => "00000000010001010100110010100101",
			4751 => "00000001011111000100110010100101",
			4752 => "0000000110000000001101111100001000",
			4753 => "0000001001000000001001111000000100",
			4754 => "11111111011110100100110010100101",
			4755 => "00000000001111110100110010100101",
			4756 => "0000000110000000000100110100000100",
			4757 => "11111110100101110100110010100101",
			4758 => "11111111110001010100110010100101",
			4759 => "00000001010010110100110010100101",
			4760 => "0000001001000000001001111000011000",
			4761 => "0000000111000000000100010100001100",
			4762 => "0000000101000000001101100000001000",
			4763 => "0000000011000000001001110000000100",
			4764 => "00000000100010000100110010100101",
			4765 => "11111111000101100100110010100101",
			4766 => "11111110100000010100110010100101",
			4767 => "0000001000000000000110001000000100",
			4768 => "11111111011100000100110010100101",
			4769 => "0000000000000000001000011000000100",
			4770 => "00000001110111000100110010100101",
			4771 => "00000000000000000100110010100101",
			4772 => "0000000100000000001010110100000100",
			4773 => "11111111110011100100110010100101",
			4774 => "0000001001000000000110101000001000",
			4775 => "0000000111000000001100001000000100",
			4776 => "00000001111111010100110010100101",
			4777 => "00000000100110000100110010100101",
			4778 => "00000000011111010100110010100101",
			4779 => "0000000010000000000101110000101000",
			4780 => "0000000101000000000101101100010000",
			4781 => "0000001101000000001100110000000100",
			4782 => "00000000101001000100110010100101",
			4783 => "0000000010000000001101000100000100",
			4784 => "00000010000101100100110010100101",
			4785 => "0000001001000000001001111000000100",
			4786 => "00000000001011000100110010100101",
			4787 => "11111101111100010100110010100101",
			4788 => "0000000101000000000101101100001000",
			4789 => "0000001111000000001011011100000100",
			4790 => "00000001101110100100110010100101",
			4791 => "00000000011000000100110010100101",
			4792 => "0000000000000000000000111000001000",
			4793 => "0000000100000000000101000000000100",
			4794 => "11111110001000110100110010100101",
			4795 => "00000000001111010100110010100101",
			4796 => "0000001100000000000100010100000100",
			4797 => "11111111100100010100110010100101",
			4798 => "11111101110110010100110010100101",
			4799 => "0000000100000000001001001100011100",
			4800 => "0000000011000000000101101100001100",
			4801 => "0000000101000000000101101100001000",
			4802 => "0000000000000000001010000000000100",
			4803 => "00000000000110000100110010100101",
			4804 => "00000010000101000100110010100101",
			4805 => "00000010011100010100110010100101",
			4806 => "0000001111000000000001001000001000",
			4807 => "0000000100000000001101001000000100",
			4808 => "11111111011110100100110010100101",
			4809 => "11111101110001100100110010100101",
			4810 => "0000001110000000000101101100000100",
			4811 => "00000001111100100100110010100101",
			4812 => "00000000000000000100110010100101",
			4813 => "0000001100000000000100010100010000",
			4814 => "0000001101000000000110000100001000",
			4815 => "0000000101000000001100110000000100",
			4816 => "00000000001001100100110010100101",
			4817 => "11111110100110010100110010100101",
			4818 => "0000001011000000001100001000000100",
			4819 => "00000010000001100100110010100101",
			4820 => "00000000000000000100110010100101",
			4821 => "0000001011000000000000101000001000",
			4822 => "0000000111000000000100010100000100",
			4823 => "11111110111011110100110010100101",
			4824 => "00000001000001100100110010100101",
			4825 => "0000000110000000001101111100000100",
			4826 => "00000001000110100100110010100101",
			4827 => "11111110001000010100110010100101",
			4828 => "0000000011000000000101101101100000",
			4829 => "0000001011000000001100001000100100",
			4830 => "0000000110000000000001111000010000",
			4831 => "0000000100000000001011110000000100",
			4832 => "11111110111100000100110010100101",
			4833 => "0000000011000000001100110000001000",
			4834 => "0000001111000000000000011100000100",
			4835 => "00000001111001000100110010100101",
			4836 => "11111111110011110100110010100101",
			4837 => "00000010001111110100110010100101",
			4838 => "0000001000000000001001101000000100",
			4839 => "11111101111101000100110010100101",
			4840 => "0000000000000000001010000000001000",
			4841 => "0000000000000000000000110000000100",
			4842 => "00000000000011000100110010100101",
			4843 => "11111101011110110100110010100101",
			4844 => "0000001100000000000000101000000100",
			4845 => "00000000111010100100110010100101",
			4846 => "11111111010110000100110010100101",
			4847 => "0000001111000000001011011100100000",
			4848 => "0000000011000000001101100000010000",
			4849 => "0000001110000000000000111000001000",
			4850 => "0000000110000000001100011000000100",
			4851 => "00000000110011100100110010100101",
			4852 => "11111110110010100100110010100101",
			4853 => "0000001110000000000111111000000100",
			4854 => "00000001110101110100110010100101",
			4855 => "00000000100101110100110010100101",
			4856 => "0000001001000000000111100100001000",
			4857 => "0000001100000000000100010100000100",
			4858 => "11111101110100110100110010100101",
			4859 => "11111111101001110100110010100101",
			4860 => "0000000100000000001010110100000100",
			4861 => "00000000001101110100110010100101",
			4862 => "00000001110110010100110010100101",
			4863 => "0000001111000000000010001000001100",
			4864 => "0000001011000000001100001000000100",
			4865 => "00000001011110110100110010100101",
			4866 => "0000001110000000001011000100000100",
			4867 => "00000001101000100100110010100101",
			4868 => "00000011001010010100110010100101",
			4869 => "0000001111000000000101110100001000",
			4870 => "0000001111000000000100010000000100",
			4871 => "00000000110101110100110010100101",
			4872 => "11111110101011110100110010100101",
			4873 => "0000000110000000001010011000000100",
			4874 => "00000010000001010100110010100101",
			4875 => "00000000110101110100110010100101",
			4876 => "0000000011000000000110000100010000",
			4877 => "0000000010000000000100101000001000",
			4878 => "0000001101000000001110001100000100",
			4879 => "00000001110100110100110010100101",
			4880 => "11111110110001110100110010100101",
			4881 => "0000001000000000000111000100000100",
			4882 => "11111101001001000100110010100101",
			4883 => "11111111100101110100110010100101",
			4884 => "0000000011000000000110000100001100",
			4885 => "0000001000000000000111000100001000",
			4886 => "0000000101000000001100101100000100",
			4887 => "00000001000000110100110010100101",
			4888 => "00000010011100000100110010100101",
			4889 => "00000000000000000100110010100101",
			4890 => "0000000010000000000101110000010000",
			4891 => "0000001000000000000110001000001000",
			4892 => "0000001110000000001011000100000100",
			4893 => "00000010000010000100110010100101",
			4894 => "11111111110101100100110010100101",
			4895 => "0000000011000000001110001100000100",
			4896 => "11111101110011110100110010100101",
			4897 => "11111111111100010100110010100101",
			4898 => "0000000111000000001100001000001000",
			4899 => "0000000011000000000000001100000100",
			4900 => "00000000110011000100110010100101",
			4901 => "00000000000010000100110010100101",
			4902 => "0000001011000000001100001000000100",
			4903 => "11111110101111010100110010100101",
			4904 => "00000000000010100100110010100101",
			4905 => "0000001001000000000010001110010100",
			4906 => "0000001110000000001111000101011100",
			4907 => "0000001010000000000101000100101100",
			4908 => "0000001000000000000111000100010100",
			4909 => "0000000001000000000110000000010000",
			4910 => "0000001100000000001010000000001000",
			4911 => "0000000110000000000001111000000100",
			4912 => "11111101001001000100111101011001",
			4913 => "11111111101001010100111101011001",
			4914 => "0000000111000000000111111000000100",
			4915 => "11111110110110000100111101011001",
			4916 => "00000001101101010100111101011001",
			4917 => "11111101011000000100111101011001",
			4918 => "0000001001000000001110100000001100",
			4919 => "0000001110000000001011010100001000",
			4920 => "0000000010000000001111010000000100",
			4921 => "00000001110101110100111101011001",
			4922 => "00000000000000000100111101011001",
			4923 => "11111101111010110100111101011001",
			4924 => "0000000010000000001111010000001000",
			4925 => "0000000001000000000000011000000100",
			4926 => "00000000100110100100111101011001",
			4927 => "00000001101101010100111101011001",
			4928 => "00000000001101110100111101011001",
			4929 => "0000000101000000000011011100011100",
			4930 => "0000000111000000000111111000001100",
			4931 => "0000000010000000001010010100000100",
			4932 => "00000001011100010100111101011001",
			4933 => "0000001111000000001010001100000100",
			4934 => "11111101110010000100111101011001",
			4935 => "00000000110110000100111101011001",
			4936 => "0000000110000000001101111100001000",
			4937 => "0000000110000000000001111000000100",
			4938 => "11111110110001100100111101011001",
			4939 => "11111100000101110100111101011001",
			4940 => "0000001100000000000111111000000100",
			4941 => "00000001011011000100111101011001",
			4942 => "00000000000000000100111101011001",
			4943 => "0000001101000000001101100000001000",
			4944 => "0000001101000000000011011100000100",
			4945 => "11111110010001100100111101011001",
			4946 => "11111011001111000100111101011001",
			4947 => "0000001100000000000100010100000100",
			4948 => "00000001010010010100111101011001",
			4949 => "0000000010000000001110101000000100",
			4950 => "00000000011111010100111101011001",
			4951 => "11111110000101010100111101011001",
			4952 => "0000001000000000001111001000100000",
			4953 => "0000001000000000001011010100010000",
			4954 => "0000000111000000000100010100001100",
			4955 => "0000001010000000001000100100000100",
			4956 => "11111111011000000100111101011001",
			4957 => "0000000101000000001000111000000100",
			4958 => "00000000000000000100111101011001",
			4959 => "11111100010011010100111101011001",
			4960 => "00000001000001100100111101011001",
			4961 => "0000000001000000000000011000000100",
			4962 => "11111101010110110100111101011001",
			4963 => "0000001011000000000111111000000100",
			4964 => "11111111111011100100111101011001",
			4965 => "0000001111000000000111010000000100",
			4966 => "00000000100001110100111101011001",
			4967 => "00000001111110110100111101011001",
			4968 => "0000001110000000000010011000000100",
			4969 => "11111101001000110100111101011001",
			4970 => "0000001001000000000010001100010000",
			4971 => "0000001000000000000010101000001000",
			4972 => "0000001010000000001010110000000100",
			4973 => "00000000001100100100111101011001",
			4974 => "11111101100001000100111101011001",
			4975 => "0000000100000000000001101100000100",
			4976 => "00000000010001110100111101011001",
			4977 => "11111101101111000100111101011001",
			4978 => "00000000001101000100111101011001",
			4979 => "0000001100000000000111111001101000",
			4980 => "0000000111000000001011000100111100",
			4981 => "0000000110000000000001111000011100",
			4982 => "0000000101000000000011011100001100",
			4983 => "0000001100000000000111111000001000",
			4984 => "0000001000000000000110001000000100",
			4985 => "11111110111011010100111101011001",
			4986 => "00000001101011110100111101011001",
			4987 => "11111011111110110100111101011001",
			4988 => "0000001110000000000100010100001000",
			4989 => "0000000101000000000101101100000100",
			4990 => "00000000111001100100111101011001",
			4991 => "11111110111111000100111101011001",
			4992 => "0000000110000000000001111000000100",
			4993 => "11111111111110000100111101011001",
			4994 => "11111110010110110100111101011001",
			4995 => "0000001100000000000111111000010000",
			4996 => "0000001010000000001001000100001000",
			4997 => "0000000001000000001110100000000100",
			4998 => "00000010110101010100111101011001",
			4999 => "00000000000000000100111101011001",
			5000 => "0000001100000000001010000000000100",
			5001 => "00000000000100100100111101011001",
			5002 => "11111110101111000100111101011001",
			5003 => "0000000110000000001101111100001000",
			5004 => "0000000111000000000100010100000100",
			5005 => "00000010011110110100111101011001",
			5006 => "00000000101000110100111101011001",
			5007 => "0000000110000000001101111100000100",
			5008 => "11111111010110100100111101011001",
			5009 => "00000000101010110100111101011001",
			5010 => "0000000111000000001100001000100000",
			5011 => "0000000110000000001100011000010000",
			5012 => "0000001100000000000111111000001000",
			5013 => "0000000001000000001110100000000100",
			5014 => "00000001000011010100111101011001",
			5015 => "00000010100011000100111101011001",
			5016 => "0000001100000000000111111000000100",
			5017 => "11111111111100010100111101011001",
			5018 => "00000001010000100100111101011001",
			5019 => "0000001010000000001010110000001000",
			5020 => "0000000101000000001100101100000100",
			5021 => "11111101010001110100111101011001",
			5022 => "11111111100111000100111101011001",
			5023 => "0000000010000000000010011100000100",
			5024 => "11111110001001000100111101011001",
			5025 => "00000001010111110100111101011001",
			5026 => "0000001010000000001001000100000100",
			5027 => "00000000001011010100111101011001",
			5028 => "0000000100000000000011001100000100",
			5029 => "11111101010100010100111101011001",
			5030 => "11111111011111010100111101011001",
			5031 => "0000001100000000000100010100101100",
			5032 => "0000000101000000001110001100011100",
			5033 => "0000001001000000000110101000010000",
			5034 => "0000000101000000000110000100001000",
			5035 => "0000000101000000001101100000000100",
			5036 => "00000000000010110100111101011001",
			5037 => "11111110110100100100111101011001",
			5038 => "0000000010000000000010011100000100",
			5039 => "00000010111100010100111101011001",
			5040 => "00000000000000000100111101011001",
			5041 => "0000000100000000001000011100000100",
			5042 => "00000000110001100100111101011001",
			5043 => "0000001011000000000000101000000100",
			5044 => "11111111001001010100111101011001",
			5045 => "11111101011101100100111101011001",
			5046 => "0000001011000000001000111100001000",
			5047 => "0000001011000000000100000000000100",
			5048 => "11111111010010010100111101011001",
			5049 => "00000011101011000100111101011001",
			5050 => "0000001000000000001011010100000100",
			5051 => "11111111010001010100111101011001",
			5052 => "11111110001010010100111101011001",
			5053 => "0000001100000000000100010100010100",
			5054 => "0000001101000000000101101100000100",
			5055 => "00000010000110010100111101011001",
			5056 => "0000001011000000000000101000001000",
			5057 => "0000001011000000000000101000000100",
			5058 => "00000000011111010100111101011001",
			5059 => "11111101101000010100111101011001",
			5060 => "0000000001000000001100110100000100",
			5061 => "00000010000011000100111101011001",
			5062 => "00000000001000000100111101011001",
			5063 => "0000001001000000000110101000010000",
			5064 => "0000001110000000000000101000001000",
			5065 => "0000001001000000000110101000000100",
			5066 => "11111111110100000100111101011001",
			5067 => "00000000100011110100111101011001",
			5068 => "0000001011000000001011000100000100",
			5069 => "00000001101001010100111101011001",
			5070 => "11111111000111100100111101011001",
			5071 => "0000001110000000001011000100001000",
			5072 => "0000000111000000001100001000000100",
			5073 => "00000010001111100100111101011001",
			5074 => "00000000101011010100111101011001",
			5075 => "0000001100000000000100010100000100",
			5076 => "00000001000110010100111101011001",
			5077 => "00000000000010110100111101011001",
			5078 => "0000001110000000001100001010111100",
			5079 => "0000001111000000000010001001101000",
			5080 => "0000000100000000000000010100111000",
			5081 => "0000000011000000000100010100011000",
			5082 => "0000001000000000001100000100001000",
			5083 => "0000001011000000000100010100000100",
			5084 => "11111101111100000101001000111101",
			5085 => "00000001010110100101001000111101",
			5086 => "0000001000000000000111000100001000",
			5087 => "0000000111000000000100010100000100",
			5088 => "00000001100001100101001000111101",
			5089 => "00000000011010010101001000111101",
			5090 => "0000001011000000000100010100000100",
			5091 => "00000001000101000101001000111101",
			5092 => "11111101110101000101001000111101",
			5093 => "0000001101000000001110001100010000",
			5094 => "0000000011000000001101100000001000",
			5095 => "0000000010000000001110101000000100",
			5096 => "11111111101111100101001000111101",
			5097 => "00000000010000100101001000111101",
			5098 => "0000001001000000000110101000000100",
			5099 => "11111101111000000101001000111101",
			5100 => "11111111110010000101001000111101",
			5101 => "0000000110000000000100110100001000",
			5102 => "0000000100000000000001011100000100",
			5103 => "11111110010010000101001000111101",
			5104 => "00000001011010110101001000111101",
			5105 => "0000000111000000001100001000000100",
			5106 => "11111110001101010101001000111101",
			5107 => "00000000010101110101001000111101",
			5108 => "0000000000000000001011000100011100",
			5109 => "0000001101000000001110001100010000",
			5110 => "0000001001000000000110101000001000",
			5111 => "0000000011000000001000111000000100",
			5112 => "11111111100100100101001000111101",
			5113 => "11111110000001110101001000111101",
			5114 => "0000001100000000000100010100000100",
			5115 => "11111111110100110101001000111101",
			5116 => "00000001100010100101001000111101",
			5117 => "0000000000000000000111111000000100",
			5118 => "00000000011000110101001000111101",
			5119 => "0000001110000000000111111000000100",
			5120 => "11111100101100010101001000111101",
			5121 => "11111111000110000101001000111101",
			5122 => "0000000100000000000010100100001000",
			5123 => "0000001111000000001011011100000100",
			5124 => "00000001110001000101001000111101",
			5125 => "00000000100000100101001000111101",
			5126 => "0000001110000000001110111100001000",
			5127 => "0000000111000000000111111000000100",
			5128 => "11111110100100000101001000111101",
			5129 => "00000000001010100101001000111101",
			5130 => "11111101110111010101001000111101",
			5131 => "0000001110000000000000101000111000",
			5132 => "0000001110000000001011000100100000",
			5133 => "0000000111000000001011000100010000",
			5134 => "0000000001000000001110100000001000",
			5135 => "0000001001000000000010001100000100",
			5136 => "11111111011001100101001000111101",
			5137 => "00000000101101100101001000111101",
			5138 => "0000000011000000000011011100000100",
			5139 => "00000001010110000101001000111101",
			5140 => "11111110101101000101001000111101",
			5141 => "0000001011000000000100000000001000",
			5142 => "0000001110000000001011000100000100",
			5143 => "00000001011110100101001000111101",
			5144 => "00000000000011000101001000111101",
			5145 => "0000000110000000001100011000000100",
			5146 => "00000001000110000101001000111101",
			5147 => "11111101101111000101001000111101",
			5148 => "0000000110000000000100110100001100",
			5149 => "0000001000000000001011010100000100",
			5150 => "11111110101110100101001000111101",
			5151 => "0000000011000000000101101100000100",
			5152 => "00000000101111010101001000111101",
			5153 => "00000010010101010101001000111101",
			5154 => "0000001011000000001000111100001000",
			5155 => "0000000100000000001111100000000100",
			5156 => "11111101111001010101001000111101",
			5157 => "00000000010000000101001000111101",
			5158 => "00000000101010000101001000111101",
			5159 => "0000000001000000001110100000000100",
			5160 => "11111101111010010101001000111101",
			5161 => "0000000011000000000101101100001100",
			5162 => "0000001011000000001100001000001000",
			5163 => "0000000000000000000100010100000100",
			5164 => "00000010010011100101001000111101",
			5165 => "00000000110111000101001000111101",
			5166 => "00000000000000000101001000111101",
			5167 => "0000001101000000001100101100000100",
			5168 => "11111110111010100101001000111101",
			5169 => "0000001111000000000100010000000100",
			5170 => "11111111101000110101001000111101",
			5171 => "00000001100100010101001000111101",
			5172 => "0000001001000000000111100101011000",
			5173 => "0000001111000000001011110100100000",
			5174 => "0000000010000000000111111100011100",
			5175 => "0000001111000000000110110100001100",
			5176 => "0000001001000000000110101000001000",
			5177 => "0000000000000000000001010100000100",
			5178 => "00000000000000000101001000111101",
			5179 => "00000000101100100101001000111101",
			5180 => "11111110000011000101001000111101",
			5181 => "0000001000000000001001101000001000",
			5182 => "0000001111000000000010001000000100",
			5183 => "11111110111111000101001000111101",
			5184 => "00000001001101110101001000111101",
			5185 => "0000000011000000000101101100000100",
			5186 => "00000000001001000101001000111101",
			5187 => "11111110110010000101001000111101",
			5188 => "11111101001111110101001000111101",
			5189 => "0000000110000000001100011000011100",
			5190 => "0000000110000000000001111000001100",
			5191 => "0000000000000000000011111100001000",
			5192 => "0000000011000000001101111000000100",
			5193 => "00000000100011100101001000111101",
			5194 => "11111110010111010101001000111101",
			5195 => "11111010001110110101001000111101",
			5196 => "0000001000000000001011010100001000",
			5197 => "0000000011000000000000001100000100",
			5198 => "00000001011100100101001000111101",
			5199 => "11111110110000100101001000111101",
			5200 => "0000000100000000001101001000000100",
			5201 => "11111111000110010101001000111101",
			5202 => "00000000001100110101001000111101",
			5203 => "0000000000000000000100010100001100",
			5204 => "0000000011000000001100101100000100",
			5205 => "00000000001001010101001000111101",
			5206 => "0000000100000000000000010100000100",
			5207 => "11111110101000000101001000111101",
			5208 => "11111101000100110101001000111101",
			5209 => "0000001001000000000110101000001000",
			5210 => "0000001011000000000000101000000100",
			5211 => "00000001110000100101001000111101",
			5212 => "11111101111001010101001000111101",
			5213 => "0000001100000000000000101000000100",
			5214 => "00000001100110100101001000111101",
			5215 => "00000000001101010101001000111101",
			5216 => "0000000011000000001110001100101100",
			5217 => "0000001001000000001101101000011100",
			5218 => "0000001011000000001100001000001100",
			5219 => "0000000110000000001101111100000100",
			5220 => "00000010110100010101001000111101",
			5221 => "0000001111000000000101110100000100",
			5222 => "11111111010100110101001000111101",
			5223 => "00000010010000000101001000111101",
			5224 => "0000000001000000001100110100001000",
			5225 => "0000001011000000000100000000000100",
			5226 => "11111111111111100101001000111101",
			5227 => "00000001111111110101001000111101",
			5228 => "0000000110000000000100110100000100",
			5229 => "11111110001010100101001000111101",
			5230 => "00000000100000100101001000111101",
			5231 => "0000001101000000001101111000000100",
			5232 => "00000011101011100101001000111101",
			5233 => "0000001110000000001000111000001000",
			5234 => "0000000000000000001111000100000100",
			5235 => "00000000100100100101001000111101",
			5236 => "00000010000110100101001000111101",
			5237 => "00000000000000000101001000111101",
			5238 => "0000000001000000001100110100011000",
			5239 => "0000000100000000001010110100001100",
			5240 => "0000001101000000000000001100001000",
			5241 => "0000001111000000001010010100000100",
			5242 => "11111111010011000101001000111101",
			5243 => "00000001010011110101001000111101",
			5244 => "11111110000110010101001000111101",
			5245 => "0000001111000000000010110100001000",
			5246 => "0000000111000000001100001000000100",
			5247 => "00000011000001010101001000111101",
			5248 => "00000001110101110101001000111101",
			5249 => "11111111000000010101001000111101",
			5250 => "0000001001000000000111100100001100",
			5251 => "0000000001000000001100110100000100",
			5252 => "11111101011001000101001000111101",
			5253 => "0000000010000000000010000100000100",
			5254 => "11111111011001010101001000111101",
			5255 => "00000010000100010101001000111101",
			5256 => "0000001011000000001100001000001000",
			5257 => "0000000111000000001100001000000100",
			5258 => "11111101101011100101001000111101",
			5259 => "11111111101001000101001000111101",
			5260 => "0000001011000000001000111100000100",
			5261 => "00000000011101110101001000111101",
			5262 => "11111111111110010101001000111101",
			5263 => "0000001111000000000000110111011000",
			5264 => "0000000011000000001001110001110100",
			5265 => "0000001001000000001001111000111100",
			5266 => "0000001011000000000000101000011100",
			5267 => "0000000011000000001000111000010000",
			5268 => "0000001011000000000100010100001000",
			5269 => "0000001111000000000110110100000100",
			5270 => "11111111110001010101010100011011",
			5271 => "00000000110101110101010100011011",
			5272 => "0000001111000000000000011100000100",
			5273 => "00000000001000110101010100011011",
			5274 => "00000001000111110101010100011011",
			5275 => "0000001100000000000000110000000100",
			5276 => "00000001111101110101010100011011",
			5277 => "0000000110000000001101111100000100",
			5278 => "11111110000010100101010100011011",
			5279 => "00000000001101000101010100011011",
			5280 => "0000001101000000000110000100010000",
			5281 => "0000001010000000001100011100001000",
			5282 => "0000001110000000001010000000000100",
			5283 => "00000000000000010101010100011011",
			5284 => "11111110010001100101010100011011",
			5285 => "0000001001000000001001111000000100",
			5286 => "00000000000000000101010100011011",
			5287 => "11111101000000100101010100011011",
			5288 => "0000001111000000000111010000001000",
			5289 => "0000001010000000001100000100000100",
			5290 => "00000001101001000101010100011011",
			5291 => "11111111000010010101010100011011",
			5292 => "0000000011000000001100001000000100",
			5293 => "00000000110100010101010100011011",
			5294 => "11111101110110010101010100011011",
			5295 => "0000001100000000000111111000011000",
			5296 => "0000000000000000000000111000001100",
			5297 => "0000000111000000000000101000001000",
			5298 => "0000001010000000001001000100000100",
			5299 => "00000000101010000101010100011011",
			5300 => "11111110011000100101010100011011",
			5301 => "00000010000110010101010100011011",
			5302 => "0000001101000000001100110000000100",
			5303 => "00000000000100110101010100011011",
			5304 => "0000001111000000000000011100000100",
			5305 => "00000001000101100101010100011011",
			5306 => "00000010000010100101010100011011",
			5307 => "0000001001000000001001111000010000",
			5308 => "0000000100000000001001001100001000",
			5309 => "0000000110000000000111101000000100",
			5310 => "00000000000000000101010100011011",
			5311 => "00000001111111010101010100011011",
			5312 => "0000000111000000000100010100000100",
			5313 => "11111110100110100101010100011011",
			5314 => "00000000111011000101010100011011",
			5315 => "0000000101000000000110000100001000",
			5316 => "0000000000000000001110111100000100",
			5317 => "11111111001011000101010100011011",
			5318 => "00000000100000100101010100011011",
			5319 => "0000000111000000001100001000000100",
			5320 => "00000001111001010101010100011011",
			5321 => "00000000000110010101010100011011",
			5322 => "0000000111000000000100010100101000",
			5323 => "0000001111000000000111110000011000",
			5324 => "0000001010000000001001000100001100",
			5325 => "0000000000000000000010111100001000",
			5326 => "0000001110000000001000111100000100",
			5327 => "11111110001111000101010100011011",
			5328 => "00000000000000000101010100011011",
			5329 => "00000001001111100101010100011011",
			5330 => "0000001110000000000100010100000100",
			5331 => "11111101100101000101010100011011",
			5332 => "0000000011000000001101100000000100",
			5333 => "11111111111010110101010100011011",
			5334 => "11111110001001010101010100011011",
			5335 => "0000000100000000001000001000000100",
			5336 => "00000010011000100101010100011011",
			5337 => "0000000011000000001101100000000100",
			5338 => "00000001100000000101010100011011",
			5339 => "0000001011000000001011000100000100",
			5340 => "11111111111100110101010100011011",
			5341 => "11111101100100010101010100011011",
			5342 => "0000001001000000000110101000100000",
			5343 => "0000001011000000001011000100010000",
			5344 => "0000001100000000000100010100001000",
			5345 => "0000001010000000000110011000000100",
			5346 => "00000001111011000101010100011011",
			5347 => "11111111101001100101010100011011",
			5348 => "0000000000000000000000110000000100",
			5349 => "00000000110111000101010100011011",
			5350 => "00000010010100100101010100011011",
			5351 => "0000000111000000001011000100001000",
			5352 => "0000001111000000000101110100000100",
			5353 => "11111110110110100101010100011011",
			5354 => "11111111110111000101010100011011",
			5355 => "0000001011000000000100000000000100",
			5356 => "11111111111110100101010100011011",
			5357 => "11111110011101110101010100011011",
			5358 => "0000000111000000000000101000001100",
			5359 => "0000001100000000000000101000001000",
			5360 => "0000000000000000000010011000000100",
			5361 => "11111111100100000101010100011011",
			5362 => "00000000101111010101010100011011",
			5363 => "11111110010111100101010100011011",
			5364 => "0000000111000000001100001000001000",
			5365 => "0000001110000000000011011100000100",
			5366 => "11111101001110000101010100011011",
			5367 => "00000000000000000101010100011011",
			5368 => "0000000111000000001000111000000100",
			5369 => "11111111110101000101010100011011",
			5370 => "00000000011000010101010100011011",
			5371 => "0000001110000000000100001001010100",
			5372 => "0000000000000000000000111000100100",
			5373 => "0000001100000000000100000000100000",
			5374 => "0000001110000000001101111000010000",
			5375 => "0000000101000000000000001100001000",
			5376 => "0000000110000000000100110100000100",
			5377 => "00000000000101110101010100011011",
			5378 => "00000011000001110101010100011011",
			5379 => "0000000111000000001100001000000100",
			5380 => "11111110010111000101010100011011",
			5381 => "00000000110110000101010100011011",
			5382 => "0000001010000000001001000100001000",
			5383 => "0000001101000000000001111100000100",
			5384 => "00000010010101000101010100011011",
			5385 => "11111111100100100101010100011011",
			5386 => "0000001111000000000110100000000100",
			5387 => "11111110010111010101010100011011",
			5388 => "00000000100111010101010100011011",
			5389 => "00000010101110110101010100011011",
			5390 => "0000000100000000001101001000010000",
			5391 => "0000001000000000000111000100001100",
			5392 => "0000000011000000000001111100001000",
			5393 => "0000001111000000001110101100000100",
			5394 => "11111110001011000101010100011011",
			5395 => "00000000110100100101010100011011",
			5396 => "11111101110100110101010100011011",
			5397 => "00000000000110010101010100011011",
			5398 => "0000001001000000001101101000010000",
			5399 => "0000001100000000000100000000001000",
			5400 => "0000001111000000001101000100000100",
			5401 => "00000000010110110101010100011011",
			5402 => "11111111001011100101010100011011",
			5403 => "0000000100000000000100001100000100",
			5404 => "11111101110001000101010100011011",
			5405 => "00000000101101100101010100011011",
			5406 => "0000000101000000001010111100001000",
			5407 => "0000001011000000000011011100000100",
			5408 => "00000000101010100101010100011011",
			5409 => "00000010000111100101010100011011",
			5410 => "0000000011000000001010111000000100",
			5411 => "11111100001010100101010100011011",
			5412 => "00000000010001110101010100011011",
			5413 => "0000001110000000000001111100100000",
			5414 => "0000001100000000000100000000010100",
			5415 => "0000000101000000001010111100010000",
			5416 => "0000000011000000001110110000001000",
			5417 => "0000000011000000000111001000000100",
			5418 => "11111111000011010101010100011011",
			5419 => "00000001100101100101010100011011",
			5420 => "0000001000000000000111000100000100",
			5421 => "11111111001110010101010100011011",
			5422 => "11111101111100100101010100011011",
			5423 => "00000001110011110101010100011011",
			5424 => "0000001001000000001111001100000100",
			5425 => "11111101100001100101010100011011",
			5426 => "0000001011000000000000001100000100",
			5427 => "00000000110010000101010100011011",
			5428 => "00000000000000000101010100011011",
			5429 => "0000000111000000000000101000000100",
			5430 => "11111110001111000101010100011011",
			5431 => "0000000101000000001100101000010000",
			5432 => "0000000100000000000011001100001000",
			5433 => "0000000100000000001000110100000100",
			5434 => "00000001101000000101010100011011",
			5435 => "11111110111110110101010100011011",
			5436 => "0000000011000000000100011000000100",
			5437 => "00000000000000000101010100011011",
			5438 => "00000010101010100101010100011011",
			5439 => "0000001101000000000111001000001000",
			5440 => "0000001111000000000101001000000100",
			5441 => "11111110101101100101010100011011",
			5442 => "00000001010001000101010100011011",
			5443 => "0000001011000000001101100000000100",
			5444 => "00000000100110010101010100011011",
			5445 => "11111111111110010101010100011011",
			5446 => "0000000111000000001110001101011000",
			5447 => "0000000100000000000110110000111100",
			5448 => "0000000011000000000010111100001000",
			5449 => "0000001101000000000100000000000100",
			5450 => "00000000110110110101011001001101",
			5451 => "00000010000111000101011001001101",
			5452 => "0000001001000000001100110100010100",
			5453 => "0000000011000000000000111000001000",
			5454 => "0000000111000000000111111000000100",
			5455 => "11111111100111010101011001001101",
			5456 => "00000001111101000101011001001101",
			5457 => "0000001111000000000110100100000100",
			5458 => "11111100100000110101011001001101",
			5459 => "0000000100000000001001001100000100",
			5460 => "00000000000001100101011001001101",
			5461 => "11111110000110000101011001001101",
			5462 => "0000000011000000000100010100010000",
			5463 => "0000001111000000000001101000001000",
			5464 => "0000000001000000000110000000000100",
			5465 => "00000000111110010101011001001101",
			5466 => "11111111100111110101011001001101",
			5467 => "0000001000000000001000101100000100",
			5468 => "00000001100011010101011001001101",
			5469 => "11111111101000110101011001001101",
			5470 => "0000001001000000000010001100001000",
			5471 => "0000000011000000001100001000000100",
			5472 => "11111111110110010101011001001101",
			5473 => "11111110011000000101011001001101",
			5474 => "0000000011000000001001110000000100",
			5475 => "00000000011101000101011001001101",
			5476 => "00000000001001000101011001001101",
			5477 => "0000000110000000001100011000001000",
			5478 => "0000001101000000000110000100000100",
			5479 => "11111110010101100101011001001101",
			5480 => "11111111111110010101011001001101",
			5481 => "0000000111000000000100010100000100",
			5482 => "00000001010001100101011001001101",
			5483 => "0000001110000000000000110000000100",
			5484 => "11111101010100010101011001001101",
			5485 => "0000000110000000001011001100001000",
			5486 => "0000001000000000001101010000000100",
			5487 => "11111111010101010101011001001101",
			5488 => "00000001000111100101011001001101",
			5489 => "11111110011001100101011001001101",
			5490 => "0000001000000000001001101000010000",
			5491 => "0000001001000000000100110100001100",
			5492 => "0000001001000000000001111000000100",
			5493 => "11111110011010110101011001001101",
			5494 => "0000001111000000000110100000000100",
			5495 => "11111110111011000101011001001101",
			5496 => "00000001110111000101011001001101",
			5497 => "11111110011001000101011001001101",
			5498 => "0000000100000000000011111000101000",
			5499 => "0000001010000000000001010100011000",
			5500 => "0000000100000000001011001000010000",
			5501 => "0000001110000000001100111000001000",
			5502 => "0000001011000000001010011100000100",
			5503 => "00000000000100010101011001001101",
			5504 => "00000001100010100101011001001101",
			5505 => "0000001011000000001110101100000100",
			5506 => "11111110011001110101011001001101",
			5507 => "00000000110111100101011001001101",
			5508 => "0000001010000000000101000100000100",
			5509 => "11111110001110110101011001001101",
			5510 => "11111111111000010101011001001101",
			5511 => "0000001111000000000000010100001000",
			5512 => "0000000000000000001011000100000100",
			5513 => "00000001001011000101011001001101",
			5514 => "00000010010001010101011001001101",
			5515 => "0000000111000000001001010100000100",
			5516 => "11111110011101010101011001001101",
			5517 => "00000010010111000101011001001101",
			5518 => "0000000100000000000000000000001000",
			5519 => "0000000000000000001010111100000100",
			5520 => "11111110100100110101011001001101",
			5521 => "00000001110001110101011001001101",
			5522 => "11111110011001110101011001001101",
			5523 => "0000000111000000001101111001100000",
			5524 => "0000000001000000000000011000100000",
			5525 => "0000000001000000001100100000000100",
			5526 => "11111110010101010101011110001001",
			5527 => "0000000011000000000000111000001100",
			5528 => "0000001011000000001110111100000100",
			5529 => "11111110110001100101011110001001",
			5530 => "0000000001000000001100100000000100",
			5531 => "00000000000011000101011110001001",
			5532 => "00000010001110110101011110001001",
			5533 => "0000001010000000001100011100001100",
			5534 => "0000001000000000000010101000001000",
			5535 => "0000000111000000000100010100000100",
			5536 => "11111110010010000101011110001001",
			5537 => "11111111110100010101011110001001",
			5538 => "00000000000000000101011110001001",
			5539 => "11111101010011110101011110001001",
			5540 => "0000000000000000000100010100100100",
			5541 => "0000000000000000000110001000000100",
			5542 => "11111110011001010101011110001001",
			5543 => "0000000110000000001101111100010000",
			5544 => "0000001101000000000100001000001000",
			5545 => "0000000011000000001100101100000100",
			5546 => "00000001000101000101011110001001",
			5547 => "11111111111101110101011110001001",
			5548 => "0000001011000000000101101100000100",
			5549 => "00000010011100010101011110001001",
			5550 => "00000000110101110101011110001001",
			5551 => "0000000100000000000110001100001000",
			5552 => "0000001100000000001001110000000100",
			5553 => "11111111101011100101011110001001",
			5554 => "00000001110110000101011110001001",
			5555 => "0000000111000000001100001000000100",
			5556 => "00000000011100110101011110001001",
			5557 => "00000000111001100101011110001001",
			5558 => "0000000100000000000100111000011000",
			5559 => "0000000100000000000011010100001100",
			5560 => "0000001001000000001011101000001000",
			5561 => "0000001111000000001001010100000100",
			5562 => "00000010010100100101011110001001",
			5563 => "00000000110001100101011110001001",
			5564 => "00000010111110010101011110001001",
			5565 => "0000000111000000000111111000000100",
			5566 => "00000000000000000101011110001001",
			5567 => "0000000100000000000000101100000100",
			5568 => "00000001011100010101011110001001",
			5569 => "00000000100001110101011110001001",
			5570 => "11111110011011110101011110001001",
			5571 => "0000001000000000001001101000001100",
			5572 => "0000000001000000001011101000001000",
			5573 => "0000000001000000001011101000000100",
			5574 => "11111110011011000101011110001001",
			5575 => "00000011011001000101011110001001",
			5576 => "11111110010101100101011110001001",
			5577 => "0000000100000000000010010000101000",
			5578 => "0000001000000000000110001000010100",
			5579 => "0000000001000000001110010100001000",
			5580 => "0000000100000000001110111000000100",
			5581 => "00000011110011000101011110001001",
			5582 => "11111110011101000101011110001001",
			5583 => "0000001100000000000001011000001000",
			5584 => "0000001000000000001001101000000100",
			5585 => "00000000111011100101011110001001",
			5586 => "11111110010101100101011110001001",
			5587 => "00000010001101000101011110001001",
			5588 => "0000001111000000001111100000010000",
			5589 => "0000001100000000001000000000001000",
			5590 => "0000001001000000001010011000000100",
			5591 => "00000010110010110101011110001001",
			5592 => "11111111100100000101011110001001",
			5593 => "0000000100000000000011110100000100",
			5594 => "00000100100011010101011110001001",
			5595 => "00000000111101100101011110001001",
			5596 => "11111110101110100101011110001001",
			5597 => "0000000100000000000000000000001000",
			5598 => "0000000100000000001010101000000100",
			5599 => "11111110011111100101011110001001",
			5600 => "11111111010001010101011110001001",
			5601 => "11111110010101010101011110001001",
			5602 => "0000000111000000001101111001100000",
			5603 => "0000000100000000000110110001000100",
			5604 => "0000000110000000000001000100001000",
			5605 => "0000000110000000000001000100000100",
			5606 => "11111110010110000101100010111101",
			5607 => "11111111101101010101100010111101",
			5608 => "0000001110000000000110000100100000",
			5609 => "0000001001000000001101101000010000",
			5610 => "0000000100000000001110111000001000",
			5611 => "0000000110000000001101111100000100",
			5612 => "00000001000011000101100010111101",
			5613 => "00000000001100110101100010111101",
			5614 => "0000001001000000000110101000000100",
			5615 => "00000001000001110101100010111101",
			5616 => "00000001101000010101100010111101",
			5617 => "0000000101000000000000001100001000",
			5618 => "0000000100000000000010111000000100",
			5619 => "00000101000011010101100010111101",
			5620 => "00000010111101000101100010111101",
			5621 => "0000000100000000000011110000000100",
			5622 => "00000001000000110101100010111101",
			5623 => "00000010010100010101100010111101",
			5624 => "0000001100000000001000111100010000",
			5625 => "0000000110000000001011001100001000",
			5626 => "0000000111000000000100000000000100",
			5627 => "11111111110000000101100010111101",
			5628 => "00000000101001000101100010111101",
			5629 => "0000000111000000001101100000000100",
			5630 => "11111110101001100101100010111101",
			5631 => "00000000010100100101100010111101",
			5632 => "0000001001000000000100110100001000",
			5633 => "0000000110000000001010011000000100",
			5634 => "00000000011011110101100010111101",
			5635 => "00000001011010100101100010111101",
			5636 => "11111110010001110101100010111101",
			5637 => "0000000110000000001100011000001000",
			5638 => "0000001011000000001100001000000100",
			5639 => "11111110010100000101100010111101",
			5640 => "11111110111101100101100010111101",
			5641 => "0000000111000000000100010100000100",
			5642 => "00000001101101000101100010111101",
			5643 => "0000000100000000000001001100000100",
			5644 => "00000000100100110101100010111101",
			5645 => "0000001001000000000010001100001000",
			5646 => "0000001001000000000000011000000100",
			5647 => "11111110011110110101100010111101",
			5648 => "11111111110011010101100010111101",
			5649 => "11111110001110100101100010111101",
			5650 => "0000001000000000001001101000001100",
			5651 => "0000001100000000000110000100001000",
			5652 => "0000000111000000000100001000000100",
			5653 => "11111110100011110101100010111101",
			5654 => "00000001100010010101100010111101",
			5655 => "11111110010100010101100010111101",
			5656 => "0000000100000000000010010000101100",
			5657 => "0000001000000000001111001000011000",
			5658 => "0000001111000000001000000100001100",
			5659 => "0000000100000000000100001100001000",
			5660 => "0000001001000000000111101100000100",
			5661 => "00000011000110110101100010111101",
			5662 => "11111111011010100101100010111101",
			5663 => "11111110011001000101100010111101",
			5664 => "0000001000000000001001101000000100",
			5665 => "00000000000000000101100010111101",
			5666 => "0000000111000000000111110000000100",
			5667 => "11111110010100000101100010111101",
			5668 => "00000000000000000101100010111101",
			5669 => "0000001100000000000110000100000100",
			5670 => "11111110101110010101100010111101",
			5671 => "0000001111000000000000010100001000",
			5672 => "0000001101000000001100000000000100",
			5673 => "00000001010110110101100010111101",
			5674 => "00000011101010110101100010111101",
			5675 => "0000000110000000000100101100000100",
			5676 => "11111110000111010101100010111101",
			5677 => "00000001011101100101100010111101",
			5678 => "11111110010101100101100010111101",
			5679 => "0000000100000000000011011001110100",
			5680 => "0000000000000000001100001001001100",
			5681 => "0000000100000000001011101100011100",
			5682 => "0000001000000000000110011100011000",
			5683 => "0000000100000000000000010000001100",
			5684 => "0000000011000000001010111000001000",
			5685 => "0000000001000000001100110100000100",
			5686 => "11111110011001000101101001100001",
			5687 => "00000001001011110101101001100001",
			5688 => "11111110010100000101101001100001",
			5689 => "0000000001000000000110101000001000",
			5690 => "0000000111000000001100001000000100",
			5691 => "00000000000011000101101001100001",
			5692 => "00000010000100000101101001100001",
			5693 => "11111110100110000101101001100001",
			5694 => "11111101110001110101101001100001",
			5695 => "0000001000000000000101000100010000",
			5696 => "0000001011000000000001111100001100",
			5697 => "0000001101000000000001111100001000",
			5698 => "0000000011000000000000001100000100",
			5699 => "00000001011010000101101001100001",
			5700 => "11111110101111110101101001100001",
			5701 => "00000010010110100101101001100001",
			5702 => "11111110011111010101101001100001",
			5703 => "0000000010000000001110101000010000",
			5704 => "0000000100000000000100001100001000",
			5705 => "0000000001000000001100110100000100",
			5706 => "11111111111010010101101001100001",
			5707 => "11111101111111010101101001100001",
			5708 => "0000000011000000000000111000000100",
			5709 => "00000001100001010101101001100001",
			5710 => "11111101010111100101101001100001",
			5711 => "0000000001000000000110000000001000",
			5712 => "0000000011000000001011000100000100",
			5713 => "11111111101010110101101001100001",
			5714 => "11111110001101110101101001100001",
			5715 => "0000000011000000001100001000000100",
			5716 => "00000000111010100101101001100001",
			5717 => "00000000000101010101101001100001",
			5718 => "0000001110000000000000101000011100",
			5719 => "0000001011000000000111111000001100",
			5720 => "0000000101000000001000111100001000",
			5721 => "0000000101000000001000111100000100",
			5722 => "00000001110100100101101001100001",
			5723 => "00000000101010000101101001100001",
			5724 => "11111110110001000101101001100001",
			5725 => "0000001000000000001000110000001100",
			5726 => "0000000111000000000000101000000100",
			5727 => "00000001111000000101101001100001",
			5728 => "0000001110000000000000111000000100",
			5729 => "11111111101111010101101001100001",
			5730 => "00000001101100010101101001100001",
			5731 => "00000000000000000101101001100001",
			5732 => "0000001110000000000100000000000100",
			5733 => "11111100101011110101101001100001",
			5734 => "0000000001000000000010001100000100",
			5735 => "00000001101111010101101001100001",
			5736 => "11111111100010100101101001100001",
			5737 => "0000001111000000001001010100110000",
			5738 => "0000000001000000001110100000100100",
			5739 => "0000000111000000000111111000010000",
			5740 => "0000001110000000000111000100001000",
			5741 => "0000000111000000000111111000000100",
			5742 => "11111110011101110101101001100001",
			5743 => "00000000000000000101101001100001",
			5744 => "0000001011000000001110111100000100",
			5745 => "11111110110110110101101001100001",
			5746 => "11111100001001000101101001100001",
			5747 => "0000000100000000001101110100000100",
			5748 => "00000001000101110101101001100001",
			5749 => "0000000010000000001001010000001000",
			5750 => "0000001110000000001011010100000100",
			5751 => "11111110011011010101101001100001",
			5752 => "00000000110011110101101001100001",
			5753 => "0000000010000000000010011100000100",
			5754 => "11111100011001100101101001100001",
			5755 => "11111111000010000101101001100001",
			5756 => "0000001100000000000000101000000100",
			5757 => "11111010101000110101101001100001",
			5758 => "0000000011000000001100101100000100",
			5759 => "00000001010011110101101001100001",
			5760 => "00000000000000000101101001100001",
			5761 => "0000000111000000001101111000011000",
			5762 => "0000000010000000001100010000001000",
			5763 => "0000000011000000001101111000000100",
			5764 => "00000010000001000101101001100001",
			5765 => "11111101111001010101101001100001",
			5766 => "0000000000000000001100001000000100",
			5767 => "11111111010000100101101001100001",
			5768 => "0000000100000000000001001100001000",
			5769 => "0000000111000000001001110000000100",
			5770 => "00000001011001100101101001100001",
			5771 => "00000010011111110101101001100001",
			5772 => "11111111011010010101101001100001",
			5773 => "0000001000000000001010101100000100",
			5774 => "11111110010111110101101001100001",
			5775 => "0000001100000000001001110100001100",
			5776 => "0000000101000000000110110100001000",
			5777 => "0000001110000000000001111100000100",
			5778 => "00000000000000000101101001100001",
			5779 => "11111110111011000101101001100001",
			5780 => "00000001100010100101101001100001",
			5781 => "0000001110000000001011111000000100",
			5782 => "00000000000000000101101001100001",
			5783 => "11111110101001110101101001100001",
			5784 => "0000000111000000001101111001100000",
			5785 => "0000000100000000000110110001001000",
			5786 => "0000000110000000000001000100001000",
			5787 => "0000000110000000000001000100000100",
			5788 => "11111110010101000101101110011101",
			5789 => "11111111100111100101101110011101",
			5790 => "0000001110000000001000111100100000",
			5791 => "0000000111000000001011000100010000",
			5792 => "0000000011000000001100001000001000",
			5793 => "0000001100000000000000110000000100",
			5794 => "11111111110111000101101110011101",
			5795 => "00000001100001100101101110011101",
			5796 => "0000001001000000000010001100000100",
			5797 => "11111110011111100101101110011101",
			5798 => "00000000111000110101101110011101",
			5799 => "0000000010000000001001011100001000",
			5800 => "0000000110000000000001111000000100",
			5801 => "00000001111000110101101110011101",
			5802 => "00000001001001100101101110011101",
			5803 => "0000000000000000000000111000000100",
			5804 => "00000011011110000101101110011101",
			5805 => "00000001111100000101101110011101",
			5806 => "0000000100000000000010111000010000",
			5807 => "0000001100000000001000111100001000",
			5808 => "0000001010000000000110011000000100",
			5809 => "00000000011100010101101110011101",
			5810 => "11111111010000110101101110011101",
			5811 => "0000001001000000001101111100000100",
			5812 => "00000001100100110101101110011101",
			5813 => "11111110010010110101101110011101",
			5814 => "0000000110000000001001100100001000",
			5815 => "0000001001000000001101101000000100",
			5816 => "00000000110000110101101110011101",
			5817 => "00000001011100110101101110011101",
			5818 => "0000001100000000001000111000000100",
			5819 => "11111110111111110101101110011101",
			5820 => "00000001010110110101101110011101",
			5821 => "0000000110000000001100011000000100",
			5822 => "11111110010011100101101110011101",
			5823 => "0000000111000000000100010100000100",
			5824 => "00000001111000110101101110011101",
			5825 => "0000000100000000000001001100000100",
			5826 => "00000000101100100101101110011101",
			5827 => "0000001001000000000010001100001000",
			5828 => "0000001001000000000000011000000100",
			5829 => "11111110011100010101101110011101",
			5830 => "11111111110000100101101110011101",
			5831 => "11111110001110100101101110011101",
			5832 => "0000001000000000001001101000001100",
			5833 => "0000001100000000000110000100001000",
			5834 => "0000000111000000000100001000000100",
			5835 => "11111110100000010101101110011101",
			5836 => "00000001110110000101101110011101",
			5837 => "11111110010011000101101110011101",
			5838 => "0000000100000000000010010000110000",
			5839 => "0000001000000000001111001000011000",
			5840 => "0000001111000000001000000100001100",
			5841 => "0000000100000000000100001100001000",
			5842 => "0000000100000000000011001100000100",
			5843 => "11111111101110100101101110011101",
			5844 => "00000011110010000101101110011101",
			5845 => "11111110010111100101101110011101",
			5846 => "0000001000000000001001101000000100",
			5847 => "00000000000000000101101110011101",
			5848 => "0000000111000000000111110000000100",
			5849 => "11111110010010110101101110011101",
			5850 => "00000000000000000101101110011101",
			5851 => "0000001000000000001010101100010000",
			5852 => "0000000100000000000011011000001000",
			5853 => "0000000100000000001001001100000100",
			5854 => "11111111010111000101101110011101",
			5855 => "00000001110010100101101110011101",
			5856 => "0000000000000000000000110000000100",
			5857 => "00000000000000000101101110011101",
			5858 => "11111101111111110101101110011101",
			5859 => "0000000001000000000000111100000100",
			5860 => "00000001011010000101101110011101",
			5861 => "00000011010001110101101110011101",
			5862 => "11111110010100010101101110011101",
			5863 => "0000001011000000000000001101101100",
			5864 => "0000000001000000000000011000011000",
			5865 => "0000000110000000001101111100001100",
			5866 => "0000000100000000001011100000001000",
			5867 => "0000000100000000000011010100000100",
			5868 => "11111110100010010101110100011001",
			5869 => "00000000000101000101110100011001",
			5870 => "11111110010001000101110100011001",
			5871 => "0000001101000000000011011100001000",
			5872 => "0000000011000000001000110000000100",
			5873 => "00000010000100000101110100011001",
			5874 => "11111111000110110101110100011001",
			5875 => "11111110010000100101110100011001",
			5876 => "0000001110000000001100001000100100",
			5877 => "0000000110000000000001000100000100",
			5878 => "11111110010010000101110100011001",
			5879 => "0000001101000000001100101100010000",
			5880 => "0000000011000000001001110000001000",
			5881 => "0000001011000000000111111000000100",
			5882 => "00000001000001100101110100011001",
			5883 => "00000001111000110101110100011001",
			5884 => "0000000000000000001011000100000100",
			5885 => "00000000101010100101110100011001",
			5886 => "00000010001111110101110100011001",
			5887 => "0000000110000000000001111000001000",
			5888 => "0000001110000000000111111000000100",
			5889 => "00000010110001010101110100011001",
			5890 => "00000011010011110101110100011001",
			5891 => "0000001111000000000100000100000100",
			5892 => "00000000111010110101110100011001",
			5893 => "00000010001010010101110100011001",
			5894 => "0000000100000000001010110100010100",
			5895 => "0000000110000000001011111100000100",
			5896 => "11111110010011100101110100011001",
			5897 => "0000000110000000001101111100001000",
			5898 => "0000001111000000000110110100000100",
			5899 => "11111111110110010101110100011001",
			5900 => "00000001101010100101110100011001",
			5901 => "0000000000000000001010000000000100",
			5902 => "00000000001000100101110100011001",
			5903 => "00000011001110000101110100011001",
			5904 => "0000000110000000001001100100010000",
			5905 => "0000001011000000001100001000001000",
			5906 => "0000000101000000001101100000000100",
			5907 => "11111110100010000101110100011001",
			5908 => "00000000110000100101110100011001",
			5909 => "0000000100000000000100001100000100",
			5910 => "00000001011101010101110100011001",
			5911 => "00000010001111100101110100011001",
			5912 => "0000001111000000000010000100001000",
			5913 => "0000001111000000001100100100000100",
			5914 => "11111111111000110101110100011001",
			5915 => "11111110100100010101110100011001",
			5916 => "00000001000000110101110100011001",
			5917 => "0000001100000000001110001100101100",
			5918 => "0000001111000000000101110000010000",
			5919 => "0000000101000000001000000000000100",
			5920 => "00000000000110010101110100011001",
			5921 => "0000001111000000001110000100000100",
			5922 => "11111110010010100101110100011001",
			5923 => "0000001011000000000100001000000100",
			5924 => "00000001001000110101110100011001",
			5925 => "11111110010010000101110100011001",
			5926 => "0000001001000000000100110100010100",
			5927 => "0000000100000000000001001100010000",
			5928 => "0000001111000000000010000100001000",
			5929 => "0000001101000000000111010000000100",
			5930 => "00000010111001010101110100011001",
			5931 => "11111111100011100101110100011001",
			5932 => "0000000000000000000000111000000100",
			5933 => "00000100010011000101110100011001",
			5934 => "00000001101111010101110100011001",
			5935 => "11111110100000010101110100011001",
			5936 => "0000000000000000000111111000000100",
			5937 => "11111110001100010101110100011001",
			5938 => "00000000011011010101110100011001",
			5939 => "0000001000000000001001101000000100",
			5940 => "11111110010000100101110100011001",
			5941 => "0000000100000000000110110000100000",
			5942 => "0000001110000000001101101100010000",
			5943 => "0000000100000000000011101100001000",
			5944 => "0000001001000000000100101100000100",
			5945 => "00000011010001000101110100011001",
			5946 => "00000000011101110101110100011001",
			5947 => "0000001010000000000110011100000100",
			5948 => "11111110101110010101110100011001",
			5949 => "00000011010111100101110100011001",
			5950 => "0000000110000000000100101100001000",
			5951 => "0000001100000000001011011100000100",
			5952 => "11111110010101000101110100011001",
			5953 => "00000001100011110101110100011001",
			5954 => "0000001000000000000001110100000100",
			5955 => "11111111011010000101110100011001",
			5956 => "00000010100001100101110100011001",
			5957 => "11111110010000100101110100011001",
			5958 => "0000000111000000001110001110000000",
			5959 => "0000000100000000000110110001100000",
			5960 => "0000000011000000000100010100100000",
			5961 => "0000001100000000000000110000010000",
			5962 => "0000000010000000000110100000000100",
			5963 => "00000000011011010101111010101101",
			5964 => "0000001111000000000100000100001000",
			5965 => "0000000101000000001000111100000100",
			5966 => "00000001010101000101111010101101",
			5967 => "11111101000110100101111010101101",
			5968 => "00000001010111100101111010101101",
			5969 => "0000001010000000000111110100000100",
			5970 => "11111110000110010101111010101101",
			5971 => "0000001111000000000111010000001000",
			5972 => "0000000010000000001001010000000100",
			5973 => "00000000111001010101111010101101",
			5974 => "11111110101100100101111010101101",
			5975 => "00000010000111000101111010101101",
			5976 => "0000001001000000000010001100100000",
			5977 => "0000000011000000001100001000010000",
			5978 => "0000001011000000001110111100001000",
			5979 => "0000000011000000001011000100000100",
			5980 => "00000001001110110101111010101101",
			5981 => "11111101010000000101111010101101",
			5982 => "0000000010000000001111010000000100",
			5983 => "11111111000110010101111010101101",
			5984 => "00000000111001100101111010101101",
			5985 => "0000001111000000000101100100001000",
			5986 => "0000000101000000000011011100000100",
			5987 => "11111011110011100101111010101101",
			5988 => "11111101111110100101111010101101",
			5989 => "0000001001000000000010001100000100",
			5990 => "11111101010101010101111010101101",
			5991 => "11111111100111110101111010101101",
			5992 => "0000000011000000001001110000010000",
			5993 => "0000001111000000000101100100001000",
			5994 => "0000001010000000001001000100000100",
			5995 => "00000000110111100101111010101101",
			5996 => "00000000000000010101111010101101",
			5997 => "0000001001000000001001111000000100",
			5998 => "00000000101010110101111010101101",
			5999 => "00000001100010010101111010101101",
			6000 => "0000001101000000001100101100001000",
			6001 => "0000001001000000000110101000000100",
			6002 => "11111111100000100101111010101101",
			6003 => "00000000110100010101111010101101",
			6004 => "0000001100000000001010000000000100",
			6005 => "00000010110101000101111010101101",
			6006 => "00000000001110010101111010101101",
			6007 => "0000000110000000001100011000001000",
			6008 => "0000001101000000000110000100000100",
			6009 => "11111110010101100101111010101101",
			6010 => "11111111110000110101111010101101",
			6011 => "0000000111000000000100010100000100",
			6012 => "00000001010111110101111010101101",
			6013 => "0000001010000000000001110000001000",
			6014 => "0000001100000000000011011100000100",
			6015 => "00000000100010110101111010101101",
			6016 => "11111111010001010101111010101101",
			6017 => "0000001100000000000000101000000100",
			6018 => "11111101000001000101111010101101",
			6019 => "0000000011000000001110001100000100",
			6020 => "00000000000001100101111010101101",
			6021 => "11111110100000010101111010101101",
			6022 => "0000001000000000001001101000010000",
			6023 => "0000000001000000001011101000001100",
			6024 => "0000001001000000000001111000000100",
			6025 => "11111110010110010101111010101101",
			6026 => "0000000010000000000111100000000100",
			6027 => "11111110110011100101111010101101",
			6028 => "00000010000101010101111010101101",
			6029 => "11111110011000110101111010101101",
			6030 => "0000000100000000000011111000101100",
			6031 => "0000001100000000000110000100010000",
			6032 => "0000000100000000000000101100001000",
			6033 => "0000001010000000000110011000000100",
			6034 => "00000000000000000101111010101101",
			6035 => "11111110000011010101111010101101",
			6036 => "0000000001000000001101011100000100",
			6037 => "11111110111111100101111010101101",
			6038 => "00000000111101100101111010101101",
			6039 => "0000000001000000001011101000001100",
			6040 => "0000000101000000001001010100001000",
			6041 => "0000001011000000001110110000000100",
			6042 => "00000001101100000101111010101101",
			6043 => "00000011100001100101111010101101",
			6044 => "11111110111000100101111010101101",
			6045 => "0000001100000000000001011000001000",
			6046 => "0000001001000000000111101100000100",
			6047 => "00000000100001000101111010101101",
			6048 => "11111111001000000101111010101101",
			6049 => "0000000001000000000100110100000100",
			6050 => "11111111100011010101111010101101",
			6051 => "00000001111001110101111010101101",
			6052 => "0000000100000000000000000000001100",
			6053 => "0000001100000000000000001100001000",
			6054 => "0000001000000000001101010000000100",
			6055 => "11111111110001110101111010101101",
			6056 => "00000010101110000101111010101101",
			6057 => "11111110100001100101111010101101",
			6058 => "11111110011001010101111010101101",
			6059 => "0000000011000000000000110001001000",
			6060 => "0000001110000000000001110100111100",
			6061 => "0000000011000000000011111100100100",
			6062 => "0000000010000000000000110100001000",
			6063 => "0000001111000000000101101100000100",
			6064 => "00000000000000000110000001100001",
			6065 => "00000001101011110110000001100001",
			6066 => "0000001111000000001010111000001100",
			6067 => "0000000110000000001100011000001000",
			6068 => "0000001111000000001010111000000100",
			6069 => "11111110011001010110000001100001",
			6070 => "00000000000000000110000001100001",
			6071 => "00000000000000000110000001100001",
			6072 => "0000001100000000000111111000001000",
			6073 => "0000000000000000000100000000000100",
			6074 => "00000000111100100110000001100001",
			6075 => "11111111000101010110000001100001",
			6076 => "0000000100000000001110011000000100",
			6077 => "00000001100001000110000001100001",
			6078 => "00000000000000000110000001100001",
			6079 => "0000001101000000001000111100001000",
			6080 => "0000001011000000001010000000000100",
			6081 => "11111110101111110110000001100001",
			6082 => "11111010100110110110000001100001",
			6083 => "0000001011000000000100010100001000",
			6084 => "0000000111000000001010000000000100",
			6085 => "00000000000000000110000001100001",
			6086 => "11111110111100000110000001100001",
			6087 => "0000000100000000001010101000000100",
			6088 => "00000001000110110110000001100001",
			6089 => "00000000000000000110000001100001",
			6090 => "0000000110000000001110010100000100",
			6091 => "11111110101000010110000001100001",
			6092 => "0000000010000000001001010000000100",
			6093 => "00000001110010000110000001100001",
			6094 => "11111111111011010110000001100001",
			6095 => "0000001111000000000110100100111000",
			6096 => "0000000110000000000001111000011000",
			6097 => "0000001101000000001100110000001000",
			6098 => "0000000011000000000111111000000100",
			6099 => "00000000011011000110000001100001",
			6100 => "11111110000100100110000001100001",
			6101 => "0000000111000000001011000100001000",
			6102 => "0000001001000000001001111000000100",
			6103 => "00000001010011010110000001100001",
			6104 => "11111110101110000110000001100001",
			6105 => "0000000000000000000110001000000100",
			6106 => "11111111101111110110000001100001",
			6107 => "00000001101100000110000001100001",
			6108 => "0000001011000000000111111000000100",
			6109 => "00000000110000000110000001100001",
			6110 => "0000000000000000001011000100001100",
			6111 => "0000000100000000000000010100001000",
			6112 => "0000000010000000001110101100000100",
			6113 => "11111101110010010110000001100001",
			6114 => "00000000000000000110000001100001",
			6115 => "11111100011011010110000001100001",
			6116 => "0000001111000000000110100100001000",
			6117 => "0000000000000000000110000100000100",
			6118 => "00000001100000100110000001100001",
			6119 => "00000000000000000110000001100001",
			6120 => "0000000110000000000100110100000100",
			6121 => "00000000000000000110000001100001",
			6122 => "11111101001110010110000001100001",
			6123 => "0000000011000000001011000100100000",
			6124 => "0000001000000000001001101000001000",
			6125 => "0000000011000000000100010100000100",
			6126 => "11111100000110110110000001100001",
			6127 => "00000000000000000110000001100001",
			6128 => "0000000100000000000000010100001000",
			6129 => "0000001100000000000100010100000100",
			6130 => "00000001110010010110000001100001",
			6131 => "11111111001000100110000001100001",
			6132 => "0000000000000000000100010100001000",
			6133 => "0000001111000000001010001100000100",
			6134 => "11111110010011000110000001100001",
			6135 => "00000000110110010110000001100001",
			6136 => "0000000111000000000111111000000100",
			6137 => "11111111100110010110000001100001",
			6138 => "00000000111111110110000001100001",
			6139 => "0000001001000000001001111000011100",
			6140 => "0000000010000000001110000100001100",
			6141 => "0000001110000000000010011000000100",
			6142 => "00000000111110100110000001100001",
			6143 => "0000000100000000001101001000000100",
			6144 => "11111111101100010110000001100001",
			6145 => "11111101110011000110000001100001",
			6146 => "0000000011000000001100001000001000",
			6147 => "0000000010000000000010011100000100",
			6148 => "00000001100110100110000001100001",
			6149 => "11111111110000010110000001100001",
			6150 => "0000001111000000000101100100000100",
			6151 => "11111110001001010110000001100001",
			6152 => "11111111101101010110000001100001",
			6153 => "0000001110000000001101111000010000",
			6154 => "0000001111000000000010110100001000",
			6155 => "0000001100000000000000110000000100",
			6156 => "11111110101001100110000001100001",
			6157 => "00000000000011110110000001100001",
			6158 => "0000001010000000000110011000000100",
			6159 => "00000010010101010110000001100001",
			6160 => "00000000010100110110000001100001",
			6161 => "0000000111000000001000111000001000",
			6162 => "0000000111000000000100000000000100",
			6163 => "11111111110101100110000001100001",
			6164 => "11111111000110000110000001100001",
			6165 => "0000001111000000000111110000000100",
			6166 => "00000010001001110110000001100001",
			6167 => "11111111111101010110000001100001",
			6168 => "0000000101000000001000000010001000",
			6169 => "0000000001000000000000011000010100",
			6170 => "0000000110000000001101111100001000",
			6171 => "0000000010000000000101110100000100",
			6172 => "11111111010011010110001000101101",
			6173 => "11111110001010100110001000101101",
			6174 => "0000000001000000001100100000000100",
			6175 => "11111110001100000110001000101101",
			6176 => "0000000111000000000111111000000100",
			6177 => "11111111100000010110001000101101",
			6178 => "00000011111100010110001000101101",
			6179 => "0000001110000000001101100000110100",
			6180 => "0000000000000000001010000000011100",
			6181 => "0000001110000000000111111000001100",
			6182 => "0000000110000000000001000100000100",
			6183 => "11111110010010110110001000101101",
			6184 => "0000001010000000000001010000000100",
			6185 => "00000011001101100110001000101101",
			6186 => "11111111100110110110001000101101",
			6187 => "0000000111000000001011000100001000",
			6188 => "0000000110000000000100110100000100",
			6189 => "00000001001011000110001000101101",
			6190 => "11111111010111010110001000101101",
			6191 => "0000000010000000000101110000000100",
			6192 => "00000001101110010110001000101101",
			6193 => "00000010111011110110001000101101",
			6194 => "0000001100000000000000110000001000",
			6195 => "0000000010000000000001000000000100",
			6196 => "00000010000111110110001000101101",
			6197 => "11111110110101100110001000101101",
			6198 => "0000000101000000000110000100001000",
			6199 => "0000001110000000000100010100000100",
			6200 => "00000011000101100110001000101101",
			6201 => "00000010000011010110001000101101",
			6202 => "0000001011000000000101101100000100",
			6203 => "00000011100011010110001000101101",
			6204 => "11111110011010110110001000101101",
			6205 => "0000000000000000000000110000100000",
			6206 => "0000000010000000001010001000010000",
			6207 => "0000000111000000000100000000001000",
			6208 => "0000001110000000001100101000000100",
			6209 => "11111111100100000110001000101101",
			6210 => "11111110000111100110001000101101",
			6211 => "0000000010000000000010110100000100",
			6212 => "11111110010001100110001000101101",
			6213 => "00000000111011000110001000101101",
			6214 => "0000000110000000000100110100001000",
			6215 => "0000000101000000001101111000000100",
			6216 => "00000000100011110110001000101101",
			6217 => "00000101011101000110001000101101",
			6218 => "0000001100000000000100000000000100",
			6219 => "00000000001101100110001000101101",
			6220 => "00000010001110110110001000101101",
			6221 => "0000000110000000001001100100010000",
			6222 => "0000001100000000000100000000001000",
			6223 => "0000000000000000000111111000000100",
			6224 => "00000001100100010110001000101101",
			6225 => "00000010110110110110001000101101",
			6226 => "0000000001000000001001111000000100",
			6227 => "00000011001111000110001000101101",
			6228 => "00000100010110100110001000101101",
			6229 => "0000000111000000001101100000001000",
			6230 => "0000000010000000001000001100000100",
			6231 => "11111110001000000110001000101101",
			6232 => "11111111100110010110001000101101",
			6233 => "0000000110000000001111000000000100",
			6234 => "00000100100001100110001000101101",
			6235 => "11111111010000100110001000101101",
			6236 => "0000000111000000001101111000111000",
			6237 => "0000001110000000000001101000010100",
			6238 => "0000000101000000001000000000001000",
			6239 => "0000000011000000001110110000000100",
			6240 => "11111110011111110110001000101101",
			6241 => "00000001110001110110001000101101",
			6242 => "0000000010000000000010000000000100",
			6243 => "11111110001111100110001000101101",
			6244 => "0000000000000000001000111100000100",
			6245 => "00000010110111110110001000101101",
			6246 => "11111110010110000110001000101101",
			6247 => "0000001001000000000001111000011000",
			6248 => "0000000111000000001101100000001100",
			6249 => "0000000110000000001011001100000100",
			6250 => "00000001110111010110001000101101",
			6251 => "0000000001000000000111100100000100",
			6252 => "00000001000011000110001000101101",
			6253 => "11111110010100110110001000101101",
			6254 => "0000000000000000001010101100000100",
			6255 => "11111110001111010110001000101101",
			6256 => "0000001000000000000010101000000100",
			6257 => "00000011100011010110001000101101",
			6258 => "11111111100010110110001000101101",
			6259 => "0000000000000000000111111000001000",
			6260 => "0000001100000000001110001100000100",
			6261 => "11111110001000110110001000101101",
			6262 => "00000001001111100110001000101101",
			6263 => "00000010000000100110001000101101",
			6264 => "0000001001000000001000010100100000",
			6265 => "0000001000000000001001101000001100",
			6266 => "0000001100000000000110000100001000",
			6267 => "0000001100000000000110000100000100",
			6268 => "11111110010011000110001000101101",
			6269 => "00000000110001110110001000101101",
			6270 => "11111110001001110110001000101101",
			6271 => "0000000000000000001000111100010000",
			6272 => "0000001000000000001111001000001000",
			6273 => "0000001001000000001010011000000100",
			6274 => "00000011101111110110001000101101",
			6275 => "11111110011010100110001000101101",
			6276 => "0000000010000000001110111000000100",
			6277 => "00000010000010000110001000101101",
			6278 => "11111111010100110110001000101101",
			6279 => "11111110001010000110001000101101",
			6280 => "0000000111000000000101110100000100",
			6281 => "11111110001100010110001000101101",
			6282 => "00000010000111110110001000101101",
			6283 => "0000000101000000001000000010001100",
			6284 => "0000000001000000000000011000011100",
			6285 => "0000000001000000001100100000000100",
			6286 => "11111110001100100110001111111001",
			6287 => "0000001111000000001000000000001100",
			6288 => "0000000111000000000111111000000100",
			6289 => "11111111110100000110001111111001",
			6290 => "0000000010000000001101000100000100",
			6291 => "00000011110100000110001111111001",
			6292 => "00000001011010000110001111111001",
			6293 => "0000000010000000001001010000001000",
			6294 => "0000000000000000000111111000000100",
			6295 => "11111110000001110110001111111001",
			6296 => "00000000010011100110001111111001",
			6297 => "11111110001010110110001111111001",
			6298 => "0000000100000000001001001100111100",
			6299 => "0000000011000000000101101100011100",
			6300 => "0000000011000000000100000000001100",
			6301 => "0000001000000000000101000100000100",
			6302 => "11111111100110010110001111111001",
			6303 => "0000001010000000000001010000000100",
			6304 => "00000010110010010110001111111001",
			6305 => "00000000011010010110001111111001",
			6306 => "0000001011000000001100001000001000",
			6307 => "0000001111000000000111110000000100",
			6308 => "00000001010000000110001111111001",
			6309 => "00000011110111000110001111111001",
			6310 => "0000001000000000000001010100000100",
			6311 => "00000100000000100110001111111001",
			6312 => "00000010001010100110001111111001",
			6313 => "0000000111000000000100000000010000",
			6314 => "0000000011000000001101111000001000",
			6315 => "0000001101000000001100101000000100",
			6316 => "00000000110111110110001111111001",
			6317 => "00000011000010110110001111111001",
			6318 => "0000001010000000000001010000000100",
			6319 => "00000000000011010110001111111001",
			6320 => "11111110110000110110001111111001",
			6321 => "0000000001000000000110101000001000",
			6322 => "0000000100000000000000010000000100",
			6323 => "11111110011011110110001111111001",
			6324 => "00000001100101110110001111111001",
			6325 => "0000000010000000000111011000000100",
			6326 => "11111110010001000110001111111001",
			6327 => "00000000000111100110001111111001",
			6328 => "0000000011000000000001101000100000",
			6329 => "0000000111000000001100001000010000",
			6330 => "0000000000000000000100010100001000",
			6331 => "0000000011000000001000111100000100",
			6332 => "00000010100110000110001111111001",
			6333 => "00000001011100000110001111111001",
			6334 => "0000000100000000000000100000000100",
			6335 => "00000010110000100110001111111001",
			6336 => "00000001011111010110001111111001",
			6337 => "0000000100000000000110110000001000",
			6338 => "0000000100000000000100001100000100",
			6339 => "00000010100100110110001111111001",
			6340 => "00000011000100110110001111111001",
			6341 => "0000000011000000000111001000000100",
			6342 => "00000000000000000110001111111001",
			6343 => "11111110011001000110001111111001",
			6344 => "0000001100000000001001110000010000",
			6345 => "0000001010000000001100011100001000",
			6346 => "0000000100000000000100001100000100",
			6347 => "11111111111010110110001111111001",
			6348 => "00000011001110100110001111111001",
			6349 => "0000001111000000000011001000000100",
			6350 => "11111110001110110110001111111001",
			6351 => "00000001011000010110001111111001",
			6352 => "00000010111111000110001111111001",
			6353 => "0000000111000000001101111000110000",
			6354 => "0000001111000000001101000100001000",
			6355 => "0000001101000000001000000000000100",
			6356 => "11111111011110100110001111111001",
			6357 => "11111110010000110110001111111001",
			6358 => "0000000001000000001011101000011100",
			6359 => "0000001010000000000101000100010000",
			6360 => "0000001100000000001000111000001000",
			6361 => "0000001001000000001011111100000100",
			6362 => "00000000100110110110001111111001",
			6363 => "11111110011110000110001111111001",
			6364 => "0000000111000000001101100000000100",
			6365 => "00000000000000010110001111111001",
			6366 => "00000010100101010110001111111001",
			6367 => "0000001101000000000001011000001000",
			6368 => "0000001100000000000110000100000100",
			6369 => "11111110010100010110001111111001",
			6370 => "00000000010110110110001111111001",
			6371 => "00000000111111000110001111111001",
			6372 => "0000001100000000001100110000000100",
			6373 => "11111110001100010110001111111001",
			6374 => "0000001111000000000010000000000100",
			6375 => "11111110011100010110001111111001",
			6376 => "00000001010000000110001111111001",
			6377 => "0000001000000000001001101000001100",
			6378 => "0000000111000000001100101000001000",
			6379 => "0000001100000000000110000100000100",
			6380 => "00000000000000000110001111111001",
			6381 => "11111110100100010110001111111001",
			6382 => "11111110001100100110001111111001",
			6383 => "0000000100000000000010010000011000",
			6384 => "0000001000000000001111001000001100",
			6385 => "0000001001000000001010011000000100",
			6386 => "00000011001010010110001111111001",
			6387 => "0000001100000000001011011100000100",
			6388 => "11111110011001110110001111111001",
			6389 => "00000000111110010110001111111001",
			6390 => "0000001000000000000111000000001000",
			6391 => "0000000100000000000001101100000100",
			6392 => "00000001101110010110001111111001",
			6393 => "11111110001001010110001111111001",
			6394 => "00000100100100000110001111111001",
			6395 => "0000000001000000001001011000000100",
			6396 => "11111110001100010110001111111001",
			6397 => "00000000000001110110001111111001",
			6398 => "0000000101000000000011100010001000",
			6399 => "0000000001000000000000011000011100",
			6400 => "0000000110000000001101111100010000",
			6401 => "0000001001000000001110100000001000",
			6402 => "0000000010000000000101110100000100",
			6403 => "11111111001100000110010111100101",
			6404 => "11111110000111010110010111100101",
			6405 => "0000000010000000001010001000000100",
			6406 => "00000000101010100110010111100101",
			6407 => "11111110011000100110010111100101",
			6408 => "0000001101000000000011011100001000",
			6409 => "0000000111000000000111111000000100",
			6410 => "11111111100110100110010111100101",
			6411 => "00000101000110010110010111100101",
			6412 => "11111110001011100110010111100101",
			6413 => "0000001110000000001000111000110100",
			6414 => "0000001110000000000111111000010100",
			6415 => "0000000110000000000001000100000100",
			6416 => "11111110001110110110010111100101",
			6417 => "0000000111000000001011000100001000",
			6418 => "0000000011000000000000101000000100",
			6419 => "00000100001111010110010111100101",
			6420 => "00000011010000100110010111100101",
			6421 => "0000000110000000000001111000000100",
			6422 => "00000101000011000110010111100101",
			6423 => "00000100010010000110010111100101",
			6424 => "0000000010000000000100101000010000",
			6425 => "0000001101000000000000001100001000",
			6426 => "0000001010000000001001000100000100",
			6427 => "00000010111110010110010111100101",
			6428 => "00000001100010000110010111100101",
			6429 => "0000001111000000001010001100000100",
			6430 => "00000001110110110110010111100101",
			6431 => "00000100101011000110010111100101",
			6432 => "0000000111000000001011000100001000",
			6433 => "0000001010000000001100011100000100",
			6434 => "00000010001110000110010111100101",
			6435 => "00000100100001000110010111100101",
			6436 => "0000001101000000001010111100000100",
			6437 => "00000100110011010110010111100101",
			6438 => "11111110001101010110010111100101",
			6439 => "0000000010000000000111111100011100",
			6440 => "0000001010000000001010110000010000",
			6441 => "0000000110000000001101111100001000",
			6442 => "0000000110000000001110010100000100",
			6443 => "11111110001110010110010111100101",
			6444 => "00000001111001010110010111100101",
			6445 => "0000000110000000001010011000000100",
			6446 => "11111111011110110110010111100101",
			6447 => "00000010010111000110010111100101",
			6448 => "0000001001000000001101101000000100",
			6449 => "00000000010010110110010111100101",
			6450 => "0000000010000000000100101000000100",
			6451 => "00000101100110010110010111100101",
			6452 => "00000011101000000110010111100101",
			6453 => "0000000110000000001001100100010000",
			6454 => "0000001100000000000100000000001000",
			6455 => "0000001110000000000110000100000100",
			6456 => "00000011010100110110010111100101",
			6457 => "00000001011011110110010111100101",
			6458 => "0000001010000000000110011000000100",
			6459 => "00000001110100100110010111100101",
			6460 => "00000100101010000110010111100101",
			6461 => "0000000111000000001101100000001000",
			6462 => "0000000011000000001001001000000100",
			6463 => "00000000000000000110010111100101",
			6464 => "11111110010011110110010111100101",
			6465 => "00000011001000100110010111100101",
			6466 => "0000000111000000001101111001000100",
			6467 => "0000001111000000001110101100001100",
			6468 => "0000001111000000000100010000000100",
			6469 => "11111110001110100110010111100101",
			6470 => "0000001111000000000001001000000100",
			6471 => "11111111100101000110010111100101",
			6472 => "11111110011000000110010111100101",
			6473 => "0000000110000000001011001100011000",
			6474 => "0000001101000000001111011100001100",
			6475 => "0000001000000000001000101100001000",
			6476 => "0000000111000000000101101100000100",
			6477 => "00000010111011000110010111100101",
			6478 => "00000101001010110110010111100101",
			6479 => "11111110100000000110010111100101",
			6480 => "0000001111000000001100010100001000",
			6481 => "0000000110000000001011001100000100",
			6482 => "11111110001101010110010111100101",
			6483 => "00000000000000000110010111100101",
			6484 => "00000001101000010110010111100101",
			6485 => "0000000111000000000101101100010000",
			6486 => "0000000001000000000110101000001000",
			6487 => "0000001110000000000110100100000100",
			6488 => "11111110100111000110010111100101",
			6489 => "00000011010100100110010111100101",
			6490 => "0000000001000000000111100100000100",
			6491 => "11111111000000110110010111100101",
			6492 => "11111110000110000110010111100101",
			6493 => "0000000010000000000000010000001000",
			6494 => "0000000001000000001101101000000100",
			6495 => "00000101000000100110010111100101",
			6496 => "00000001010001010110010111100101",
			6497 => "0000001111000000001001100000000100",
			6498 => "11111110010100100110010111100101",
			6499 => "00000000011111110110010111100101",
			6500 => "0000001001000000001000010100100100",
			6501 => "0000001000000000001001101000001100",
			6502 => "0000001100000000000110000100001000",
			6503 => "0000000010000000000111010100000100",
			6504 => "11111110010010000110010111100101",
			6505 => "00000000110010110110010111100101",
			6506 => "11111110000110100110010111100101",
			6507 => "0000001000000000001101010000010000",
			6508 => "0000001000000000001111001000001000",
			6509 => "0000001001000000001010011000000100",
			6510 => "00000100110100110110010111100101",
			6511 => "11111110010110010110010111100101",
			6512 => "0000000001000000001001011000000100",
			6513 => "11111111011101110110010111100101",
			6514 => "00000010100001110110010111100101",
			6515 => "0000001010000000001100000100000100",
			6516 => "11111111000000100110010111100101",
			6517 => "11111110000110010110010111100101",
			6518 => "0000000111000000000101110100000100",
			6519 => "11111110001000010110010111100101",
			6520 => "00000010100100000110010111100101",
			6521 => "0000000100000000001011101100100000",
			6522 => "0000001000000000000110011100011100",
			6523 => "0000000100000000000000010000010100",
			6524 => "0000001111000000000100000100001100",
			6525 => "0000001111000000001001110100000100",
			6526 => "11111110001001100110011101010001",
			6527 => "0000000110000000000001000100000100",
			6528 => "00000000000000000110011101010001",
			6529 => "00000001101100110110011101010001",
			6530 => "0000000110000000001110010100000100",
			6531 => "11111111100100100110011101010001",
			6532 => "11111110010010100110011101010001",
			6533 => "0000000110000000000001111000000100",
			6534 => "00000001111010110110011101010001",
			6535 => "11111110011101010110011101010001",
			6536 => "11111101110101100110011101010001",
			6537 => "0000001000000000000101000100011000",
			6538 => "0000001011000000000001111100010100",
			6539 => "0000001101000000000001111100010000",
			6540 => "0000000011000000000000001100001100",
			6541 => "0000001101000000000110000100001000",
			6542 => "0000001111000000001010001100000100",
			6543 => "00000000101111100110011101010001",
			6544 => "11111101000111110110011101010001",
			6545 => "00000001111010100110011101010001",
			6546 => "11111110110101100110011101010001",
			6547 => "00000010001111110110011101010001",
			6548 => "11111110100001000110011101010001",
			6549 => "0000000010000000000111111101000000",
			6550 => "0000000010000000000111111100100000",
			6551 => "0000000010000000000100101000010000",
			6552 => "0000000110000000001101111100001000",
			6553 => "0000001100000000000100010100000100",
			6554 => "11111111111010000110011101010001",
			6555 => "00000000011011100110011101010001",
			6556 => "0000001100000000000111111000000100",
			6557 => "00000000010000100110011101010001",
			6558 => "11111111110001000110011101010001",
			6559 => "0000001111000000000110110100001000",
			6560 => "0000000101000000000110000100000100",
			6561 => "00000000000000000110011101010001",
			6562 => "11111100100111000110011101010001",
			6563 => "0000000110000000001100011000000100",
			6564 => "00000001110000100110011101010001",
			6565 => "00000000010001010110011101010001",
			6566 => "0000000001000000001100110100010000",
			6567 => "0000000111000000000100010100001000",
			6568 => "0000000100000000000011010100000100",
			6569 => "11111101111110010110011101010001",
			6570 => "00000001001100010110011101010001",
			6571 => "0000001011000000001100001000000100",
			6572 => "00000010100110100110011101010001",
			6573 => "00000000000000000110011101010001",
			6574 => "0000001001000000000111100100001000",
			6575 => "0000000110000000000100110100000100",
			6576 => "11111100011101010110011101010001",
			6577 => "11111110100101000110011101010001",
			6578 => "0000001000000000000110001000000100",
			6579 => "11111110011011100110011101010001",
			6580 => "11111111110100010110011101010001",
			6581 => "0000000110000000001100011000100000",
			6582 => "0000000101000000000000001100010000",
			6583 => "0000000011000000001001110000001000",
			6584 => "0000000001000000000110000000000100",
			6585 => "11111110011100010110011101010001",
			6586 => "00000001011000000110011101010001",
			6587 => "0000000101000000000011011100000100",
			6588 => "11111101111010100110011101010001",
			6589 => "00000000001110100110011101010001",
			6590 => "0000000111000000001001110000001000",
			6591 => "0000001000000000001001101000000100",
			6592 => "00000000000110000110011101010001",
			6593 => "00000001011110010110011101010001",
			6594 => "0000000011000000000111001000000100",
			6595 => "11111101000001100110011101010001",
			6596 => "00000000100100000110011101010001",
			6597 => "0000001001000000001101101000010000",
			6598 => "0000000100000000001111100000001000",
			6599 => "0000001000000000000010101000000100",
			6600 => "11111111101011110110011101010001",
			6601 => "11111101111000100110011101010001",
			6602 => "0000001001000000000110101000000100",
			6603 => "11111111111001100110011101010001",
			6604 => "00000000111000110110011101010001",
			6605 => "0000000101000000001010111100001000",
			6606 => "0000000100000000000011001100000100",
			6607 => "11111111100111000110011101010001",
			6608 => "00000000111100110110011101010001",
			6609 => "0000000001000000000010001100000100",
			6610 => "11111111010110000110011101010001",
			6611 => "00000000001001010110011101010001",
			6612 => "0000001110000000001000000010011000",
			6613 => "0000001001000000001111001101011000",
			6614 => "0000001011000000000101101100111100",
			6615 => "0000001110000000000100001000100000",
			6616 => "0000001001000000001011101000010000",
			6617 => "0000001011000000000101101100001000",
			6618 => "0000001001000000000111100100000100",
			6619 => "11111111111110100110100101011101",
			6620 => "00000000001110110110100101011101",
			6621 => "0000000110000000001100011000000100",
			6622 => "00000001100010100110100101011101",
			6623 => "11111101010101110110100101011101",
			6624 => "0000000100000000000011110000001000",
			6625 => "0000000001000000000010001100000100",
			6626 => "00000000011100100110100101011101",
			6627 => "11111110000101110110100101011101",
			6628 => "0000001111000000001101000100000100",
			6629 => "00000010000101100110100101011101",
			6630 => "11111110010010000110100101011101",
			6631 => "0000001111000000001101000100010000",
			6632 => "0000000111000000001000111000001000",
			6633 => "0000000000000000000010011000000100",
			6634 => "11111111100011000110100101011101",
			6635 => "11111110010001110110100101011101",
			6636 => "0000001011000000001101100000000100",
			6637 => "11111111111010100110100101011101",
			6638 => "00000001100111100110100101011101",
			6639 => "0000001110000000000100001000000100",
			6640 => "00000001110111000110100101011101",
			6641 => "0000000000000000000000111000000100",
			6642 => "00000000101110010110100101011101",
			6643 => "11111111101001000110100101011101",
			6644 => "0000000100000000000100001100001100",
			6645 => "0000000110000000001100011000001000",
			6646 => "0000001101000000000100011000000100",
			6647 => "00000000110100000110100101011101",
			6648 => "11111111010000110110100101011101",
			6649 => "11111100111100110110100101011101",
			6650 => "0000000100000000000011101100000100",
			6651 => "00000001010001010110100101011101",
			6652 => "0000001100000000001000111000000100",
			6653 => "11111101111111010110100101011101",
			6654 => "0000000001000000001100110100000100",
			6655 => "11111111001010000110100101011101",
			6656 => "00000001000110110110100101011101",
			6657 => "0000000000000000000000110000110000",
			6658 => "0000000111000000001000111000010100",
			6659 => "0000001011000000000011011100001000",
			6660 => "0000000011000000001001001000000100",
			6661 => "00000000111010110110100101011101",
			6662 => "11111110110101100110100101011101",
			6663 => "0000000001000000001001111000000100",
			6664 => "00000011000000010110100101011101",
			6665 => "0000000001000000001001111000000100",
			6666 => "00000000000000000110100101011101",
			6667 => "00000010011100110110100101011101",
			6668 => "0000001000000000001011010100010000",
			6669 => "0000000010000000001001010000001000",
			6670 => "0000001110000000000100011000000100",
			6671 => "00000001100100010110100101011101",
			6672 => "00000000000000000110100101011101",
			6673 => "0000001101000000000011100000000100",
			6674 => "11111101110011010110100101011101",
			6675 => "11111111001110100110100101011101",
			6676 => "0000000100000000001010110100001000",
			6677 => "0000000110000000001101011000000100",
			6678 => "00000001100111010110100101011101",
			6679 => "11111111100101100110100101011101",
			6680 => "11111110001110010110100101011101",
			6681 => "0000001101000000000110100100001100",
			6682 => "0000000110000000001001100100000100",
			6683 => "00000001110001110110100101011101",
			6684 => "0000000110000000001111000000000100",
			6685 => "00000000000010100110100101011101",
			6686 => "11111111011010010110100101011101",
			6687 => "11111110011100010110100101011101",
			6688 => "0000001111000000001110110100111100",
			6689 => "0000001100000000001000111100100000",
			6690 => "0000001011000000001000111000000100",
			6691 => "00000001010010110110100101011101",
			6692 => "0000000010000000001100010100001100",
			6693 => "0000000110000000001010011000001000",
			6694 => "0000001111000000001101000100000100",
			6695 => "11111111100110110110100101011101",
			6696 => "11111110000011000110100101011101",
			6697 => "00000001101000110110100101011101",
			6698 => "0000000111000000001001110000001000",
			6699 => "0000001100000000000000101000000100",
			6700 => "11111111010100110110100101011101",
			6701 => "11111101111111010110100101011101",
			6702 => "0000001001000000001001011000000100",
			6703 => "00000000011110110110100101011101",
			6704 => "11111110101000010110100101011101",
			6705 => "0000000011000000001010011100000100",
			6706 => "00000010000010100110100101011101",
			6707 => "0000001100000000001000111100001000",
			6708 => "0000001101000000000110100100000100",
			6709 => "00000001100000000110100101011101",
			6710 => "11111110111011000110100101011101",
			6711 => "0000001100000000001000111000001000",
			6712 => "0000001111000000001110010000000100",
			6713 => "11111101101100000110100101011101",
			6714 => "00000000000000000110100101011101",
			6715 => "0000000001000000001001111000000100",
			6716 => "00000001000000100110100101011101",
			6717 => "11111111100011100110100101011101",
			6718 => "0000000011000000001100010100010100",
			6719 => "0000001001000000001100011000001100",
			6720 => "0000000110000000001000010000000100",
			6721 => "00000001111100110110100101011101",
			6722 => "0000001001000000001110010100000100",
			6723 => "00000000000000000110100101011101",
			6724 => "00000001010100000110100101011101",
			6725 => "0000000111000000000011100000000100",
			6726 => "11111110110000100110100101011101",
			6727 => "00000000101010100110100101011101",
			6728 => "0000000100000000000011001100000100",
			6729 => "11111110011110010110100101011101",
			6730 => "0000000001000000000101011100001100",
			6731 => "0000001000000000001000110000000100",
			6732 => "11111110011001000110100101011101",
			6733 => "0000000000000000001000111000000100",
			6734 => "00000000000000000110100101011101",
			6735 => "11111111100100000110100101011101",
			6736 => "0000001000000000000001110100001000",
			6737 => "0000001111000000001011110000000100",
			6738 => "00000001100110110110100101011101",
			6739 => "11111111010100100110100101011101",
			6740 => "0000000010000000001101001000000100",
			6741 => "00000000000000000110100101011101",
			6742 => "00000001100000110110100101011101",
			6743 => "0000000100000000000000101110111000",
			6744 => "0000000101000000000100011001100100",
			6745 => "0000001001000000001111001100111100",
			6746 => "0000000011000000001011000000100000",
			6747 => "0000001001000000001101101000010000",
			6748 => "0000001110000000000110000100001000",
			6749 => "0000001001000000001101101000000100",
			6750 => "00000000000001110110101101000001",
			6751 => "00000000101010010110101101000001",
			6752 => "0000000010000000001001100000000100",
			6753 => "11111110110001000110101101000001",
			6754 => "00000000010010000110101101000001",
			6755 => "0000001110000000001101111000001000",
			6756 => "0000001011000000001001110000000100",
			6757 => "00000000001111010110101101000001",
			6758 => "00000000111100110110101101000001",
			6759 => "0000000110000000000100110100000100",
			6760 => "00000001000001110110101101000001",
			6761 => "11111111111001010110101101000001",
			6762 => "0000000110000000001010011000010000",
			6763 => "0000000101000000000100001000001000",
			6764 => "0000001011000000001001110000000100",
			6765 => "00000001001010100110101101000001",
			6766 => "00000011100000110110101101000001",
			6767 => "0000000111000000001000111000000100",
			6768 => "11111110110001100110101101000001",
			6769 => "00000000010000010110101101000001",
			6770 => "0000000001000000000010001100000100",
			6771 => "00000001010001010110101101000001",
			6772 => "0000001100000000001000111000000100",
			6773 => "11111110101011000110101101000001",
			6774 => "00000000011110000110101101000001",
			6775 => "0000001110000000000100011000010100",
			6776 => "0000001100000000001100001000000100",
			6777 => "00000100001001100110101101000001",
			6778 => "0000001000000000001001101000001000",
			6779 => "0000001011000000000101101100000100",
			6780 => "11111110011101000110101101000001",
			6781 => "00000010100000010110101101000001",
			6782 => "0000001100000000001000111000000100",
			6783 => "00000010010011100110101101000001",
			6784 => "00000000011110100110101101000001",
			6785 => "0000001100000000000000101000000100",
			6786 => "00000010101100000110101101000001",
			6787 => "0000001100000000001000111100001000",
			6788 => "0000000100000000001001001100000100",
			6789 => "11111110110110110110101101000001",
			6790 => "00000001000011010110101101000001",
			6791 => "0000000111000000001001110000000100",
			6792 => "11111111010000100110101101000001",
			6793 => "00000001101010000110101101000001",
			6794 => "0000001000000000001001101000011000",
			6795 => "0000001001000000000100110100010100",
			6796 => "0000001011000000001100101100000100",
			6797 => "11111101101101010110101101000001",
			6798 => "0000001110000000000001101000001000",
			6799 => "0000000100000000000110111000000100",
			6800 => "00000000001110010110101101000001",
			6801 => "11111101111110110110101101000001",
			6802 => "0000001010000000000110011000000100",
			6803 => "00000000011111100110101101000001",
			6804 => "11111110010010110110101101000001",
			6805 => "11111110011001110110101101000001",
			6806 => "0000001100000000001100110000100000",
			6807 => "0000000100000000001000001000010000",
			6808 => "0000001011000000001110001100001000",
			6809 => "0000000010000000000111011000000100",
			6810 => "11111110011000010110101101000001",
			6811 => "00000000101001100110101101000001",
			6812 => "0000000001000000001101101000000100",
			6813 => "00000001010001100110101101000001",
			6814 => "11111111001011100110101101000001",
			6815 => "0000001110000000001001001000001000",
			6816 => "0000001011000000001110001100000100",
			6817 => "11111111110110110110101101000001",
			6818 => "11111100110101010110101101000001",
			6819 => "0000001111000000000100101000000100",
			6820 => "00000001010110110110101101000001",
			6821 => "11111111000000010110101101000001",
			6822 => "0000000100000000001110111000010000",
			6823 => "0000000110000000000101010000001000",
			6824 => "0000000100000000001101001000000100",
			6825 => "00000001010011110110101101000001",
			6826 => "00000011000110100110101101000001",
			6827 => "0000001011000000000110100000000100",
			6828 => "11111110101010000110101101000001",
			6829 => "00000001110001100110101101000001",
			6830 => "0000001000000000001111001000000100",
			6831 => "11111110011111000110101101000001",
			6832 => "0000001100000000000110000100000100",
			6833 => "11111111011000010110101101000001",
			6834 => "00000000110110010110101101000001",
			6835 => "0000001000000000001101010000011100",
			6836 => "0000000001000000000110000000001100",
			6837 => "0000000100000000000110110000001000",
			6838 => "0000001001000000001110100000000100",
			6839 => "11111111011101000110101101000001",
			6840 => "00000001100010000110101101000001",
			6841 => "11111110101000110110101101000001",
			6842 => "0000001111000000001001010100000100",
			6843 => "11111011101011000110101101000001",
			6844 => "0000000110000000001011001100001000",
			6845 => "0000001010000000000101000100000100",
			6846 => "11111111010110000110101101000001",
			6847 => "00000000111010000110101101000001",
			6848 => "11111110010111110110101101000001",
			6849 => "0000000100000000000101100000011100",
			6850 => "0000001100000000000111111000001000",
			6851 => "0000001100000000000111111000000100",
			6852 => "00000001001110100110101101000001",
			6853 => "11111110010111100110101101000001",
			6854 => "0000001011000000000000101000000100",
			6855 => "00000001100111000110101101000001",
			6856 => "0000000010000000000010010100001000",
			6857 => "0000000010000000001100010000000100",
			6858 => "00000000000000000110101101000001",
			6859 => "11111110010001100110101101000001",
			6860 => "0000000100000000000011111000000100",
			6861 => "00000001101011000110101101000001",
			6862 => "11111111010010110110101101000001",
			6863 => "11111110100011110110101101000001",
			6864 => "0000001000000000001011010110001000",
			6865 => "0000000000000000000011010001010100",
			6866 => "0000000110000000001010011000111000",
			6867 => "0000000001000000001001111000011100",
			6868 => "0000000110000000000100110100010000",
			6869 => "0000001011000000000011011100001000",
			6870 => "0000000001000000000010001100000100",
			6871 => "00000000000101100110110101111101",
			6872 => "11111111100011010110110101111101",
			6873 => "0000000001000000000010001100000100",
			6874 => "00000001110100100110110101111101",
			6875 => "11111111110010100110110101111101",
			6876 => "0000000000000000001101010000000100",
			6877 => "00000011110100000110110101111101",
			6878 => "0000000000000000000011111100000100",
			6879 => "00000000100111000110110101111101",
			6880 => "11111110000100110110110101111101",
			6881 => "0000000110000000000100110100010000",
			6882 => "0000000001000000001001111000001000",
			6883 => "0000000101000000001010111100000100",
			6884 => "11111101110110000110110101111101",
			6885 => "11111111111001100110110101111101",
			6886 => "0000001011000000000101101100000100",
			6887 => "00000010010001100110110101111101",
			6888 => "11111111101010110110110101111101",
			6889 => "0000000100000000000011110000001000",
			6890 => "0000000111000000001101100000000100",
			6891 => "11111110011011000110110101111101",
			6892 => "00000000000110000110110101111101",
			6893 => "00000000001100110110110101111101",
			6894 => "0000001000000000000001010100000100",
			6895 => "11111110011000100110110101111101",
			6896 => "0000001111000000000110100000001000",
			6897 => "0000000100000000001000000100000100",
			6898 => "00000000111111100110110101111101",
			6899 => "00000010100010100110110101111101",
			6900 => "0000001000000000000001010100001000",
			6901 => "0000000000000000001000101100000100",
			6902 => "00000000000000000110110101111101",
			6903 => "00000111110000110110110101111101",
			6904 => "0000001110000000001000000000000100",
			6905 => "11111110111100100110110101111101",
			6906 => "00000000100011010110110101111101",
			6907 => "0000000111000000000111111000010100",
			6908 => "0000000011000000001100001000001000",
			6909 => "0000001000000000001001101000000100",
			6910 => "00000000000000000110110101111101",
			6911 => "00000001001100100110110101111101",
			6912 => "0000000101000000001001110000001000",
			6913 => "0000001100000000000000111000000100",
			6914 => "00000000000000000110110101111101",
			6915 => "00000000111000010110110101111101",
			6916 => "11111101010011000110110101111101",
			6917 => "0000000010000000001111010000010000",
			6918 => "0000001000000000001001101000001000",
			6919 => "0000000101000000001101100000000100",
			6920 => "00000001100100110110110101111101",
			6921 => "11111111001101110110110101111101",
			6922 => "0000001111000000000001011000000100",
			6923 => "00000001111001100110110101111101",
			6924 => "00000010110110110110110101111101",
			6925 => "0000000001000000001100110100001100",
			6926 => "0000001000000000001001101000000100",
			6927 => "00000010000110110110110101111101",
			6928 => "0000000111000000001100001000000100",
			6929 => "11111111011101010110110101111101",
			6930 => "00000000110000110110110101111101",
			6931 => "11111101111110010110110101111101",
			6932 => "0000000011000000001011000101001100",
			6933 => "0000000100000000000100001100100000",
			6934 => "0000001010000000001010110000010100",
			6935 => "0000001111000000001011000000001000",
			6936 => "0000001110000000001010101100000100",
			6937 => "00000001011110000110110101111101",
			6938 => "11111110011110000110110101111101",
			6939 => "0000000101000000001000111100000100",
			6940 => "00000000000001110110110101111101",
			6941 => "0000001010000000000110011000000100",
			6942 => "00000000000000000110110101111101",
			6943 => "00000001011110010110110101111101",
			6944 => "0000001110000000001111000100001000",
			6945 => "0000000101000000001001110000000100",
			6946 => "00000001010000100110110101111101",
			6947 => "11111101011101110110110101111101",
			6948 => "00000001100111010110110101111101",
			6949 => "0000000000000000000100010100001100",
			6950 => "0000001011000000000100010100001000",
			6951 => "0000000011000000001110111100000100",
			6952 => "00000000011110010110110101111101",
			6953 => "11111100110100100110110101111101",
			6954 => "00000000001011110110110101111101",
			6955 => "0000000001000000000110000000010000",
			6956 => "0000001111000000001110110000001000",
			6957 => "0000000100000000000110110000000100",
			6958 => "00000001100110000110110101111101",
			6959 => "11111111000101110110110101111101",
			6960 => "0000001111000000000000011100000100",
			6961 => "11111110100100110110110101111101",
			6962 => "00000001100101010110110101111101",
			6963 => "0000000100000000000000100000001000",
			6964 => "0000000101000000001001110000000100",
			6965 => "00000001110001110110110101111101",
			6966 => "00000000010010000110110101111101",
			6967 => "0000001000000000001101010000000100",
			6968 => "11111110100110100110110101111101",
			6969 => "00000000011110110110110101111101",
			6970 => "0000001111000000001000011000001100",
			6971 => "0000001100000000001011000100001000",
			6972 => "0000001100000000000111111000000100",
			6973 => "11111110111011110110110101111101",
			6974 => "11111101100010010110110101111101",
			6975 => "00000000101011010110110101111101",
			6976 => "0000000011000000001100001000100000",
			6977 => "0000000001000000000110000000010000",
			6978 => "0000000101000000000011011100001000",
			6979 => "0000000101000000001000111100000100",
			6980 => "00000000100001000110110101111101",
			6981 => "11111110001110010110110101111101",
			6982 => "0000001011000000001011000000000100",
			6983 => "00000001000010010110110101111101",
			6984 => "00000000000000000110110101111101",
			6985 => "0000000010000000000111100000001000",
			6986 => "0000001100000000000111111000000100",
			6987 => "00000000001011000110110101111101",
			6988 => "00000001111001010110110101111101",
			6989 => "0000000001000000000110000000000100",
			6990 => "00000001010001100110110101111101",
			6991 => "11111111001000110110110101111101",
			6992 => "0000001111000000000110110100010000",
			6993 => "0000001110000000000111111000001000",
			6994 => "0000000000000000000011010000000100",
			6995 => "11111101111110110110110101111101",
			6996 => "11111111111001100110110101111101",
			6997 => "0000001100000000000000101000000100",
			6998 => "11111110110111000110110101111101",
			6999 => "00000000110010110110110101111101",
			7000 => "0000001110000000001100001000001000",
			7001 => "0000000111000000001011000100000100",
			7002 => "11111111111010110110110101111101",
			7003 => "00000000101000010110110101111101",
			7004 => "0000001111000000001011110100000100",
			7005 => "11111111010001000110110101111101",
			7006 => "11111111111010100110110101111101",
			7007 => "0000000101000000001010111110101100",
			7008 => "0000001100000000000000101001001100",
			7009 => "0000001100000000000100010100110000",
			7010 => "0000001001000000001011101000100000",
			7011 => "0000000111000000000100000000010000",
			7012 => "0000000111000000001100001000001000",
			7013 => "0000000111000000000000101000000100",
			7014 => "00000000000100110110111110110001",
			7015 => "11111111101011100110111110110001",
			7016 => "0000001100000000000100010100000100",
			7017 => "00000000010000010110111110110001",
			7018 => "00000001101010110110111110110001",
			7019 => "0000000101000000000100001000001000",
			7020 => "0000000110000000000100110100000100",
			7021 => "11111111111010110110111110110001",
			7022 => "11111110111000110110111110110001",
			7023 => "0000000000000000000000110000000100",
			7024 => "00000010001000000110111110110001",
			7025 => "00000000000000000110111110110001",
			7026 => "0000000110000000000100110100000100",
			7027 => "11111110100100010110111110110001",
			7028 => "0000001110000000001010111100000100",
			7029 => "00000010101010010110111110110001",
			7030 => "0000001101000000001010111100000100",
			7031 => "11111111010000010110111110110001",
			7032 => "00000001111000110110111110110001",
			7033 => "0000000111000000000000101000001100",
			7034 => "0000000010000000000111100000000100",
			7035 => "00000000000000000110111110110001",
			7036 => "0000000100000000001001001100000100",
			7037 => "11111110001110000110111110110001",
			7038 => "11111101000111010110111110110001",
			7039 => "0000001110000000001100101100001100",
			7040 => "0000001111000000001010010100001000",
			7041 => "0000000001000000001100110100000100",
			7042 => "00000000000001010110111110110001",
			7043 => "11111101111011110110111110110001",
			7044 => "00000001111011000110111110110001",
			7045 => "11111110000011010110111110110001",
			7046 => "0000001100000000000000101000101000",
			7047 => "0000000111000000000100010100001000",
			7048 => "0000000100000000000101010100000100",
			7049 => "11111101101110100110111110110001",
			7050 => "11111111100111100110111110110001",
			7051 => "0000001011000000000100000000010000",
			7052 => "0000001011000000001100001000001000",
			7053 => "0000000111000000001011000100000100",
			7054 => "00000001101100100110111110110001",
			7055 => "00000000010110100110111110110001",
			7056 => "0000000010000000000011001000000100",
			7057 => "00000001111101010110111110110001",
			7058 => "00000000010001110110111110110001",
			7059 => "0000001010000000001001000100001000",
			7060 => "0000000100000000001000110100000100",
			7061 => "00000000000101010110111110110001",
			7062 => "00000001000001100110111110110001",
			7063 => "0000000010000000001110010000000100",
			7064 => "11111111100100100110111110110001",
			7065 => "00000000011101100110111110110001",
			7066 => "0000001100000000000000101000011000",
			7067 => "0000001011000000001100001000001000",
			7068 => "0000000101000000001100101100000100",
			7069 => "11111111001000010110111110110001",
			7070 => "00000010101110000110111110110001",
			7071 => "0000000101000000001100101000001000",
			7072 => "0000000000000000000111111000000100",
			7073 => "11111101100111110110111110110001",
			7074 => "11111111000011010110111110110001",
			7075 => "0000000111000000000100000000000100",
			7076 => "00000001000111110110111110110001",
			7077 => "11111110010000110110111110110001",
			7078 => "0000001100000000000100000000010000",
			7079 => "0000000111000000000100000000001000",
			7080 => "0000000100000000000110001100000100",
			7081 => "11111110000001110110111110110001",
			7082 => "00000000001010010110111110110001",
			7083 => "0000001001000000001011101000000100",
			7084 => "00000010000010010110111110110001",
			7085 => "00000000000000000110111110110001",
			7086 => "0000000110000000001100011000001000",
			7087 => "0000001111000000000010001000000100",
			7088 => "00000000011111010110111110110001",
			7089 => "11111111001001100110111110110001",
			7090 => "0000001010000000000110011000000100",
			7091 => "00000001110110100110111110110001",
			7092 => "00000000000011000110111110110001",
			7093 => "0000000111000000001000111000100000",
			7094 => "0000001100000000001000111100011100",
			7095 => "0000000100000000001110100100001000",
			7096 => "0000000000000000000111000000000100",
			7097 => "11111111011100000110111110110001",
			7098 => "11111101101111010110111110110001",
			7099 => "0000001011000000001101100000001000",
			7100 => "0000001001000000001111001100000100",
			7101 => "00000001100011100110111110110001",
			7102 => "11111111011000110110111110110001",
			7103 => "0000001001000000001101011100001000",
			7104 => "0000001001000000001011101000000100",
			7105 => "11111101000111010110111110110001",
			7106 => "11111110001101010110111110110001",
			7107 => "00000000001101000110111110110001",
			7108 => "00000000101011000110111110110001",
			7109 => "0000001111000000000001000000100000",
			7110 => "0000001101000000001101010100000100",
			7111 => "11111110010000000110111110110001",
			7112 => "0000000100000000001111100000001100",
			7113 => "0000001111000000000001000000001000",
			7114 => "0000000100000000001001001100000100",
			7115 => "00000000001000010110111110110001",
			7116 => "00000001000111010110111110110001",
			7117 => "00000010000110110110111110110001",
			7118 => "0000001001000000001011101000001000",
			7119 => "0000000110000000001101011000000100",
			7120 => "11111110000000000110111110110001",
			7121 => "00000001001101010110111110110001",
			7122 => "0000000110000000001011001100000100",
			7123 => "11111001010101100110111110110001",
			7124 => "11111111001011000110111110110001",
			7125 => "0000001110000000000100011000010100",
			7126 => "0000000110000000001011001100001100",
			7127 => "0000001001000000001101011100001000",
			7128 => "0000001011000000000110000100000100",
			7129 => "11111101001010000110111110110001",
			7130 => "11111111100111010110111110110001",
			7131 => "00000001000011010110111110110001",
			7132 => "0000000110000000001001100100000100",
			7133 => "00000001011110010110111110110001",
			7134 => "00000000000000000110111110110001",
			7135 => "0000000010000000000110010000001100",
			7136 => "0000001101000000001011000000000100",
			7137 => "11111111110111010110111110110001",
			7138 => "0000000110000000001011001100000100",
			7139 => "11111110001010100110111110110001",
			7140 => "11111111111011110110111110110001",
			7141 => "0000000110000000001010011000001000",
			7142 => "0000001100000000001000111100000100",
			7143 => "00000001110101010110111110110001",
			7144 => "00000000000110010110111110110001",
			7145 => "0000000111000000001001110000000100",
			7146 => "11111110101110010110111110110001",
			7147 => "00000000000001110110111110110001",
			7148 => "0000001100000000000100000010100000",
			7149 => "0000000111000000001001110001110000",
			7150 => "0000000101000000001010111100111100",
			7151 => "0000001100000000000100000000100000",
			7152 => "0000000011000000000011100000010000",
			7153 => "0000000011000000000100011000001000",
			7154 => "0000001101000000000111001000000100",
			7155 => "00000000000001100111000111100101",
			7156 => "00000001110111100111000111100101",
			7157 => "0000001011000000001001110000000100",
			7158 => "11111111111111010111000111100101",
			7159 => "11111110101011000111000111100101",
			7160 => "0000001100000000000000101000001000",
			7161 => "0000001000000000000111000100000100",
			7162 => "11111110101101100111000111100101",
			7163 => "00000000111000000111000111100101",
			7164 => "0000000111000000001100001000000100",
			7165 => "11111110111000100111000111100101",
			7166 => "00000001001110010111000111100101",
			7167 => "0000000111000000000100000000001100",
			7168 => "0000000111000000000100000000001000",
			7169 => "0000001001000000000111100100000100",
			7170 => "11111111100101100111000111100101",
			7171 => "00000001101110110111000111100101",
			7172 => "11111110010110100111000111100101",
			7173 => "0000001010000000001100011100001000",
			7174 => "0000000111000000001000111000000100",
			7175 => "00000010001101100111000111100101",
			7176 => "00000000100011110111000111100101",
			7177 => "0000000010000000001001100000000100",
			7178 => "00000001011000000111000111100101",
			7179 => "11111111100011010111000111100101",
			7180 => "0000001001000000001101011100100000",
			7181 => "0000001011000000001101100000010000",
			7182 => "0000001100000000000100000000001000",
			7183 => "0000000111000000000100000000000100",
			7184 => "11111110011100110111000111100101",
			7185 => "00000000000000000111000111100101",
			7186 => "0000000111000000001000111000000100",
			7187 => "00000010000101110111000111100101",
			7188 => "11111111000000000111000111100101",
			7189 => "0000000110000000000100110100001000",
			7190 => "0000000100000000001000000100000100",
			7191 => "11111111001010100111000111100101",
			7192 => "00000000111100010111000111100101",
			7193 => "0000000100000000000100001100000100",
			7194 => "11111110010100110111000111100101",
			7195 => "11111111111110100111000111100101",
			7196 => "0000001100000000000000101000000100",
			7197 => "00000010000011110111000111100101",
			7198 => "0000001110000000001000000000001000",
			7199 => "0000000010000000000010000000000100",
			7200 => "11111111111100000111000111100101",
			7201 => "00000010000000110111000111100101",
			7202 => "0000000010000000001110110100000100",
			7203 => "11111110100101100111000111100101",
			7204 => "00000000101111100111000111100101",
			7205 => "0000001000000000000001110100101000",
			7206 => "0000000101000000001010111000001100",
			7207 => "0000000010000000000101110000000100",
			7208 => "11111111011001100111000111100101",
			7209 => "0000001000000000000111000100000100",
			7210 => "00000010000111100111000111100101",
			7211 => "00000000111100000111000111100101",
			7212 => "0000001101000000000110100100010000",
			7213 => "0000000110000000001101011000001000",
			7214 => "0000000010000000001100010100000100",
			7215 => "11111111001101110111000111100101",
			7216 => "00000001111001010111000111100101",
			7217 => "0000000100000000001110100100000100",
			7218 => "00000000101011000111000111100101",
			7219 => "11111110001000100111000111100101",
			7220 => "0000001001000000001011111100001000",
			7221 => "0000000010000000001100010000000100",
			7222 => "00000000110001100111000111100101",
			7223 => "00000010000011000111000111100101",
			7224 => "11111111110011000111000111100101",
			7225 => "0000001000000000000010101000000100",
			7226 => "11111101110001000111000111100101",
			7227 => "00000000100111110111000111100101",
			7228 => "0000001100000000000100000000011100",
			7229 => "0000000101000000001010111000010100",
			7230 => "0000001011000000001000111000000100",
			7231 => "00000000001100110111000111100101",
			7232 => "0000001010000000001100011100001100",
			7233 => "0000000001000000001001111000001000",
			7234 => "0000000010000000000100101000000100",
			7235 => "11111111001010110111000111100101",
			7236 => "11111101101110100111000111100101",
			7237 => "11111111100111110111000111100101",
			7238 => "11111111100101100111000111100101",
			7239 => "0000001110000000001000011000000100",
			7240 => "00000001110011110111000111100101",
			7241 => "11111110111110010111000111100101",
			7242 => "0000001100000000001000111100101000",
			7243 => "0000001100000000001000111100011000",
			7244 => "0000000111000000001001110000010000",
			7245 => "0000001110000000001101100000001000",
			7246 => "0000000001000000000010001100000100",
			7247 => "00000000001100000111000111100101",
			7248 => "00000010000101100111000111100101",
			7249 => "0000001110000000001100101100000100",
			7250 => "11111101110010010111000111100101",
			7251 => "00000000010010100111000111100101",
			7252 => "0000001000000000000111000100000100",
			7253 => "11111101110001010111000111100101",
			7254 => "00000000100010110111000111100101",
			7255 => "0000000001000000001001111000000100",
			7256 => "00000010001010010111000111100101",
			7257 => "0000001110000000001001001000000100",
			7258 => "11111111111001110111000111100101",
			7259 => "0000001010000000000001010000000100",
			7260 => "00000001111011100111000111100101",
			7261 => "00000000000000000111000111100101",
			7262 => "0000000110000000001010011000011100",
			7263 => "0000000100000000000000010100001100",
			7264 => "0000001000000000001111001000001000",
			7265 => "0000001101000000001110110000000100",
			7266 => "00000000000000000111000111100101",
			7267 => "11111110011001010111000111100101",
			7268 => "11111101101010100111000111100101",
			7269 => "0000001101000000001011000000001000",
			7270 => "0000000001000000001110100000000100",
			7271 => "00000000000000000111000111100101",
			7272 => "00000001101100000111000111100101",
			7273 => "0000000110000000001010011000000100",
			7274 => "11111111011000000111000111100101",
			7275 => "00000000000000000111000111100101",
			7276 => "0000000010000000000100101000001100",
			7277 => "0000001101000000001001001000001000",
			7278 => "0000001011000000000000001100000100",
			7279 => "00000001110101010111000111100101",
			7280 => "00000000000000000111000111100101",
			7281 => "00000000000000000111000111100101",
			7282 => "0000001001000000001101101000001000",
			7283 => "0000000100000000001101001100000100",
			7284 => "00000001100101010111000111100101",
			7285 => "00000000000000000111000111100101",
			7286 => "0000001101000000001010111000000100",
			7287 => "11111111000000110111000111100101",
			7288 => "11111111111110110111000111100101",
			7289 => "0000001001000000001001111001111000",
			7290 => "0000001100000000000100010100111100",
			7291 => "0000001100000000000100010100111000",
			7292 => "0000000100000000000001101100011100",
			7293 => "0000001110000000001111000100001100",
			7294 => "0000001011000000000100010100001000",
			7295 => "0000001111000000000111010000000100",
			7296 => "11111111111110110111010001000001",
			7297 => "00000001110111110111010001000001",
			7298 => "00000001101001000111010001000001",
			7299 => "0000001111000000000000011100001000",
			7300 => "0000000000000000001110111100000100",
			7301 => "11111111101000000111010001000001",
			7302 => "11111110101000100111010001000001",
			7303 => "0000001100000000000111111000000100",
			7304 => "00000000000111010111010001000001",
			7305 => "11111101101110000111010001000001",
			7306 => "0000001010000000000001010100010000",
			7307 => "0000000011000000000010111100001000",
			7308 => "0000000011000000000010011000000100",
			7309 => "00000000000000000111010001000001",
			7310 => "11110110101100010111010001000001",
			7311 => "0000000000000000001100001000000100",
			7312 => "00000000000000000111010001000001",
			7313 => "11111110000110010111010001000001",
			7314 => "0000001010000000000001110000000100",
			7315 => "00000001101000000111010001000001",
			7316 => "0000001110000000001011010100000100",
			7317 => "11111110110000000111010001000001",
			7318 => "00000000000000000111010001000001",
			7319 => "00000001101110010111010001000001",
			7320 => "0000000011000000000100000000101100",
			7321 => "0000000001000000000110000000010100",
			7322 => "0000001111000000000101100100001100",
			7323 => "0000000001000000000000011000001000",
			7324 => "0000001110000000000010101000000100",
			7325 => "11111111101000100111010001000001",
			7326 => "00000000000001000111010001000001",
			7327 => "00000001101111100111010001000001",
			7328 => "0000001111000000001011011100000100",
			7329 => "11111110110111000111010001000001",
			7330 => "00000000100001110111010001000001",
			7331 => "0000001101000000001100110000010000",
			7332 => "0000001001000000000010001100001000",
			7333 => "0000001101000000001101100000000100",
			7334 => "11111110101110110111010001000001",
			7335 => "11111100110010000111010001000001",
			7336 => "0000001011000000000100010100000100",
			7337 => "11111110110010100111010001000001",
			7338 => "00000001011100110111010001000001",
			7339 => "0000000101000000001100110000000100",
			7340 => "00000001110011000111010001000001",
			7341 => "11111110001000000111010001000001",
			7342 => "0000001100000000000100010100000100",
			7343 => "11111100110011000111010001000001",
			7344 => "0000001110000000001110111100001000",
			7345 => "0000001111000000000110110100000100",
			7346 => "00000000000000000111010001000001",
			7347 => "00000001001000110111010001000001",
			7348 => "11111110001001110111010001000001",
			7349 => "0000000011000000000101101101001000",
			7350 => "0000000011000000000101101100110100",
			7351 => "0000000011000000001100110000100000",
			7352 => "0000001001000000000111100100010000",
			7353 => "0000000001000000001100110100001000",
			7354 => "0000000111000000000111111000000100",
			7355 => "11111111011001110111010001000001",
			7356 => "00000000001110000111010001000001",
			7357 => "0000000111000000000000101000000100",
			7358 => "00000000101011000111010001000001",
			7359 => "11111110111111100111010001000001",
			7360 => "0000000001000000001100110100001000",
			7361 => "0000000101000000001101111000000100",
			7362 => "00000001110001110111010001000001",
			7363 => "11111111011000010111010001000001",
			7364 => "0000001001000000000111100100000100",
			7365 => "11111111001111100111010001000001",
			7366 => "00000001110110110111010001000001",
			7367 => "0000000110000000000100110100001100",
			7368 => "0000001100000000000100010100001000",
			7369 => "0000001100000000000100010100000100",
			7370 => "11111111100110110111010001000001",
			7371 => "00000001100101010111010001000001",
			7372 => "11111110100001000111010001000001",
			7373 => "0000001111000000001011110100000100",
			7374 => "11111101110110000111010001000001",
			7375 => "11111110111000010111010001000001",
			7376 => "0000001011000000001100001000001100",
			7377 => "0000000111000000001011000100000100",
			7378 => "00000001000010100111010001000001",
			7379 => "0000001110000000001011000100000100",
			7380 => "00000001001100000111010001000001",
			7381 => "00000010011111110111010001000001",
			7382 => "0000001101000000001110001100000100",
			7383 => "11111111110111000111010001000001",
			7384 => "00000001011111010111010001000001",
			7385 => "0000001001000000000110101000110000",
			7386 => "0000001111000000000101110100010100",
			7387 => "0000001111000000001011011100001000",
			7388 => "0000000100000000001000011100000100",
			7389 => "11111110101001100111010001000001",
			7390 => "00000000011111000111010001000001",
			7391 => "0000000111000000001100001000001000",
			7392 => "0000001010000000000001010000000100",
			7393 => "11111110010010010111010001000001",
			7394 => "11111111010100000111010001000001",
			7395 => "11111101010011110111010001000001",
			7396 => "0000000101000000001100101100010000",
			7397 => "0000001100000000000111111000001000",
			7398 => "0000000011000000001100101100000100",
			7399 => "11111101100100000111010001000001",
			7400 => "11111111100011110111010001000001",
			7401 => "0000001100000000000100010100000100",
			7402 => "00000000010000010111010001000001",
			7403 => "11111110101000000111010001000001",
			7404 => "0000001001000000000110101000000100",
			7405 => "11111111111001000111010001000001",
			7406 => "0000001110000000001000111000000100",
			7407 => "00000010011010000111010001000001",
			7408 => "00000000101100010111010001000001",
			7409 => "0000001100000000000000101000100000",
			7410 => "0000001100000000000000101000010000",
			7411 => "0000001100000000000000101000001000",
			7412 => "0000001001000000001111001100000100",
			7413 => "11111111110011000111010001000001",
			7414 => "00000001101000010111010001000001",
			7415 => "0000000111000000000100000000000100",
			7416 => "00000001000011000111010001000001",
			7417 => "11111111111010000111010001000001",
			7418 => "0000001101000000000001111100001000",
			7419 => "0000000111000000000100000000000100",
			7420 => "11111111000110100111010001000001",
			7421 => "00000000011110000111010001000001",
			7422 => "0000000111000000001000111000000100",
			7423 => "11111101111110010111010001000001",
			7424 => "11111111011110110111010001000001",
			7425 => "0000000111000000001100001000010000",
			7426 => "0000000111000000001100001000001000",
			7427 => "0000001011000000001100001000000100",
			7428 => "00000010001110110111010001000001",
			7429 => "11111111110100110111010001000001",
			7430 => "0000001100000000000000101000000100",
			7431 => "00000001010110100111010001000001",
			7432 => "00000000011000010111010001000001",
			7433 => "0000001001000000001101101000001000",
			7434 => "0000000001000000001100110100000100",
			7435 => "00000000011000000111010001000001",
			7436 => "11111111010001100111010001000001",
			7437 => "0000000001000000001100110100000100",
			7438 => "00000010011100100111010001000001",
			7439 => "00000000000011000111010001000001",
			7440 => "0000001100000000000111111011000000",
			7441 => "0000001001000000000110101001101100",
			7442 => "0000000011000000001001110000111100",
			7443 => "0000001001000000001001111000100000",
			7444 => "0000000001000000001110100000010000",
			7445 => "0000000110000000000111101000001000",
			7446 => "0000001011000000000100010100000100",
			7447 => "11111110000000110111011011000101",
			7448 => "00000000111100110111011011000101",
			7449 => "0000000001000000000110000000000100",
			7450 => "11111111101001000111011011000101",
			7451 => "00000000010111100111011011000101",
			7452 => "0000001011000000000100010100001000",
			7453 => "0000000101000000000011011100000100",
			7454 => "11111101100111000111011011000101",
			7455 => "11111111110110010111011011000101",
			7456 => "0000000111000000000100010100000100",
			7457 => "00000001111010000111011011000101",
			7458 => "11111111101011100111011011000101",
			7459 => "0000000100000000000011110000001100",
			7460 => "0000001110000000000000110000001000",
			7461 => "0000000011000000001100001000000100",
			7462 => "00000001110010110111011011000101",
			7463 => "11111111101100000111011011000101",
			7464 => "11111110010110000111011011000101",
			7465 => "0000001010000000000001010000001000",
			7466 => "0000001011000000000100010100000100",
			7467 => "11111111101000110111011011000101",
			7468 => "00000001110110000111011011000101",
			7469 => "0000000000000000000100010100000100",
			7470 => "11111111010110010111011011000101",
			7471 => "00000001100101010111011011000101",
			7472 => "0000000010000000000101110000010100",
			7473 => "0000000110000000001101111100001100",
			7474 => "0000000001000000001110100000000100",
			7475 => "11111101011011100111011011000101",
			7476 => "0000000010000000000101001000000100",
			7477 => "11111110111111110111011011000101",
			7478 => "00000001010010110111011011000101",
			7479 => "0000000111000000000100010100000100",
			7480 => "11111110101001010111011011000101",
			7481 => "11111101101101100111011011000101",
			7482 => "0000001010000000000001010000010000",
			7483 => "0000000011000000000101101100001000",
			7484 => "0000000101000000001101100000000100",
			7485 => "11111111100111100111011011000101",
			7486 => "00000010000001000111011011000101",
			7487 => "0000000100000000001001001100000100",
			7488 => "11111101111111110111011011000101",
			7489 => "00000001110010000111011011000101",
			7490 => "0000001010000000001100011100001000",
			7491 => "0000001100000000000111111000000100",
			7492 => "11111110000100110111011011000101",
			7493 => "11111111011111000111011011000101",
			7494 => "00000001010110000111011011000101",
			7495 => "0000000101000000001100110000011000",
			7496 => "0000001011000000000000101000010000",
			7497 => "0000001100000000000111111000001100",
			7498 => "0000001110000000000000101000001000",
			7499 => "0000000010000000000010011100000100",
			7500 => "00000010011100110111011011000101",
			7501 => "00000001011010100111011011000101",
			7502 => "00000000000100010111011011000101",
			7503 => "11111111000101000111011011000101",
			7504 => "0000001001000000000110101000000100",
			7505 => "00000001011110110111011011000101",
			7506 => "00000011011100100111011011000101",
			7507 => "0000001010000000001001000100100000",
			7508 => "0000000100000000001000110100010000",
			7509 => "0000001010000000001000100100001000",
			7510 => "0000000100000000000010010100000100",
			7511 => "11111111110100000111011011000101",
			7512 => "00000001111010110111011011000101",
			7513 => "0000001100000000000111111000000100",
			7514 => "11111111011100100111011011000101",
			7515 => "11111110001010010111011011000101",
			7516 => "0000000001000000001100110100001000",
			7517 => "0000000011000000000110000100000100",
			7518 => "00000001100110000111011011000101",
			7519 => "11111111000000100111011011000101",
			7520 => "0000000101000000001110001100000100",
			7521 => "00000011010101110111011011000101",
			7522 => "00000000110001110111011011000101",
			7523 => "0000001100000000000111111000001100",
			7524 => "0000000101000000001100101100001000",
			7525 => "0000001000000000000110001000000100",
			7526 => "11111111111101110111011011000101",
			7527 => "11111101110001110111011011000101",
			7528 => "00000001001100100111011011000101",
			7529 => "0000000001000000001100110100001000",
			7530 => "0000001010000000000110011000000100",
			7531 => "11111111001110000111011011000101",
			7532 => "00000001010000010111011011000101",
			7533 => "0000001110000000000000101000000100",
			7534 => "11111101010110010111011011000101",
			7535 => "00000000000111100111011011000101",
			7536 => "0000001100000000000100010100111100",
			7537 => "0000000100000000001000001000010100",
			7538 => "0000000001000000001100110100001100",
			7539 => "0000000111000000000100010100000100",
			7540 => "11111110101000000111011011000101",
			7541 => "0000000111000000000000101000000100",
			7542 => "00000000101010100111011011000101",
			7543 => "00000010011100010111011011000101",
			7544 => "0000001100000000000111111000000100",
			7545 => "00000000010001000111011011000101",
			7546 => "11111101111010010111011011000101",
			7547 => "0000000000000000001011000100011000",
			7548 => "0000001110000000000100010100001100",
			7549 => "0000000010000000000110100000000100",
			7550 => "11111101000101100111011011000101",
			7551 => "0000001000000000000111000100000100",
			7552 => "00000000011101100111011011000101",
			7553 => "11111110000010010111011011000101",
			7554 => "0000000010000000000011001000000100",
			7555 => "11111101011111100111011011000101",
			7556 => "0000001110000000001001110000000100",
			7557 => "00000000110010100111011011000101",
			7558 => "11111110101000010111011011000101",
			7559 => "0000001000000000001010101100000100",
			7560 => "00000001101100100111011011000101",
			7561 => "0000000010000000001100100100001000",
			7562 => "0000001001000000000000011000000100",
			7563 => "00000000000000000111011011000101",
			7564 => "00000001100111000111011011000101",
			7565 => "11111110011111110111011011000101",
			7566 => "0000000101000000001001110000001000",
			7567 => "0000000000000000000110000100000100",
			7568 => "00000001101110000111011011000101",
			7569 => "00000000000000000111011011000101",
			7570 => "0000000111000000001000111000100000",
			7571 => "0000000111000000000100000000010000",
			7572 => "0000000111000000000100000000001000",
			7573 => "0000000111000000001100001000000100",
			7574 => "00000000000100010111011011000101",
			7575 => "11111111100101000111011011000101",
			7576 => "0000000111000000000100000000000100",
			7577 => "00000000101101110111011011000101",
			7578 => "00000010001100100111011011000101",
			7579 => "0000001011000000000011011100001000",
			7580 => "0000000000000000000011111100000100",
			7581 => "11111111111000100111011011000101",
			7582 => "11111110101000110111011011000101",
			7583 => "0000000100000000001001001100000100",
			7584 => "00000000000000110111011011000101",
			7585 => "00000010000100000111011011000101",
			7586 => "0000000011000000001000011000010000",
			7587 => "0000000110000000001100011000001000",
			7588 => "0000001001000000000111100100000100",
			7589 => "11111110010100110111011011000101",
			7590 => "00000000000110010111011011000101",
			7591 => "0000000101000000001000000000000100",
			7592 => "00000000110010100111011011000101",
			7593 => "11111101010010010111011011000101",
			7594 => "0000000111000000001101100000001000",
			7595 => "0000000001000000000110101000000100",
			7596 => "11111111110011100111011011000101",
			7597 => "11111110011100110111011011000101",
			7598 => "0000001110000000001110110000000100",
			7599 => "11111101111100010111011011000101",
			7600 => "00000000001001100111011011000101",
			7601 => "0000001010000000001010110010010000",
			7602 => "0000001000000000000111000101101100",
			7603 => "0000000010000000001110110100111000",
			7604 => "0000001011000000000111111000011000",
			7605 => "0000001011000000001110111100001100",
			7606 => "0000001011000000001110111100001000",
			7607 => "0000001010000000001001000100000100",
			7608 => "11111101011000000111100101010001",
			7609 => "00000000111010110111100101010001",
			7610 => "11111101100100000111100101010001",
			7611 => "0000001000000000000001110000000100",
			7612 => "11111110111000100111100101010001",
			7613 => "0000000010000000000101110000000100",
			7614 => "00000001110100100111100101010001",
			7615 => "00000000010111110111100101010001",
			7616 => "0000001010000000001001000100010000",
			7617 => "0000001000000000001011010100001000",
			7618 => "0000000001000000000110000000000100",
			7619 => "11111110101111000111100101010001",
			7620 => "00000000000010010111100101010001",
			7621 => "0000001001000000001101101000000100",
			7622 => "00000000010101100111100101010001",
			7623 => "00000011000010100111100101010001",
			7624 => "0000000010000000000111111100001000",
			7625 => "0000000000000000000010111100000100",
			7626 => "00000001101011000111100101010001",
			7627 => "11111111101010010111100101010001",
			7628 => "0000001000000000001111001000000100",
			7629 => "11111111111010100111100101010001",
			7630 => "00000000111011100111100101010001",
			7631 => "0000001000000000001001101000010100",
			7632 => "0000001000000000001001101000010000",
			7633 => "0000001011000000000100001000001000",
			7634 => "0000000001000000000010001100000100",
			7635 => "00000000000000000111100101010001",
			7636 => "00000001101011000111100101010001",
			7637 => "0000000100000000001100001100000100",
			7638 => "11111110110100100111100101010001",
			7639 => "00000000010101100111100101010001",
			7640 => "11111101111111010111100101010001",
			7641 => "0000001010000000000110011000010000",
			7642 => "0000001010000000001001000100001000",
			7643 => "0000001000000000001001101000000100",
			7644 => "11111111011000010111100101010001",
			7645 => "00000000000000000111100101010001",
			7646 => "0000001001000000000111101000000100",
			7647 => "00000010100001000111100101010001",
			7648 => "00000000000000000111100101010001",
			7649 => "0000001010000000000001010000001000",
			7650 => "0000000100000000001000001000000100",
			7651 => "00000000001101100111100101010001",
			7652 => "11111110101100010111100101010001",
			7653 => "0000000010000000001100000000000100",
			7654 => "00000000100111100111100101010001",
			7655 => "00000001101100110111100101010001",
			7656 => "0000000100000000000000010100010000",
			7657 => "0000001010000000000001010000001000",
			7658 => "0000001100000000000111111000000100",
			7659 => "00000000010001100111100101010001",
			7660 => "00000010010100000111100101010001",
			7661 => "0000000011000000001000111100000100",
			7662 => "00000010000010010111100101010001",
			7663 => "11111111101001110111100101010001",
			7664 => "0000000000000000001110111100000100",
			7665 => "11111110101011000111100101010001",
			7666 => "0000001001000000001001111000001100",
			7667 => "0000000111000000000100010100001000",
			7668 => "0000001001000000001100110100000100",
			7669 => "11111111101000010111100101010001",
			7670 => "00000001110110010111100101010001",
			7671 => "11111110111010000111100101010001",
			7672 => "00000001111100100111100101010001",
			7673 => "0000000100000000000000010101010000",
			7674 => "0000000000000000000111111000111100",
			7675 => "0000001000000000000111000100100000",
			7676 => "0000001000000000000111000100010000",
			7677 => "0000000100000000001001001100001000",
			7678 => "0000000100000000001010110100000100",
			7679 => "11111111110011000111100101010001",
			7680 => "11111111001010000111100101010001",
			7681 => "0000000111000000001100001000000100",
			7682 => "11111111100000110111100101010001",
			7683 => "00000000110000110111100101010001",
			7684 => "0000000010000000001100010100001000",
			7685 => "0000000111000000001011000100000100",
			7686 => "00000010100010100111100101010001",
			7687 => "11111111101010110111100101010001",
			7688 => "0000000100000000001010110100000100",
			7689 => "11111110111101100111100101010001",
			7690 => "00000010011100100111100101010001",
			7691 => "0000000100000000001010110100001100",
			7692 => "0000001100000000000000101000000100",
			7693 => "11111110111001010111100101010001",
			7694 => "0000000000000000000000110000000100",
			7695 => "00000000000000000111100101010001",
			7696 => "00000010001001000111100101010001",
			7697 => "0000000101000000000101101100001000",
			7698 => "0000001000000000000111000100000100",
			7699 => "00000010000100000111100101010001",
			7700 => "11111111001010110111100101010001",
			7701 => "0000001001000000001011101000000100",
			7702 => "11111110101100110111100101010001",
			7703 => "11111111101010000111100101010001",
			7704 => "0000000001000000001110100000000100",
			7705 => "11111111001010000111100101010001",
			7706 => "0000000100000000000000010100001100",
			7707 => "0000001110000000001110001100001000",
			7708 => "0000001010000000001100011100000100",
			7709 => "00000010011100110111100101010001",
			7710 => "00000001011100110111100101010001",
			7711 => "00000000000000000111100101010001",
			7712 => "00000000000101100111100101010001",
			7713 => "0000001001000000000110101000110000",
			7714 => "0000000001000000001100110100100000",
			7715 => "0000000001000000001110100000010000",
			7716 => "0000000000000000001011000100001000",
			7717 => "0000000100000000001111100000000100",
			7718 => "11111111111101000111100101010001",
			7719 => "11111110110100110111100101010001",
			7720 => "0000000100000000000010100100000100",
			7721 => "00000000101100110111100101010001",
			7722 => "11111111110100010111100101010001",
			7723 => "0000000101000000001100110000001000",
			7724 => "0000000101000000001100110000000100",
			7725 => "00000001100010000111100101010001",
			7726 => "11111110101010100111100101010001",
			7727 => "0000001110000000000000101000000100",
			7728 => "00000001101000100111100101010001",
			7729 => "00000000001110000111100101010001",
			7730 => "0000001011000000001000111100001100",
			7731 => "0000001110000000001000111000001000",
			7732 => "0000001111000000001001010100000100",
			7733 => "11111110100111010111100101010001",
			7734 => "00000001000000000111100101010001",
			7735 => "11111101001110100111100101010001",
			7736 => "00000001010100000111100101010001",
			7737 => "0000001111000000001110101100011100",
			7738 => "0000001111000000000001001000010000",
			7739 => "0000000100000000001011100000001000",
			7740 => "0000001111000000001001010100000100",
			7741 => "00000000100110010111100101010001",
			7742 => "11111110010101110111100101010001",
			7743 => "0000001111000000001010010100000100",
			7744 => "11111101101101000111100101010001",
			7745 => "00000000101011110111100101010001",
			7746 => "0000001010000000001010110000000100",
			7747 => "00000000100001110111100101010001",
			7748 => "0000001010000000000101000100000100",
			7749 => "00000010000101100111100101010001",
			7750 => "00000000011010000111100101010001",
			7751 => "0000000000000000001110111100001100",
			7752 => "0000001011000000000011011100000100",
			7753 => "00000010001101000111100101010001",
			7754 => "0000001100000000001000111000000100",
			7755 => "11111110011110110111100101010001",
			7756 => "00000000011111000111100101010001",
			7757 => "0000000100000000000100001100001000",
			7758 => "0000000111000000000100000000000100",
			7759 => "11111101111011100111100101010001",
			7760 => "11111111011010000111100101010001",
			7761 => "0000001010000000001100011100000100",
			7762 => "00000000110101100111100101010001",
			7763 => "11111111101110010111100101010001",
			7764 => "0000001001000000000110101011000100",
			7765 => "0000000011000000000011011101101100",
			7766 => "0000001111000000000110110101000000",
			7767 => "0000001110000000000011111100100000",
			7768 => "0000000011000000000000101000010000",
			7769 => "0000000001000000001110100000001000",
			7770 => "0000001001000000000010001100000100",
			7771 => "11111111111010110111101111010101",
			7772 => "00000000100111010111101111010101",
			7773 => "0000000110000000000111101000000100",
			7774 => "00000000010110100111101111010101",
			7775 => "11111100111010010111101111010101",
			7776 => "0000001111000000000001011000001000",
			7777 => "0000001010000000001100011100000100",
			7778 => "00000001110111110111101111010101",
			7779 => "00000000001001100111101111010101",
			7780 => "0000000110000000001101111100000100",
			7781 => "11111110001001000111101111010101",
			7782 => "00000001011100010111101111010101",
			7783 => "0000001001000000000010001100010000",
			7784 => "0000000011000000000000101000001000",
			7785 => "0000001000000000000001110100000100",
			7786 => "00000001100111100111101111010101",
			7787 => "11111110111011010111101111010101",
			7788 => "0000001111000000000101100100000100",
			7789 => "11111101011110000111101111010101",
			7790 => "11111111101000000111101111010101",
			7791 => "0000001111000000001010011100001000",
			7792 => "0000000110000000000111101000000100",
			7793 => "00000000111010000111101111010101",
			7794 => "11111110011001000111101111010101",
			7795 => "0000000111000000000111111000000100",
			7796 => "11111110100011100111101111010101",
			7797 => "00000000000110110111101111010101",
			7798 => "0000001001000000001001111000011000",
			7799 => "0000000011000000001000111000001100",
			7800 => "0000000101000000001101100000001000",
			7801 => "0000000001000000000110000000000100",
			7802 => "11111111010000010111101111010101",
			7803 => "00000001001101100111101111010101",
			7804 => "11111101001111000111101111010101",
			7805 => "0000001110000000000000110000000100",
			7806 => "11111011110011100111101111010101",
			7807 => "0000001111000000001011110100000100",
			7808 => "11111110000111000111101111010101",
			7809 => "00000000111010100111101111010101",
			7810 => "0000000101000000001001110000000100",
			7811 => "11111110111100100111101111010101",
			7812 => "0000000110000000001101111100001000",
			7813 => "0000001001000000001001111000000100",
			7814 => "00000000111101100111101111010101",
			7815 => "00000010000001100111101111010101",
			7816 => "0000001110000000000100010100000100",
			7817 => "00000001001000010111101111010101",
			7818 => "11111111010110010111101111010101",
			7819 => "0000000010000000001010001000110000",
			7820 => "0000001011000000001011000100010100",
			7821 => "0000000011000000001101100000001000",
			7822 => "0000000000000000000000110000000100",
			7823 => "11111101101110010111101111010101",
			7824 => "11111111101001000111101111010101",
			7825 => "0000000111000000000100010100001000",
			7826 => "0000001110000000001011000100000100",
			7827 => "00000001110011000111101111010101",
			7828 => "11111110011111100111101111010101",
			7829 => "00000010110010100111101111010101",
			7830 => "0000000101000000001100101100010000",
			7831 => "0000000111000000001011000100001000",
			7832 => "0000000101000000001100110000000100",
			7833 => "11111100110101110111101111010101",
			7834 => "11111110011101110111101111010101",
			7835 => "0000000111000000000000101000000100",
			7836 => "11111111101011110111101111010101",
			7837 => "11111110011010100111101111010101",
			7838 => "0000001001000000000110101000001000",
			7839 => "0000001110000000001011000100000100",
			7840 => "00000000000001110111101111010101",
			7841 => "00000010101101010111101111010101",
			7842 => "11111110001010110111101111010101",
			7843 => "0000001100000000000111111000010000",
			7844 => "0000000010000000000011001000000100",
			7845 => "00000000100001100111101111010101",
			7846 => "0000000010000000001100010100000100",
			7847 => "11111100110011110111101111010101",
			7848 => "0000001110000000001100001000000100",
			7849 => "00000001101110100111101111010101",
			7850 => "11111110101011010111101111010101",
			7851 => "0000000000000000000000110000001000",
			7852 => "0000001000000000001001101000000100",
			7853 => "00000000000000000111101111010101",
			7854 => "00000010100110110111101111010101",
			7855 => "0000001011000000000000101000001000",
			7856 => "0000000110000000001101111100000100",
			7857 => "11111111010110110111101111010101",
			7858 => "00000001101000110111101111010101",
			7859 => "0000000110000000000100110100000100",
			7860 => "00000001001000110111101111010101",
			7861 => "11111111000000010111101111010101",
			7862 => "0000000001000000001110100000001100",
			7863 => "0000001011000000001100001000001000",
			7864 => "0000000011000000000110000100000100",
			7865 => "00000010000101010111101111010101",
			7866 => "11111111111100100111101111010101",
			7867 => "00000011000011110111101111010101",
			7868 => "0000001110000000000100010100110100",
			7869 => "0000001011000000000000101000010100",
			7870 => "0000000000000000000010111100000100",
			7871 => "00000001011000000111101111010101",
			7872 => "0000000000000000000000110000001000",
			7873 => "0000000001000000001110100000000100",
			7874 => "11111111111111000111101111010101",
			7875 => "11111101010111100111101111010101",
			7876 => "0000001110000000000111111000000100",
			7877 => "00000010001000100111101111010101",
			7878 => "00000000001000000111101111010101",
			7879 => "0000001111000000000001011000010000",
			7880 => "0000000011000000001001110000001000",
			7881 => "0000000000000000001101010000000100",
			7882 => "11111111000000110111101111010101",
			7883 => "00000001100011100111101111010101",
			7884 => "0000001000000000001111001000000100",
			7885 => "00000000010011110111101111010101",
			7886 => "11111101100011010111101111010101",
			7887 => "0000000010000000001110000100001000",
			7888 => "0000001111000000000101100100000100",
			7889 => "00000001101000000111101111010101",
			7890 => "00000010111110010111101111010101",
			7891 => "0000000000000000000000111000000100",
			7892 => "11111111010100100111101111010101",
			7893 => "00000001011001110111101111010101",
			7894 => "0000000010000000001110000100100000",
			7895 => "0000000110000000000001111000010000",
			7896 => "0000001110000000000100000000001000",
			7897 => "0000001010000000000111110100000100",
			7898 => "00000000000000000111101111010101",
			7899 => "00000010010010010111101111010101",
			7900 => "0000001010000000000011101000000100",
			7901 => "00000000110011010111101111010101",
			7902 => "11111111000100000111101111010101",
			7903 => "0000000110000000000100110100001000",
			7904 => "0000000011000000001010111100000100",
			7905 => "11111111000011000111101111010101",
			7906 => "00000000100010000111101111010101",
			7907 => "0000000011000000001101111000000100",
			7908 => "11111101011001100111101111010101",
			7909 => "11111110011101010111101111010101",
			7910 => "0000000111000000001100001000010000",
			7911 => "0000000111000000001100001000001000",
			7912 => "0000000010000000000111011000000100",
			7913 => "00000000001010000111101111010101",
			7914 => "11111110000111000111101111010101",
			7915 => "0000000111000000001100001000000100",
			7916 => "00000001110001010111101111010101",
			7917 => "00000000010000110111101111010101",
			7918 => "0000001011000000000100000000001000",
			7919 => "0000000111000000000100000000000100",
			7920 => "11111110011101010111101111010101",
			7921 => "00000000000000000111101111010101",
			7922 => "0000001001000000001101101000000100",
			7923 => "11111111110000000111101111010101",
			7924 => "00000000001100110111101111010101",
			7925 => "0000001110000000000101101111001100",
			7926 => "0000001111000000000101110101110000",
			7927 => "0000000011000000000110000101000000",
			7928 => "0000001001000000000111100100100000",
			7929 => "0000000001000000001100110100010000",
			7930 => "0000001001000000000110101000001000",
			7931 => "0000000000000000000011111100000100",
			7932 => "00000000011001010111111010101011",
			7933 => "11111111111100100111111010101011",
			7934 => "0000000111000000001011000100000100",
			7935 => "11111111010001000111111010101011",
			7936 => "00000001010011010111111010101011",
			7937 => "0000000011000000000011011100001000",
			7938 => "0000000010000000001101000100000100",
			7939 => "11111110100111110111111010101011",
			7940 => "00000000100011000111111010101011",
			7941 => "0000000111000000000000101000000100",
			7942 => "11111111111110000111111010101011",
			7943 => "11111110010010100111111010101011",
			7944 => "0000001111000000000100000100010000",
			7945 => "0000001100000000000000101000001000",
			7946 => "0000001111000000001010011100000100",
			7947 => "00000001111010010111111010101011",
			7948 => "11111111101110100111111010101011",
			7949 => "0000000111000000001100001000000100",
			7950 => "11111101010101100111111010101011",
			7951 => "11111111010001110111111010101011",
			7952 => "0000001111000000000100010000001000",
			7953 => "0000000010000000001100100100000100",
			7954 => "00000010101010010111111010101011",
			7955 => "00000000100111110111111010101011",
			7956 => "0000000010000000000101110000000100",
			7957 => "00000011100100110111111010101011",
			7958 => "00000001011101010111111010101011",
			7959 => "0000001101000000000001111100100000",
			7960 => "0000001110000000001000111100010000",
			7961 => "0000000001000000001100110100001000",
			7962 => "0000000010000000000010011100000100",
			7963 => "11111111110100010111111010101011",
			7964 => "11111101110101000111111010101011",
			7965 => "0000001111000000000101100100000100",
			7966 => "11111110000100000111111010101011",
			7967 => "00000000110010110111111010101011",
			7968 => "0000001100000000000000101000001000",
			7969 => "0000000000000000000010111100000100",
			7970 => "11111111101111010111111010101011",
			7971 => "11111110100111110111111010101011",
			7972 => "0000001110000000000011011100000100",
			7973 => "11111101101011000111111010101011",
			7974 => "11111111000101110111111010101011",
			7975 => "0000000100000000001101001000001100",
			7976 => "0000000100000000001110100100001000",
			7977 => "0000000101000000001010111100000100",
			7978 => "00000000111101110111111010101011",
			7979 => "11111110111011110111111010101011",
			7980 => "00000010011110100111111010101011",
			7981 => "11111111001110010111111010101011",
			7982 => "0000000000000000000000110000111000",
			7983 => "0000001101000000001100101100011100",
			7984 => "0000000111000000000100010100001100",
			7985 => "0000000101000000001100110000001000",
			7986 => "0000001100000000001110111100000100",
			7987 => "11111110110011110111111010101011",
			7988 => "00000010001111010111111010101011",
			7989 => "11111110001111000111111010101011",
			7990 => "0000000100000000001000001000001000",
			7991 => "0000000110000000001101111100000100",
			7992 => "00000001110110110111111010101011",
			7993 => "00000011111100110111111010101011",
			7994 => "0000000100000000000011001100000100",
			7995 => "11111111110111010111111010101011",
			7996 => "00000001101010110111111010101011",
			7997 => "0000001011000000001100001000001100",
			7998 => "0000000011000000001101111000001000",
			7999 => "0000001101000000001110001100000100",
			8000 => "11111110110010000111111010101011",
			8001 => "00000000101110110111111010101011",
			8002 => "11111101100010010111111010101011",
			8003 => "0000000010000000000010011100001000",
			8004 => "0000001001000000001101101000000100",
			8005 => "11111110101011110111111010101011",
			8006 => "00000000001011010111111010101011",
			8007 => "0000000111000000001000111000000100",
			8008 => "00000000100111010111111010101011",
			8009 => "00000010001000010111111010101011",
			8010 => "0000001011000000000101101100011100",
			8011 => "0000001001000000000111100100001100",
			8012 => "0000000001000000001100110100001000",
			8013 => "0000000100000000000101010100000100",
			8014 => "11111110110100000111111010101011",
			8015 => "00000000000111010111111010101011",
			8016 => "11111101001111010111111010101011",
			8017 => "0000000111000000001011000100001000",
			8018 => "0000001110000000001101100000000100",
			8019 => "00000010110010100111111010101011",
			8020 => "00000000100101010111111010101011",
			8021 => "0000000000000000001010000000000100",
			8022 => "11111111010110110111111010101011",
			8023 => "00000000011111010111111010101011",
			8024 => "0000000111000000001101100000000100",
			8025 => "11111011111101010111111010101011",
			8026 => "00000000000000000111111010101011",
			8027 => "0000001001000000001101101000111000",
			8028 => "0000001111000000000111100000110000",
			8029 => "0000000110000000001100011000011100",
			8030 => "0000001111000000000010110100010000",
			8031 => "0000000100000000000010111000001000",
			8032 => "0000000011000000001101111000000100",
			8033 => "00000000011110000111111010101011",
			8034 => "11111110001011000111111010101011",
			8035 => "0000001110000000000110000100000100",
			8036 => "00000001000011010111111010101011",
			8037 => "11111110011011110111111010101011",
			8038 => "0000001101000000001100101000001000",
			8039 => "0000000000000000000011010000000100",
			8040 => "00000001011101010111111010101011",
			8041 => "11111111000111000111111010101011",
			8042 => "00000010010101100111111010101011",
			8043 => "0000000100000000001111100000001100",
			8044 => "0000000010000000001110010000000100",
			8045 => "00000000101010010111111010101011",
			8046 => "0000000101000000000000001100000100",
			8047 => "11111110101101000111111010101011",
			8048 => "11111101100101100111111010101011",
			8049 => "0000001110000000000110000100000100",
			8050 => "00000001010011100111111010101011",
			8051 => "11111111101110000111111010101011",
			8052 => "0000000011000000001010111000000100",
			8053 => "00000010001010000111111010101011",
			8054 => "00000000001111000111111010101011",
			8055 => "0000000000000000001111000100110100",
			8056 => "0000000001000000001001111000011100",
			8057 => "0000000111000000000100000000001100",
			8058 => "0000000010000000000100101000001000",
			8059 => "0000000110000000000100110100000100",
			8060 => "11111110110001100111111010101011",
			8061 => "00000001011101110111111010101011",
			8062 => "00000010000010010111111010101011",
			8063 => "0000000111000000001000111000001000",
			8064 => "0000000100000000001011110000000100",
			8065 => "00000000111010010111111010101011",
			8066 => "00000011000011100111111010101011",
			8067 => "0000000101000000001010111100000100",
			8068 => "11111110011001000111111010101011",
			8069 => "00000001010101110111111010101011",
			8070 => "0000001001000000001111001100001000",
			8071 => "0000000000000000001000101100000100",
			8072 => "00000000000000000111111010101011",
			8073 => "11111110000001100111111010101011",
			8074 => "0000001001000000000100110100001000",
			8075 => "0000000100000000001000000100000100",
			8076 => "00000000000110000111111010101011",
			8077 => "00000010001011010111111010101011",
			8078 => "0000000110000000001001111100000100",
			8079 => "11111110011100110111111010101011",
			8080 => "00000000000000000111111010101011",
			8081 => "0000000100000000001100001100010100",
			8082 => "0000001100000000001001110000010000",
			8083 => "0000000111000000000100000000001000",
			8084 => "0000001100000000000100000000000100",
			8085 => "11111111001000010111111010101011",
			8086 => "00000010010011110111111010101011",
			8087 => "0000001100000000001000111100000100",
			8088 => "11111110001110100111111010101011",
			8089 => "11111111011111110111111010101011",
			8090 => "00000010001001010111111010101011",
			8091 => "0000001001000000001011101000010000",
			8092 => "0000000001000000000010001100001000",
			8093 => "0000000101000000000001111100000100",
			8094 => "11111111110110010111111010101011",
			8095 => "00000001011111010111111010101011",
			8096 => "0000001100000000000000101000000100",
			8097 => "11111111110110010111111010101011",
			8098 => "11111111000010100111111010101011",
			8099 => "0000000011000000001000000000001000",
			8100 => "0000000100000000001111100000000100",
			8101 => "00000001010101000111111010101011",
			8102 => "11111101101100110111111010101011",
			8103 => "0000000100000000001000001000000100",
			8104 => "00000000100101000111111010101011",
			8105 => "11111111101000000111111010101011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(2753, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(5446, initial_addr_3'length));
	end generate gen_rom_7;

	gen_rom_8: if SELECT_ROM = 8 generate
		bank <= (
			0 => "00000000000000000000000000000101",
			1 => "00000000000000000000000000001001",
			2 => "0000000101000000001111010100000100",
			3 => "00000000000000000000000000010101",
			4 => "11111110110100000000000000010101",
			5 => "0000000100000000000101010100000100",
			6 => "11111111111111010000000000101001",
			7 => "0000000100000000000001100100000100",
			8 => "00000000001001110000000000101001",
			9 => "00000000000000000000000000101001",
			10 => "0000000100000000000011010100000100",
			11 => "11111111111111010000000000111101",
			12 => "0000000100000000000001100100000100",
			13 => "00000000000011100000000000111101",
			14 => "00000000000000000000000000111101",
			15 => "0000001000000000000110001000001000",
			16 => "0000001000000000000001010100000100",
			17 => "00000000000000000000000001010001",
			18 => "00000000000011100000000001010001",
			19 => "00000000000000000000000001010001",
			20 => "0000001011000000000010011100001000",
			21 => "0000001001000000001001111100000100",
			22 => "00000000000000000000000001100101",
			23 => "00000000000000010000000001100101",
			24 => "11111111010101000000000001100101",
			25 => "0000000111000000000001001000001100",
			26 => "0000000100000000000100001100000100",
			27 => "00000000000000000000000010000001",
			28 => "0000000100000000000001100100000100",
			29 => "00000000001011110000000010000001",
			30 => "00000000000000000000000010000001",
			31 => "11111111011101000000000010000001",
			32 => "0000000111000000000001001000001100",
			33 => "0000000100000000000000010100000100",
			34 => "00000000000000000000000010011101",
			35 => "0000000100000000000001100100000100",
			36 => "00000000000110010000000010011101",
			37 => "00000000000000000000000010011101",
			38 => "11111111100110100000000010011101",
			39 => "0000001010000000000110011000001100",
			40 => "0000001010000000001001000100000100",
			41 => "00000000000000000000000011000001",
			42 => "0000000110000000001111000000000100",
			43 => "00000000000000000000000011000001",
			44 => "00000000000110000000000011000001",
			45 => "0000001010000000000110011100000100",
			46 => "11111111110110010000000011000001",
			47 => "00000000000000000000000011000001",
			48 => "0000000001000000001100011000001100",
			49 => "0000001010000000000110011100001000",
			50 => "0000001010000000001000010100000100",
			51 => "00000000000000000000000011100101",
			52 => "11111111110111110000000011100101",
			53 => "00000000000000000000000011100101",
			54 => "0000001010000000001010110000000100",
			55 => "00000000001101100000000011100101",
			56 => "00000000000000000000000011100101",
			57 => "0000001100000000001011011100001100",
			58 => "0000001001000000001001111100000100",
			59 => "00000000000000000000000100001001",
			60 => "0000001001000000001000010100000100",
			61 => "00000000000010100000000100001001",
			62 => "00000000000000000000000100001001",
			63 => "0000001100000000001011011100000100",
			64 => "11111111010101100000000100001001",
			65 => "00000000000000000000000100001001",
			66 => "0000001010000000000110011000001100",
			67 => "0000000000000000000010101000000100",
			68 => "00000000000000000000000100110101",
			69 => "0000000110000000001111000000000100",
			70 => "00000000000000000000000100110101",
			71 => "00000000010101110000000100110101",
			72 => "0000000110000000001000010000000100",
			73 => "00000000000000000000000100110101",
			74 => "0000000000000000001000110000000100",
			75 => "00000000000000000000000100110101",
			76 => "11111111110110110000000100110101",
			77 => "0000001000000000001011010100001100",
			78 => "0000000100000000000011110000000100",
			79 => "00000000000000000000000101100001",
			80 => "0000000100000000001111100000000100",
			81 => "00000000000110100000000101100001",
			82 => "00000000000000000000000101100001",
			83 => "0000001110000000000011010100001000",
			84 => "0000000100000000000000101100000100",
			85 => "11111111100100100000000101100001",
			86 => "00000000000000000000000101100001",
			87 => "00000000000000000000000101100001",
			88 => "0000000111000000000001001000010000",
			89 => "0000001001000000001001111100000100",
			90 => "00000000000000000000000110000101",
			91 => "0000000100000000000011110000000100",
			92 => "00000000000000000000000110000101",
			93 => "0000001100000000001000000000000100",
			94 => "00000000000000000000000110000101",
			95 => "00000000010010100000000110000101",
			96 => "11111111000000100000000110000101",
			97 => "0000000101000000000000010000010000",
			98 => "0000000111000000000001011000000100",
			99 => "00000000000000000000000110101001",
			100 => "0000000101000000001110010000000100",
			101 => "00000000000000000000000110101001",
			102 => "0000001011000000000001001000000100",
			103 => "00000000000000000000000110101001",
			104 => "00000000001100010000000110101001",
			105 => "11111111111110110000000110101001",
			106 => "0000001111000000001110100100000100",
			107 => "00000000000000000000000111001101",
			108 => "0000000001000000001111000000001100",
			109 => "0000000110000000000100111100000100",
			110 => "00000000000000000000000111001101",
			111 => "0000000011000000000011101100000100",
			112 => "11111111100100000000000111001101",
			113 => "00000000000000000000000111001101",
			114 => "00000000000000000000000111001101",
			115 => "0000001100000000001011011100010000",
			116 => "0000001001000000001001111100000100",
			117 => "00000000000000000000000111111001",
			118 => "0000001100000000001001110100000100",
			119 => "00000000000000000000000111111001",
			120 => "0000001001000000001000010100000100",
			121 => "00000000001000000000000111111001",
			122 => "00000000000000000000000111111001",
			123 => "0000001100000000001011011100000100",
			124 => "11111111010010110000000111111001",
			125 => "00000000000000000000000111111001",
			126 => "0000000111000000000001001000010100",
			127 => "0000000100000000000000010100001000",
			128 => "0000000001000000001101011000000100",
			129 => "11111111111110000000001000100101",
			130 => "00000000000000000000001000100101",
			131 => "0000001001000000001001111100000100",
			132 => "00000000000000000000001000100101",
			133 => "0000001100000000001001110100000100",
			134 => "00000000000000000000001000100101",
			135 => "00000000010101100000001000100101",
			136 => "11111111000110110000001000100101",
			137 => "0000000100000000000000010100001100",
			138 => "0000000100000000001110100100000100",
			139 => "00000000000000000000001001011001",
			140 => "0000001111000000001010110100000100",
			141 => "11111111111011000000001001011001",
			142 => "00000000000000000000001001011001",
			143 => "0000000100000000000001100100001100",
			144 => "0000000010000000001101101100000100",
			145 => "00000000000000000000001001011001",
			146 => "0000000010000000001110100100000100",
			147 => "00000000001100110000001001011001",
			148 => "00000000000000000000001001011001",
			149 => "00000000000000000000001001011001",
			150 => "0000001011000000000110100000010100",
			151 => "0000000101000000001001010100000100",
			152 => "00000000000000000000001010001101",
			153 => "0000001010000000000101000100001100",
			154 => "0000001010000000001000010100000100",
			155 => "00000000000000000000001010001101",
			156 => "0000000011000000000010111000000100",
			157 => "00000000010100110000001010001101",
			158 => "00000000000000000000001010001101",
			159 => "00000000000000000000001010001101",
			160 => "0000001101000000001111010100000100",
			161 => "00000000000000000000001010001101",
			162 => "11111111111011010000001010001101",
			163 => "0000001000000000001111001000010100",
			164 => "0000000010000000000110111000000100",
			165 => "00000000000000000000001011000001",
			166 => "0000001100000000001000000000000100",
			167 => "00000000000000000000001011000001",
			168 => "0000001100000000001011011100001000",
			169 => "0000000000000000000001110100000100",
			170 => "00000000000000000000001011000001",
			171 => "00000000000111000000001011000001",
			172 => "00000000000000000000001011000001",
			173 => "0000000010000000001110000000000100",
			174 => "00000000000000000000001011000001",
			175 => "11111111100111110000001011000001",
			176 => "0000000111000000000001001000010100",
			177 => "0000001100000000000100011000000100",
			178 => "00000000000000000000001011101101",
			179 => "0000000110000000000100101100001100",
			180 => "0000000010000000001101101100000100",
			181 => "00000000000000000000001011101101",
			182 => "0000000110000000001111000000000100",
			183 => "00000000000000000000001011101101",
			184 => "00000000000110100000001011101101",
			185 => "00000000000000000000001011101101",
			186 => "11111111110100100000001011101101",
			187 => "0000000100000000000000010100001100",
			188 => "0000000110000000000100111100000100",
			189 => "00000000000000000000001100101001",
			190 => "0000001111000000001010110100000100",
			191 => "11111111110110010000001100101001",
			192 => "00000000000000000000001100101001",
			193 => "0000000110000000001001111100010000",
			194 => "0000000101000000001001010100000100",
			195 => "00000000000000000000001100101001",
			196 => "0000001101000000001100010000001000",
			197 => "0000000100000000000001100100000100",
			198 => "00000000010100010000001100101001",
			199 => "00000000000000000000001100101001",
			200 => "00000000000000000000001100101001",
			201 => "00000000000000000000001100101001",
			202 => "0000000111000000001011110100010100",
			203 => "0000001001000000001001111100000100",
			204 => "00000000000000000000001101100101",
			205 => "0000000010000000000110111000000100",
			206 => "00000000000000000000001101100101",
			207 => "0000001000000000000111000100001000",
			208 => "0000001100000000001001110100000100",
			209 => "00000000000000000000001101100101",
			210 => "00000000010010000000001101100101",
			211 => "00000000000000000000001101100101",
			212 => "0000000110000000001000010000000100",
			213 => "00000000000000000000001101100101",
			214 => "0000001011000000001101000100000100",
			215 => "00000000000000000000001101100101",
			216 => "11111111001101000000001101100101",
			217 => "0000000111000000001000011000010100",
			218 => "0000000111000000001011000000000100",
			219 => "00000000000000000000001110101001",
			220 => "0000000100000000001000001000000100",
			221 => "00000000000000000000001110101001",
			222 => "0000001010000000000001010100001000",
			223 => "0000001111000000001000110100000100",
			224 => "00000001010010100000001110101001",
			225 => "00000000000000000000001110101001",
			226 => "00000000000000000000001110101001",
			227 => "0000001000000000000110001000000100",
			228 => "00000000000000000000001110101001",
			229 => "0000001110000000000011010100001000",
			230 => "0000000110000000001000010000000100",
			231 => "00000000000000000000001110101001",
			232 => "11111111011011110000001110101001",
			233 => "00000000000000000000001110101001",
			234 => "0000000010000000001011110000010000",
			235 => "0000000010000000001101101100000100",
			236 => "00000000000000000000001111101101",
			237 => "0000000110000000001000010000001000",
			238 => "0000000110000000001111000000000100",
			239 => "00000000000000000000001111101101",
			240 => "00000000010011110000001111101101",
			241 => "00000000000000000000001111101101",
			242 => "0000001000000000000001010100000100",
			243 => "00000000000000000000001111101101",
			244 => "0000000110000000000100111100000100",
			245 => "00000000000000000000001111101101",
			246 => "0000000100000000001110100100000100",
			247 => "00000000000000000000001111101101",
			248 => "0000001010000000001000010100000100",
			249 => "00000000000000000000001111101101",
			250 => "11111111110011110000001111101101",
			251 => "0000001001000000001010100000001100",
			252 => "0000001111000000001110100100001000",
			253 => "0000000100000000000111011100000100",
			254 => "11111111011101110000010000111001",
			255 => "00000000000000000000010000111001",
			256 => "00000000000000000000010000111001",
			257 => "0000001111000000001100001100001100",
			258 => "0000001100000000000100000100001000",
			259 => "0000000111000000000111010000000100",
			260 => "00000000000000000000010000111001",
			261 => "00000000110100010000010000111001",
			262 => "00000000000000000000010000111001",
			263 => "0000000100000000000000010100001100",
			264 => "0000001001000000001000100100001000",
			265 => "0000000100000000000011110000000100",
			266 => "00000000000000000000010000111001",
			267 => "11111111110001000000010000111001",
			268 => "00000000000000000000010000111001",
			269 => "00000000000000000000010000111001",
			270 => "0000001010000000000110011000010100",
			271 => "0000001010000000001000010100000100",
			272 => "00000000000000000000010010001101",
			273 => "0000000010000000000110111000000100",
			274 => "00000000000000000000010010001101",
			275 => "0000000101000000001100010000001000",
			276 => "0000001100000000001001110100000100",
			277 => "00000000000000000000010010001101",
			278 => "00000001000100110000010010001101",
			279 => "00000000000000000000010010001101",
			280 => "0000000100000000001011001000001100",
			281 => "0000001001000000001000100100001000",
			282 => "0000001000000000001100000100000100",
			283 => "00000000000000000000010010001101",
			284 => "11111111110000010000010010001101",
			285 => "00000000000000000000010010001101",
			286 => "0000001010000000000101000100001000",
			287 => "0000001010000000001100011100000100",
			288 => "00000000000000000000010010001101",
			289 => "00000000000111000000010010001101",
			290 => "00000000000000000000010010001101",
			291 => "0000000110000000000101010000011000",
			292 => "0000001101000000001010000100010100",
			293 => "0000000110000000001111000000000100",
			294 => "00000000000000000000010011001001",
			295 => "0000001101000000001110101100000100",
			296 => "00000000000000000000010011001001",
			297 => "0000001010000000001000100100000100",
			298 => "00000000000000000000010011001001",
			299 => "0000000110000000001000010000000100",
			300 => "00000000010111100000010011001001",
			301 => "00000000000000000000010011001001",
			302 => "00000000000000000000010011001001",
			303 => "0000001000000000001001101000000100",
			304 => "00000000000000000000010011001001",
			305 => "11111111111111110000010011001001",
			306 => "0000001000000000000110001000011000",
			307 => "0000000100000000001110100100000100",
			308 => "00000000000000000000010100000101",
			309 => "0000001100000000001001110100000100",
			310 => "00000000000000000000010100000101",
			311 => "0000000111000000001011110100001100",
			312 => "0000000001000000001110010100000100",
			313 => "00000000000000000000010100000101",
			314 => "0000001000000000000101000100000100",
			315 => "00000000000000000000010100000101",
			316 => "00000000011000000000010100000101",
			317 => "00000000000000000000010100000101",
			318 => "0000000100000000001001000000000100",
			319 => "11111111010001000000010100000101",
			320 => "00000000000000000000010100000101",
			321 => "0000000100000000000000101100100000",
			322 => "0000001001000000000111101100001000",
			323 => "0000000100000000000111011100000100",
			324 => "11111111101110010000010101011001",
			325 => "00000000000000000000010101011001",
			326 => "0000000110000000001000010000001000",
			327 => "0000001001000000001010100100000100",
			328 => "00000000000000000000010101011001",
			329 => "00000000011001000000010101011001",
			330 => "0000000100000000000000010100001000",
			331 => "0000001001000000000011101000000100",
			332 => "11111111101111010000010101011001",
			333 => "00000000000000000000010101011001",
			334 => "0000001001000000001000010100000100",
			335 => "00000000000111110000010101011001",
			336 => "00000000000000000000010101011001",
			337 => "0000001010000000000101000100001000",
			338 => "0000001100000000000001111100000100",
			339 => "00000000000000000000010101011001",
			340 => "00000001110110110000010101011001",
			341 => "00000000000000000000010101011001",
			342 => "0000000100000000000100001100011000",
			343 => "0000000001000000001101011000010100",
			344 => "0000001000000000000101000100000100",
			345 => "00000000000000000000010110100101",
			346 => "0000000101000000001110110100001100",
			347 => "0000000000000000000001110100000100",
			348 => "00000000000000000000010110100101",
			349 => "0000001011000000001101000100000100",
			350 => "11111111100000100000010110100101",
			351 => "00000000000000000000010110100101",
			352 => "00000000000000000000010110100101",
			353 => "00000000000000000000010110100101",
			354 => "0000001000000000000111000100001100",
			355 => "0000000001000000001011111100000100",
			356 => "00000000000000000000010110100101",
			357 => "0000000000000000000010111100000100",
			358 => "00000000000000000000010110100101",
			359 => "00000000011010100000010110100101",
			360 => "00000000000000000000010110100101",
			361 => "0000000100000000000000010100011000",
			362 => "0000001011000000000000110100010100",
			363 => "0000000111000000001011011100010000",
			364 => "0000001100000000001111011100001100",
			365 => "0000000001000000001011001100001000",
			366 => "0000001000000000000101000100000100",
			367 => "00000000000000000000010111110001",
			368 => "11111111101011010000010111110001",
			369 => "00000000000000000000010111110001",
			370 => "00000000000000000000010111110001",
			371 => "00000000000000000000010111110001",
			372 => "00000000000000000000010111110001",
			373 => "0000001000000000001111001000001100",
			374 => "0000000001000000001011111100000100",
			375 => "00000000000000000000010111110001",
			376 => "0000000111000000000111110000000100",
			377 => "00000000101101110000010111110001",
			378 => "00000000000000000000010111110001",
			379 => "00000000000000000000010111110001",
			380 => "0000000101000000001001100000011100",
			381 => "0000001100000000001001110100001000",
			382 => "0000000100000000000000101100000100",
			383 => "11111111111011100000011001000101",
			384 => "00000000000000000000011001000101",
			385 => "0000001000000000000111000100010000",
			386 => "0000001110000000001000011100001100",
			387 => "0000000100000000001110100100000100",
			388 => "00000000000000000000011001000101",
			389 => "0000001001000000001001111100000100",
			390 => "00000000000000000000011001000101",
			391 => "00000000110110000000011001000101",
			392 => "00000000000000000000011001000101",
			393 => "00000000000000000000011001000101",
			394 => "0000000110000000001000010000000100",
			395 => "00000000000000000000011001000101",
			396 => "0000001011000000000110100000000100",
			397 => "00000000000000000000011001000101",
			398 => "0000000111000000000100010000000100",
			399 => "00000000000000000000011001000101",
			400 => "11111111110001010000011001000101",
			401 => "0000000101000000001110000100010000",
			402 => "0000000001000000001001011000000100",
			403 => "00000000000000000000011010100001",
			404 => "0000000100000000001111100000000100",
			405 => "00000000000000000000011010100001",
			406 => "0000001100000000001010111100000100",
			407 => "00000000000000000000011010100001",
			408 => "00000001101001110000011010100001",
			409 => "0000000001000000001010011000010000",
			410 => "0000000111000000001111011100000100",
			411 => "00000000000000000000011010100001",
			412 => "0000001010000000001000010100000100",
			413 => "00000000000000000000011010100001",
			414 => "0000001000000000000001010100000100",
			415 => "00000000000000000000011010100001",
			416 => "11111111100101110000011010100001",
			417 => "0000001000000000000001110100001100",
			418 => "0000000111000000000111010000000100",
			419 => "00000000000000000000011010100001",
			420 => "0000000000000000001010101100000100",
			421 => "00000000000000000000011010100001",
			422 => "00000000010100100000011010100001",
			423 => "00000000000000000000011010100001",
			424 => "0000001001000000001010100000001100",
			425 => "0000001111000000001110100100001000",
			426 => "0000000100000000000111011100000100",
			427 => "11111111100000000000011011111101",
			428 => "00000000000000000000011011111101",
			429 => "00000000000000000000011011111101",
			430 => "0000001110000000001000011100010100",
			431 => "0000001100000000000100000100010000",
			432 => "0000000110000000001001111100001100",
			433 => "0000000101000000001001010000000100",
			434 => "00000000000000000000011011111101",
			435 => "0000001011000000000100010000000100",
			436 => "00000000000000000000011011111101",
			437 => "00000000110001000000011011111101",
			438 => "00000000000000000000011011111101",
			439 => "00000000000000000000011011111101",
			440 => "0000001001000000001000100100001100",
			441 => "0000001100000000001001110100000100",
			442 => "00000000000000000000011011111101",
			443 => "0000000111000000000111110000000100",
			444 => "11111111101110100000011011111101",
			445 => "00000000000000000000011011111101",
			446 => "00000000000000000000011011111101",
			447 => "0000000010000000001011110000010100",
			448 => "0000000010000000001101101100000100",
			449 => "00000000000000000000011101100001",
			450 => "0000001100000000001010111000000100",
			451 => "00000000000000000000011101100001",
			452 => "0000001001000000001011001100000100",
			453 => "00000000000000000000011101100001",
			454 => "0000001111000000000010010100000100",
			455 => "00000001011110000000011101100001",
			456 => "00000000000000000000011101100001",
			457 => "0000001101000000000110111100001100",
			458 => "0000000001000000001100011000000100",
			459 => "00000000000000000000011101100001",
			460 => "0000001000000000001111001000000100",
			461 => "00000000001011110000011101100001",
			462 => "00000000000000000000011101100001",
			463 => "0000001001000000001000100100010000",
			464 => "0000001100000000001111011100000100",
			465 => "00000000000000000000011101100001",
			466 => "0000000011000000001110100100000100",
			467 => "00000000000000000000011101100001",
			468 => "0000000001000000001010011000000100",
			469 => "00000000000000000000011101100001",
			470 => "11111111101010000000011101100001",
			471 => "00000000000000000000011101100001",
			472 => "0000001101000000001010000100100000",
			473 => "0000001100000000001001110100001000",
			474 => "0000000100000000000000101100000100",
			475 => "11111111111100010000011110101101",
			476 => "00000000000000000000011110101101",
			477 => "0000000100000000001110100100000100",
			478 => "00000000000000000000011110101101",
			479 => "0000001000000000000111000100010000",
			480 => "0000001110000000001000011100001100",
			481 => "0000001100000000000001011000001000",
			482 => "0000000001000000001110010100000100",
			483 => "00000000000000000000011110101101",
			484 => "00000000110010110000011110101101",
			485 => "00000000000000000000011110101101",
			486 => "00000000000000000000011110101101",
			487 => "00000000000000000000011110101101",
			488 => "0000000001000000001101011000000100",
			489 => "00000000000000000000011110101101",
			490 => "11111111110101110000011110101101",
			491 => "0000001101000000000110111100011100",
			492 => "0000000111000000001011000000000100",
			493 => "00000000000000000000011111111001",
			494 => "0000000110000000000101010000010100",
			495 => "0000001001000000000011101000010000",
			496 => "0000000110000000001001100100000100",
			497 => "00000000000000000000011111111001",
			498 => "0000001001000000001011001100000100",
			499 => "00000000000000000000011111111001",
			500 => "0000000010000000001100111000000100",
			501 => "00000000000000000000011111111001",
			502 => "00000000100001000000011111111001",
			503 => "00000000000000000000011111111001",
			504 => "00000000000000000000011111111001",
			505 => "0000000010000000001000000100000100",
			506 => "00000000000000000000011111111001",
			507 => "0000000110000000001000010000000100",
			508 => "00000000000000000000011111111001",
			509 => "11111111111100100000011111111001",
			510 => "0000000100000000000011011000100100",
			511 => "0000001000000000000110001000011000",
			512 => "0000001001000000000111101100000100",
			513 => "00000000000000000000100001010101",
			514 => "0000001011000000000110100000010000",
			515 => "0000001110000000001000011100001100",
			516 => "0000000011000000000001011100000100",
			517 => "00000000000000000000100001010101",
			518 => "0000001011000000000100010000000100",
			519 => "00000000000000000000100001010101",
			520 => "00000000101010000000100001010101",
			521 => "00000000000000000000100001010101",
			522 => "00000000000000000000100001010101",
			523 => "0000000100000000001001000000001000",
			524 => "0000000011000000001110111000000100",
			525 => "11111111100010000000100001010101",
			526 => "00000000000000000000100001010101",
			527 => "00000000000000000000100001010101",
			528 => "0000001000000000001010101100001000",
			529 => "0000000110000000001000010000000100",
			530 => "00000000000000000000100001010101",
			531 => "00000001100100010000100001010101",
			532 => "00000000000000000000100001010101",
			533 => "0000001110000000000110111000011100",
			534 => "0000001100000000001001110100000100",
			535 => "00000000000000000000100010101001",
			536 => "0000001000000000000111000100010100",
			537 => "0000000011000000001011111000000100",
			538 => "00000000000000000000100010101001",
			539 => "0000001100000000000111010000001100",
			540 => "0000000010000000000010010100000100",
			541 => "00000000000000000000100010101001",
			542 => "0000001101000000001100010000000100",
			543 => "00000000110011010000100010101001",
			544 => "00000000000000000000100010101001",
			545 => "00000000000000000000100010101001",
			546 => "00000000000000000000100010101001",
			547 => "0000000100000000000110001100000100",
			548 => "00000000000000000000100010101001",
			549 => "0000001010000000001000010100000100",
			550 => "00000000000000000000100010101001",
			551 => "0000001111000000001000110100000100",
			552 => "00000000000000000000100010101001",
			553 => "11111111110001100000100010101001",
			554 => "0000000100000000000011011000101000",
			555 => "0000000001000000001010011000010100",
			556 => "0000000011000000000101000000010000",
			557 => "0000001000000000000101000100000100",
			558 => "00000000000000000000100100001101",
			559 => "0000000100000000000011101100001000",
			560 => "0000001001000000000011101000000100",
			561 => "11111111011110100000100100001101",
			562 => "00000000000000000000100100001101",
			563 => "00000000000000000000100100001101",
			564 => "00000000000000000000100100001101",
			565 => "0000001101000000001010000100010000",
			566 => "0000001111000000001001001100001100",
			567 => "0000000100000000001110100100000100",
			568 => "00000000000000000000100100001101",
			569 => "0000000101000000000101110000000100",
			570 => "00000000000000000000100100001101",
			571 => "00000000110000000000100100001101",
			572 => "00000000000000000000100100001101",
			573 => "00000000000000000000100100001101",
			574 => "0000001010000000000101000100001000",
			575 => "0000000001000000001001011000000100",
			576 => "00000000000000000000100100001101",
			577 => "00000010011001000000100100001101",
			578 => "00000000000000000000100100001101",
			579 => "0000000001000000000100110100010100",
			580 => "0000000100000000000111011100000100",
			581 => "11111111000000100000100110000001",
			582 => "0000001000000000000001110100001100",
			583 => "0000000000000000000000111000000100",
			584 => "00000000000000000000100110000001",
			585 => "0000000001000000001001011000000100",
			586 => "00000000000000000000100110000001",
			587 => "00000000100101100000100110000001",
			588 => "00000000000000000000100110000001",
			589 => "0000000011000000000110001100001100",
			590 => "0000001100000000000100000100001000",
			591 => "0000000111000000000111010000000100",
			592 => "00000000000000000000100110000001",
			593 => "00000000111101010000100110000001",
			594 => "00000000000000000000100110000001",
			595 => "0000001100000000000111010000010000",
			596 => "0000001111000000000110001100000100",
			597 => "00000000000000000000100110000001",
			598 => "0000001010000000001001000100000100",
			599 => "00000000000000000000100110000001",
			600 => "0000000111000000000100010000000100",
			601 => "11111111011010110000100110000001",
			602 => "00000000000000000000100110000001",
			603 => "0000000001000000000100111100001000",
			604 => "0000001100000000000100000100000100",
			605 => "00000000000000000000100110000001",
			606 => "00000000010111000000100110000001",
			607 => "00000000000000000000100110000001",
			608 => "0000000100000000000011011000101100",
			609 => "0000000001000000001010011000011000",
			610 => "0000001011000000001110101100010000",
			611 => "0000001000000000000101000100000100",
			612 => "00000000000000000000100111101101",
			613 => "0000000111000000001011011100001000",
			614 => "0000001000000000001100000100000100",
			615 => "11111111011001110000100111101101",
			616 => "00000000000000000000100111101101",
			617 => "00000000000000000000100111101101",
			618 => "0000001000000000001100000100000100",
			619 => "00000000000100010000100111101101",
			620 => "00000000000000000000100111101101",
			621 => "0000001101000000001010000100010000",
			622 => "0000001110000000001000001000001100",
			623 => "0000000101000000001110110100001000",
			624 => "0000000111000000000111010000000100",
			625 => "00000000000000000000100111101101",
			626 => "00000000101011000000100111101101",
			627 => "00000000000000000000100111101101",
			628 => "00000000000000000000100111101101",
			629 => "00000000000000000000100111101101",
			630 => "0000001010000000000101000100001000",
			631 => "0000000001000000001001011000000100",
			632 => "00000000000000000000100111101101",
			633 => "00000010001110010000100111101101",
			634 => "00000000000000000000100111101101",
			635 => "0000001000000000001100000100011100",
			636 => "0000001011000000001110101100010000",
			637 => "0000000001000000001010011000001100",
			638 => "0000000000000000001010101100000100",
			639 => "00000000000000000000101001100001",
			640 => "0000000000000000001000110000000100",
			641 => "11111111101011000000101001100001",
			642 => "00000000000000000000101001100001",
			643 => "00000000000000000000101001100001",
			644 => "0000000001000000001101011000001000",
			645 => "0000001001000000001010100100000100",
			646 => "00000000000000000000101001100001",
			647 => "00000000101111000000101001100001",
			648 => "00000000000000000000101001100001",
			649 => "0000000100000000000000010100001000",
			650 => "0000001001000000001000100100000100",
			651 => "11111111011101010000101001100001",
			652 => "00000000000000000000101001100001",
			653 => "0000000000000000000111111000010100",
			654 => "0000000110000000000100101100010000",
			655 => "0000000000000000000010011000000100",
			656 => "00000000000000000000101001100001",
			657 => "0000000110000000000100111100000100",
			658 => "00000000000000000000101001100001",
			659 => "0000000110000000001001111100000100",
			660 => "00000000010110010000101001100001",
			661 => "00000000000000000000101001100001",
			662 => "00000000000000000000101001100001",
			663 => "00000000000000000000101001100001",
			664 => "0000000000000000001011000100101000",
			665 => "0000000111000000001011011100011000",
			666 => "0000000001000000001010011000010100",
			667 => "0000001010000000000001010000010000",
			668 => "0000001000000000000101000100000100",
			669 => "00000000000000000000101010111101",
			670 => "0000001011000000001110101100001000",
			671 => "0000000000000000000001110100000100",
			672 => "00000000000000000000101010111101",
			673 => "11111111011101010000101010111101",
			674 => "00000000000000000000101010111101",
			675 => "00000000000000000000101010111101",
			676 => "00000000000000000000101010111101",
			677 => "0000000111000000001011110100001100",
			678 => "0000001000000000000111000100001000",
			679 => "0000000110000000001111000000000100",
			680 => "00000000000000000000101010111101",
			681 => "00000000001110010000101010111101",
			682 => "00000000000000000000101010111101",
			683 => "00000000000000000000101010111101",
			684 => "0000000000000000000000101000000100",
			685 => "00000000111101110000101010111101",
			686 => "00000000000000000000101010111101",
			687 => "0000000001000000000100110100010100",
			688 => "0000000100000000000111011100000100",
			689 => "11111111000101110000101100111001",
			690 => "0000001000000000000001110100001100",
			691 => "0000000000000000000000111000000100",
			692 => "00000000000000000000101100111001",
			693 => "0000000001000000001001011000000100",
			694 => "00000000000000000000101100111001",
			695 => "00000000011111110000101100111001",
			696 => "00000000000000000000101100111001",
			697 => "0000001110000000001000011100010100",
			698 => "0000001100000000000100000100010000",
			699 => "0000000111000000000111010000000100",
			700 => "00000000000000000000101100111001",
			701 => "0000001011000000000110100000001000",
			702 => "0000001100000000001001110100000100",
			703 => "00000000000000000000101100111001",
			704 => "00000000111111000000101100111001",
			705 => "00000000000000000000101100111001",
			706 => "00000000000000000000101100111001",
			707 => "0000001100000000000100000100010000",
			708 => "0000001001000000000111110100001100",
			709 => "0000001010000000001001000100000100",
			710 => "00000000000000000000101100111001",
			711 => "0000000001000000001011001100000100",
			712 => "11111111011000010000101100111001",
			713 => "00000000000000000000101100111001",
			714 => "00000000000000000000101100111001",
			715 => "0000000001000000000100111100000100",
			716 => "00000000010011100000101100111001",
			717 => "00000000000000000000101100111001",
			718 => "0000000100000000000000101100110000",
			719 => "0000000110000000000101010000100100",
			720 => "0000000010000000001000110100010100",
			721 => "0000000100000000000111011100010000",
			722 => "0000001000000000000001010100000100",
			723 => "00000000000000000000101110101101",
			724 => "0000000001000000001101011000001000",
			725 => "0000001111000000001000011100000100",
			726 => "11111111100001110000101110101101",
			727 => "00000000000000000000101110101101",
			728 => "00000000000000000000101110101101",
			729 => "00000000000000000000101110101101",
			730 => "0000001101000000001010000100001100",
			731 => "0000000001000000000111101000000100",
			732 => "00000000000000000000101110101101",
			733 => "0000001111000000000011001100000100",
			734 => "00000000110000000000101110101101",
			735 => "00000000000000000000101110101101",
			736 => "00000000000000000000101110101101",
			737 => "0000001001000000000111110100001000",
			738 => "0000000100000000000011101100000100",
			739 => "11111111100111000000101110101101",
			740 => "00000000000000000000101110101101",
			741 => "00000000000000000000101110101101",
			742 => "0000001010000000000101000100001000",
			743 => "0000000001000000001001011000000100",
			744 => "00000000000000000000101110101101",
			745 => "00000010001110110000101110101101",
			746 => "00000000000000000000101110101101",
			747 => "0000001100000000001001110100010000",
			748 => "0000000101000000000111111100001100",
			749 => "0000001010000000000110011100000100",
			750 => "11111110101000000000110000111001",
			751 => "0000001010000000000110011100000100",
			752 => "00000000000000000000110000111001",
			753 => "11111111101011110000110000111001",
			754 => "00000000000000000000110000111001",
			755 => "0000001001000000001010100100010100",
			756 => "0000000010000000001100001100001100",
			757 => "0000000011000000001000000100001000",
			758 => "0000000110000000000100111100000100",
			759 => "00000000000000000000110000111001",
			760 => "11111111010101100000110000111001",
			761 => "00000000000000000000110000111001",
			762 => "0000001101000000001110110100000100",
			763 => "00000000010010010000110000111001",
			764 => "00000000000000000000110000111001",
			765 => "0000001101000000000110111100001100",
			766 => "0000000011000000000010111000001000",
			767 => "0000000001000000001100011000000100",
			768 => "00000000000000000000110000111001",
			769 => "00000001001110100000110000111001",
			770 => "00000000000000000000110000111001",
			771 => "0000000111000000000100010000001100",
			772 => "0000000011000000001100001100000100",
			773 => "00000000000000000000110000111001",
			774 => "0000001000000000000001010100000100",
			775 => "11111111001011010000110000111001",
			776 => "00000000000000000000110000111001",
			777 => "0000000110000000000100101100001000",
			778 => "0000001110000000001110000000000100",
			779 => "00000000000000000000110000111001",
			780 => "00000001001010000000110000111001",
			781 => "11111111101010100000110000111001",
			782 => "0000000010000000000011000000001100",
			783 => "0000000000000000000001110100000100",
			784 => "00000000000000000000110010110101",
			785 => "0000000101000000000111111100000100",
			786 => "11111111011101110000110010110101",
			787 => "00000000000000000000110010110101",
			788 => "0000001110000000000110111000011000",
			789 => "0000001100000000000001011000010100",
			790 => "0000000000000000000111111000010000",
			791 => "0000000010000000000010010100000100",
			792 => "00000000000000000000110010110101",
			793 => "0000000001000000000101011100000100",
			794 => "00000000000000000000110010110101",
			795 => "0000001100000000001010111000000100",
			796 => "00000000000000000000110010110101",
			797 => "00000000100000110000110010110101",
			798 => "00000000000000000000110010110101",
			799 => "00000000000000000000110010110101",
			800 => "0000000001000000001101011000010000",
			801 => "0000001001000000000011101000000100",
			802 => "00000000000000000000110010110101",
			803 => "0000001111000000001000011100000100",
			804 => "00000000000000000000110010110101",
			805 => "0000000000000000000111000000000100",
			806 => "11111111011100000000110010110101",
			807 => "00000000000000000000110010110101",
			808 => "0000000000000000000011010000001000",
			809 => "0000000000000000001010101100000100",
			810 => "00000000000000000000110010110101",
			811 => "00000000001101000000110010110101",
			812 => "00000000000000000000110010110101",
			813 => "0000000001000000000101011100000100",
			814 => "11111110101110110000110100100001",
			815 => "0000000110000000000101010000100100",
			816 => "0000001001000000000011101000011000",
			817 => "0000001001000000001010100100010000",
			818 => "0000000000000000000010011000001100",
			819 => "0000000110000000000100111100000100",
			820 => "00000000000000000000110100100001",
			821 => "0000000011000000001000000100000100",
			822 => "11111111011011000000110100100001",
			823 => "00000000000000000000110100100001",
			824 => "00000000110001100000110100100001",
			825 => "0000000101000000000010011100000100",
			826 => "00000000000000000000110100100001",
			827 => "00000001000111100000110100100001",
			828 => "0000001010000000001000010100001000",
			829 => "0000000011000000000101000000000100",
			830 => "00000000000000000000110100100001",
			831 => "11111110110101000000110100100001",
			832 => "00000000101111010000110100100001",
			833 => "0000000111000000001111011100000100",
			834 => "00000000000000000000110100100001",
			835 => "0000000001000000001101011000000100",
			836 => "11111111000101000000110100100001",
			837 => "0000001000000000000111000100000100",
			838 => "00000000010110000000110100100001",
			839 => "11111111101011100000110100100001",
			840 => "0000001001000000001010100100100100",
			841 => "0000001001000000001010100100011100",
			842 => "0000001001000000000100111100000100",
			843 => "11111110010100010000110110111101",
			844 => "0000000111000000001000011000001000",
			845 => "0000001001000000001000010000000100",
			846 => "11111111010000110000110110111101",
			847 => "11111110010110100000110110111101",
			848 => "0000001110000000001111101000001100",
			849 => "0000000110000000001000010000000100",
			850 => "11111110011000000000110110111101",
			851 => "0000000110000000000101010000000100",
			852 => "00000100001110100000110110111101",
			853 => "11111111110110000000110110111101",
			854 => "11111110011000010000110110111101",
			855 => "0000000111000000001111011100000100",
			856 => "11111110011001000000110110111101",
			857 => "00000010101001100000110110111101",
			858 => "0000000111000000000111010000010000",
			859 => "0000000101000000000111111100001100",
			860 => "0000001100000000001001110100000100",
			861 => "11111110010011100000110110111101",
			862 => "0000001011000000000101110100000100",
			863 => "00000000011000000000110110111101",
			864 => "11111110011010100000110110111101",
			865 => "00000001010111010000110110111101",
			866 => "0000001000000000000111000100011000",
			867 => "0000001010000000001010110000010000",
			868 => "0000000111000000000000011100001000",
			869 => "0000000000000000001000101100000100",
			870 => "00000010100110110000110110111101",
			871 => "00000001001001010000110110111101",
			872 => "0000000000000000000010011000000100",
			873 => "00000010101000000000110110111101",
			874 => "00000011000101010000110110111101",
			875 => "0000000000000000000011111100000100",
			876 => "00000000100000100000110110111101",
			877 => "00000010100010100000110110111101",
			878 => "11111110011101100000110110111101",
			879 => "0000001001000000000100111100000100",
			880 => "11111110111111110000111000110001",
			881 => "0000000100000000000011010100100100",
			882 => "0000000110000000000100111100001100",
			883 => "0000001001000000001010100100000100",
			884 => "00000000000000000000111000110001",
			885 => "0000001011000000000100010000000100",
			886 => "00000000000000000000111000110001",
			887 => "00000000100111100000111000110001",
			888 => "0000000001000000001101011000010000",
			889 => "0000000111000000000111110000001100",
			890 => "0000000100000000000000010100001000",
			891 => "0000001000000000000101000100000100",
			892 => "00000000000000000000111000110001",
			893 => "11111111011010100000111000110001",
			894 => "00000000000000000000111000110001",
			895 => "00000000000000000000111000110001",
			896 => "0000001000000000001001101000000100",
			897 => "00000000000010010000111000110001",
			898 => "00000000000000000000111000110001",
			899 => "0000001010000000000101000100010000",
			900 => "0000001101000000001001100000000100",
			901 => "00000001000011110000111000110001",
			902 => "0000001101000000001010000100000100",
			903 => "00000000000000000000111000110001",
			904 => "0000000001000000001010011000000100",
			905 => "00000000000000000000111000110001",
			906 => "00000000011001110000111000110001",
			907 => "00000000000000000000111000110001",
			908 => "0000000001000000001100011000101100",
			909 => "0000001001000000001010100000011000",
			910 => "0000000001000000001011111100000100",
			911 => "11111110010111100000111011000101",
			912 => "0000000111000000000001101000000100",
			913 => "11111110011000110000111011000101",
			914 => "0000001101000000001001010000000100",
			915 => "00000010100110010000111011000101",
			916 => "0000001110000000001011101100001000",
			917 => "0000001100000000001001110100000100",
			918 => "11111110011110100000111011000101",
			919 => "00000000111010000000111011000101",
			920 => "11111110011010110000111011000101",
			921 => "0000000111000000001111011100000100",
			922 => "11111110011000100000111011000101",
			923 => "0000001110000000000010010100001000",
			924 => "0000000001000000000100110100000100",
			925 => "00000010101000100000111011000101",
			926 => "00000001000111010000111011000101",
			927 => "0000000110000000000101010000000100",
			928 => "00000000000000000000111011000101",
			929 => "11111110010111100000111011000101",
			930 => "0000001101000000000011001000000100",
			931 => "11111110011101100000111011000101",
			932 => "0000001000000000000110001000010100",
			933 => "0000000111000000000111010000000100",
			934 => "00000000010011000000111011000101",
			935 => "0000001100000000000101100100001100",
			936 => "0000001011000000001110101000001000",
			937 => "0000001011000000000000110100000100",
			938 => "00000001011111000000111011000101",
			939 => "00000001110100110000111011000101",
			940 => "00000000110100110000111011000101",
			941 => "00000000010000110000111011000101",
			942 => "0000000100000000000111011100000100",
			943 => "11111110110000100000111011000101",
			944 => "00000000101100010000111011000101",
			945 => "0000001001000000000100111100000100",
			946 => "11111110101100100000111101001001",
			947 => "0000001100000000000001101000011100",
			948 => "0000001010000000000001010000001100",
			949 => "0000000101000000000111111100001000",
			950 => "0000001000000000000101000100000100",
			951 => "00000000000000000000111101001001",
			952 => "11111111000010000000111101001001",
			953 => "00000000000000000000111101001001",
			954 => "0000000010000000000011110000001000",
			955 => "0000000100000000001111100000000100",
			956 => "00000000000000000000111101001001",
			957 => "00000000100100110000111101001001",
			958 => "0000001000000000001011010100000100",
			959 => "00000000000000000000111101001001",
			960 => "11111111110010110000111101001001",
			961 => "0000000100000000001100001100001000",
			962 => "0000001001000000001010100100000100",
			963 => "00000000000000000000111101001001",
			964 => "00000001000000100000111101001001",
			965 => "0000000010000000001000110100001100",
			966 => "0000000111000000001011011100000100",
			967 => "00000000000000000000111101001001",
			968 => "0000000001000000001101011000000100",
			969 => "11111111001100000000111101001001",
			970 => "00000000000000000000111101001001",
			971 => "0000001000000000000111000100001100",
			972 => "0000000000000000001010101100000100",
			973 => "00000000000000000000111101001001",
			974 => "0000000001000000000100110100000100",
			975 => "00000000000000000000111101001001",
			976 => "00000000111110010000111101001001",
			977 => "11111111110000000000111101001001",
			978 => "0000000001000000001100011000110100",
			979 => "0000001001000000001010100100101100",
			980 => "0000001001000000001010100100100000",
			981 => "0000000001000000000101011100000100",
			982 => "11111110001111010000111111100101",
			983 => "0000001100000000001001110100001100",
			984 => "0000001001000000001000010000000100",
			985 => "11111111101001000000111111100101",
			986 => "0000001001000000001001111100000100",
			987 => "11111110100010000000111111100101",
			988 => "11111110010000110000111111100101",
			989 => "0000001110000000001011101100001000",
			990 => "0000000010000000001000000100000100",
			991 => "11111110011000000000111111100101",
			992 => "00000100011111110000111111100101",
			993 => "0000001001000000001010100000000100",
			994 => "11111110010101110000111111100101",
			995 => "11111111010111100000111111100101",
			996 => "0000001100000000000001101000001000",
			997 => "0000000101000000001001010000000100",
			998 => "11111110010000110000111111100101",
			999 => "00000000011010100000111111100101",
			1000 => "00000100111110000000111111100101",
			1001 => "0000000110000000001000010000000100",
			1002 => "00000110010111000000111111100101",
			1003 => "11111110011000110000111111100101",
			1004 => "0000000101000000000111111100001000",
			1005 => "0000000111000000000111010000000100",
			1006 => "11111110010001000000111111100101",
			1007 => "00000100000000100000111111100101",
			1008 => "0000001000000000001111001000001100",
			1009 => "0000001000000000000110001000001000",
			1010 => "0000001001000000001010100100000100",
			1011 => "00000101010111110000111111100101",
			1012 => "00000110001110110000111111100101",
			1013 => "00000100011100100000111111100101",
			1014 => "0000000111000000000101110100000100",
			1015 => "11111110011000000000111111100101",
			1016 => "00000001000110000000111111100101",
			1017 => "0000000010000000000011000000001000",
			1018 => "0000001100000000001001110100000100",
			1019 => "11111111010111100001000001111001",
			1020 => "00000000000000000001000001111001",
			1021 => "0000000101000000000110010000100100",
			1022 => "0000000001000000001100011000011000",
			1023 => "0000000100000000001001000000010000",
			1024 => "0000001111000000001000001000001100",
			1025 => "0000000000000000001010101100000100",
			1026 => "00000000000000000001000001111001",
			1027 => "0000001111000000000010010100000100",
			1028 => "00000000000000000001000001111001",
			1029 => "11111111110000000001000001111001",
			1030 => "00000000000000000001000001111001",
			1031 => "0000000000000000000111111000000100",
			1032 => "00000000011010100001000001111001",
			1033 => "00000000000000000001000001111001",
			1034 => "0000001110000000000011110000001000",
			1035 => "0000001100000000001001110100000100",
			1036 => "00000000000000000001000001111001",
			1037 => "00000000110010100001000001111001",
			1038 => "00000000000000000001000001111001",
			1039 => "0000001100000000000111010000010100",
			1040 => "0000001001000000000011101000000100",
			1041 => "00000000000000000001000001111001",
			1042 => "0000000011000000000101000000000100",
			1043 => "00000000000000000001000001111001",
			1044 => "0000000111000000000101110100001000",
			1045 => "0000001101000000000110111100000100",
			1046 => "00000000000000000001000001111001",
			1047 => "11111111001111000001000001111001",
			1048 => "00000000000000000001000001111001",
			1049 => "0000000110000000000100101100001000",
			1050 => "0000001110000000001110000000000100",
			1051 => "00000000000000000001000001111001",
			1052 => "00000000101101100001000001111001",
			1053 => "00000000000000000001000001111001",
			1054 => "0000001001000000000100101100000100",
			1055 => "11111110111101100001000011101101",
			1056 => "0000000100000000000011110000100000",
			1057 => "0000000111000000001011011100010100",
			1058 => "0000000001000000001010011000010000",
			1059 => "0000000110000000000100111100000100",
			1060 => "00000000000000000001000011101101",
			1061 => "0000001011000000001110101100001000",
			1062 => "0000001010000000001000100100000100",
			1063 => "00000000000000000001000011101101",
			1064 => "11111110111011100001000011101101",
			1065 => "00000000000000000001000011101101",
			1066 => "00000000000000000001000011101101",
			1067 => "0000001101000000001111010100001000",
			1068 => "0000000000000000000111000000000100",
			1069 => "00000000101001110001000011101101",
			1070 => "00000000000000000001000011101101",
			1071 => "00000000000000000001000011101101",
			1072 => "0000000110000000000100101100010100",
			1073 => "0000001100000000001011011100010000",
			1074 => "0000001100000000001001110100000100",
			1075 => "00000000000000000001000011101101",
			1076 => "0000001110000000000110001100001000",
			1077 => "0000000111000000001000011000000100",
			1078 => "00000000000000000001000011101101",
			1079 => "00000000110001010001000011101101",
			1080 => "00000000000000000001000011101101",
			1081 => "00000000000000000001000011101101",
			1082 => "11111111110101100001000011101101",
			1083 => "0000000010000000000011000000001100",
			1084 => "0000001000000000000101000100000100",
			1085 => "00000000000000000001000101110001",
			1086 => "0000001100000000000001101000000100",
			1087 => "11111111011001010001000101110001",
			1088 => "00000000000000000001000101110001",
			1089 => "0000000110000000000100101100110100",
			1090 => "0000000000000000000111000000011000",
			1091 => "0000001000000000000001010100001000",
			1092 => "0000001001000000001010100100000100",
			1093 => "00000000000000000001000101110001",
			1094 => "00000000010001100001000101110001",
			1095 => "0000001001000000000011101000000100",
			1096 => "00000000000000000001000101110001",
			1097 => "0000000011000000001110100100000100",
			1098 => "00000000000000000001000101110001",
			1099 => "0000001001000000000011101000000100",
			1100 => "11111111010001110001000101110001",
			1101 => "00000000000000000001000101110001",
			1102 => "0000001001000000000010101100010100",
			1103 => "0000000100000000001001000000001100",
			1104 => "0000001111000000001000001000001000",
			1105 => "0000001111000000000010010100000100",
			1106 => "00000000000000000001000101110001",
			1107 => "11111111110110100001000101110001",
			1108 => "00000000000000000001000101110001",
			1109 => "0000000100000000000000101100000100",
			1110 => "00000000001100110001000101110001",
			1111 => "00000000000000000001000101110001",
			1112 => "0000001100000000001000011000000100",
			1113 => "00000000000000000001000101110001",
			1114 => "00000000110010000001000101110001",
			1115 => "11111111110101100001000101110001",
			1116 => "0000001001000000000111101100001000",
			1117 => "0000000100000000000000100000000100",
			1118 => "11111110100101100001001000010101",
			1119 => "00000000000000000001001000010101",
			1120 => "0000001110000000001000011100110100",
			1121 => "0000000100000000000110001100100000",
			1122 => "0000000110000000001000010000010000",
			1123 => "0000000101000000000111111100001000",
			1124 => "0000000110000000001111000000000100",
			1125 => "00000000000000000001001000010101",
			1126 => "11111111001111000001001000010101",
			1127 => "0000000100000000000110001100000100",
			1128 => "00000001000110010001001000010101",
			1129 => "00000000000000000001001000010101",
			1130 => "0000000111000000000100010000001100",
			1131 => "0000000100000000001100001100001000",
			1132 => "0000001100000000001010001100000100",
			1133 => "11111111000110100001001000010101",
			1134 => "00000000000000000001001000010101",
			1135 => "00000000000000000001001000010101",
			1136 => "00000000000000000001001000010101",
			1137 => "0000000110000000000101010000001100",
			1138 => "0000001011000000000100010000000100",
			1139 => "00000000000000000001001000010101",
			1140 => "0000001100000000000001011000000100",
			1141 => "00000001000110000001001000010101",
			1142 => "00000000000000000001001000010101",
			1143 => "0000001100000000000111010000000100",
			1144 => "00000000000000000001001000010101",
			1145 => "11111111110010110001001000010101",
			1146 => "0000001001000000000111110100001100",
			1147 => "0000000111000000000100010000001000",
			1148 => "0000001100000000000111010000000100",
			1149 => "11111110111001110001001000010101",
			1150 => "00000000000000000001001000010101",
			1151 => "00000000000000000001001000010101",
			1152 => "0000000110000000000100101100001000",
			1153 => "0000001100000000001111011100000100",
			1154 => "00000000000000000001001000010101",
			1155 => "00000000111001010001001000010101",
			1156 => "11111111100111010001001000010101",
			1157 => "0000001001000000001010100100011100",
			1158 => "0000000010000000001101101100000100",
			1159 => "11111110011000110001001011001001",
			1160 => "0000001110000000001111101000010100",
			1161 => "0000001100000000000100011000000100",
			1162 => "11111110100001100001001011001001",
			1163 => "0000000111000000001001001000000100",
			1164 => "00000011110101100001001011001001",
			1165 => "0000001001000000000101010000000100",
			1166 => "11111110011111100001001011001001",
			1167 => "0000000110000000000101010000000100",
			1168 => "00000001001110100001001011001001",
			1169 => "11111111010011100001001011001001",
			1170 => "11111110011010100001001011001001",
			1171 => "0000000101000000000111111100010100",
			1172 => "0000000100000000001000001000001000",
			1173 => "0000001000000000000101000100000100",
			1174 => "00000000000010100001001011001001",
			1175 => "11111110001101000001001011001001",
			1176 => "0000000100000000000011001100000100",
			1177 => "00001001100111000001001011001001",
			1178 => "0000001111000000001100001100000100",
			1179 => "00000001100110110001001011001001",
			1180 => "11111110111001110001001011001001",
			1181 => "0000000110000000001001111100011100",
			1182 => "0000001001000000001010100100001000",
			1183 => "0000001010000000001001000100000100",
			1184 => "00000001100100100001001011001001",
			1185 => "11111111011000110001001011001001",
			1186 => "0000001101000000001010000100001100",
			1187 => "0000001101000000000110111100000100",
			1188 => "00000001101001110001001011001001",
			1189 => "0000000111000000001011011100000100",
			1190 => "11111111000100000001001011001001",
			1191 => "00000001011011010001001011001001",
			1192 => "0000000000000000000111000000000100",
			1193 => "11111110111011010001001011001001",
			1194 => "00000001100011000001001011001001",
			1195 => "0000000100000000000000010100000100",
			1196 => "11111110110001100001001011001001",
			1197 => "0000001000000000000111000100001000",
			1198 => "0000001100000000001111011100000100",
			1199 => "11111111110100000001001011001001",
			1200 => "00000001111011000001001011001001",
			1201 => "11111110110000100001001011001001",
			1202 => "0000001100000000001011000000000100",
			1203 => "11111111010111010001001101001101",
			1204 => "0000000110000000001001111100101100",
			1205 => "0000000100000000000011110000011100",
			1206 => "0000001011000000000000110100010000",
			1207 => "0000000110000000000100111100000100",
			1208 => "00000000000000000001001101001101",
			1209 => "0000000001000000001010011000001000",
			1210 => "0000000111000000001011011100000100",
			1211 => "11111111001111010001001101001101",
			1212 => "00000000000000000001001101001101",
			1213 => "00000000000000000001001101001101",
			1214 => "0000001011000000000110100000001000",
			1215 => "0000000001000000000100110100000100",
			1216 => "00000000000000000001001101001101",
			1217 => "00000000011011100001001101001101",
			1218 => "00000000000000000001001101001101",
			1219 => "0000001001000000000100101100000100",
			1220 => "00000000000000000001001101001101",
			1221 => "0000000010000000001101001000001000",
			1222 => "0000000111000000001000011000000100",
			1223 => "00000000000000000001001101001101",
			1224 => "00000000101101100001001101001101",
			1225 => "00000000000000000001001101001101",
			1226 => "0000001110000000000011010100010000",
			1227 => "0000000001000000000100111100001100",
			1228 => "0000000010000000000110001100000100",
			1229 => "00000000000000000001001101001101",
			1230 => "0000001010000000001010110000000100",
			1231 => "00000000000000000001001101001101",
			1232 => "11111111010010000001001101001101",
			1233 => "00000000000000000001001101001101",
			1234 => "00000000000000000001001101001101",
			1235 => "0000000001000000000111101000001000",
			1236 => "0000000100000000000000100000000100",
			1237 => "11111110100100000001001111111001",
			1238 => "00000000000000000001001111111001",
			1239 => "0000000000000000000111000000100100",
			1240 => "0000001111000000001000011100010100",
			1241 => "0000000111000000000001011000010000",
			1242 => "0000001000000000000101000100000100",
			1243 => "00000000000000000001001111111001",
			1244 => "0000000100000000001110100100001000",
			1245 => "0000001011000000000000110100000100",
			1246 => "11111110111011110001001111111001",
			1247 => "00000000000000000001001111111001",
			1248 => "00000000000000000001001111111001",
			1249 => "00000001000001110001001111111001",
			1250 => "0000000001000000001010011000001000",
			1251 => "0000000101000000000010000000000100",
			1252 => "00000000000000000001001111111001",
			1253 => "00000000001000000001001111111001",
			1254 => "0000001101000000000110111100000100",
			1255 => "00000000000000000001001111111001",
			1256 => "11111110101110000001001111111001",
			1257 => "0000000110000000000101010000010000",
			1258 => "0000001011000000000100010000000100",
			1259 => "00000000000000000001001111111001",
			1260 => "0000000100000000000011110000000100",
			1261 => "00000000000000000001001111111001",
			1262 => "0000000101000000001100010000000100",
			1263 => "00000001001100110001001111111001",
			1264 => "00000000000000000001001111111001",
			1265 => "0000000100000000000000010100001100",
			1266 => "0000001010000000000110011000000100",
			1267 => "00000000000000000001001111111001",
			1268 => "0000000001000000001001100100000100",
			1269 => "11111110111110110001001111111001",
			1270 => "00000000000000000001001111111001",
			1271 => "0000000000000000000011010000001000",
			1272 => "0000001000000000001011010100000100",
			1273 => "00000000000000000001001111111001",
			1274 => "00000000110000000001001111111001",
			1275 => "0000000100000000001011001000000100",
			1276 => "11111111001011010001001111111001",
			1277 => "00000000000100100001001111111001",
			1278 => "0000001100000000001011000000000100",
			1279 => "11111111010010010001010001111101",
			1280 => "0000001110000000000110111000011000",
			1281 => "0000000010000000000010010100000100",
			1282 => "00000000000000000001010001111101",
			1283 => "0000001000000000000111000100010000",
			1284 => "0000000001000000001011111100000100",
			1285 => "00000000000000000001010001111101",
			1286 => "0000001100000000000111010000001000",
			1287 => "0000001010000000001000100100000100",
			1288 => "00000000000000000001010001111101",
			1289 => "00000000110000010001010001111101",
			1290 => "00000000000000000001010001111101",
			1291 => "00000000000000000001010001111101",
			1292 => "0000001100000000001010001100010100",
			1293 => "0000001000000000000001010100000100",
			1294 => "00000000000000000001010001111101",
			1295 => "0000001001000000000111110100001100",
			1296 => "0000000111000000000101110100001000",
			1297 => "0000000001000000000100110100000100",
			1298 => "00000000000000000001010001111101",
			1299 => "11111111010101110001010001111101",
			1300 => "00000000000000000001010001111101",
			1301 => "00000000000000000001010001111101",
			1302 => "0000001000000000000110001000001100",
			1303 => "0000000111000000001011110100001000",
			1304 => "0000000001000000001100011000000100",
			1305 => "00000000000000000001010001111101",
			1306 => "00000000100110010001010001111101",
			1307 => "00000000000000000001010001111101",
			1308 => "0000000001000000001001100100000100",
			1309 => "11111111101101010001010001111101",
			1310 => "00000000000000000001010001111101",
			1311 => "0000000001000000000100110100100000",
			1312 => "0000000110000000000100111100000100",
			1313 => "11111110011001010001010101010001",
			1314 => "0000001111000000000110111000010000",
			1315 => "0000000100000000000111011100001000",
			1316 => "0000001111000000000110111000000100",
			1317 => "11111110110010010001010101010001",
			1318 => "00000000000000000001010101010001",
			1319 => "0000000001000000001101011100000100",
			1320 => "11111111100010100001010101010001",
			1321 => "00000010000110010001010101010001",
			1322 => "0000000110000000001000010000001000",
			1323 => "0000000010000000001000011100000100",
			1324 => "11111111011010100001010101010001",
			1325 => "00000000100110010001010101010001",
			1326 => "11111110100011100001010101010001",
			1327 => "0000000001000000001100011000101000",
			1328 => "0000000110000000000100111100010100",
			1329 => "0000000011000000000001011100000100",
			1330 => "11111110110010100001010101010001",
			1331 => "0000000100000000000011110000001100",
			1332 => "0000000100000000001110100100000100",
			1333 => "00000001011111000001010101010001",
			1334 => "0000000100000000000101000000000100",
			1335 => "11111111110101010001010101010001",
			1336 => "00000000101001010001010101010001",
			1337 => "00000011011010100001010101010001",
			1338 => "0000000100000000001110111000010000",
			1339 => "0000001110000000001000101000001000",
			1340 => "0000001011000000000010001000000100",
			1341 => "11111111110111000001010101010001",
			1342 => "00000000110111100001010101010001",
			1343 => "0000000100000000001000011100000100",
			1344 => "00000000000000000001010101010001",
			1345 => "11111101101101000001010101010001",
			1346 => "00000000111111010001010101010001",
			1347 => "0000001000000000000110001000011100",
			1348 => "0000001101000000001010000100010100",
			1349 => "0000000111000000000111010000001100",
			1350 => "0000001110000000000110111000001000",
			1351 => "0000000010000000001011110000000100",
			1352 => "00000000000000000001010101010001",
			1353 => "00000001001100000001010101010001",
			1354 => "11111110110100100001010101010001",
			1355 => "0000000111000000000111110000000100",
			1356 => "00000001100101000001010101010001",
			1357 => "00000000000000000001010101010001",
			1358 => "0000001110000000001110100100000100",
			1359 => "11111110011001000001010101010001",
			1360 => "00000001100100110001010101010001",
			1361 => "0000000111000000000101110100000100",
			1362 => "11111110101100010001010101010001",
			1363 => "00000000000000000001010101010001",
			1364 => "0000001001000000001010100000100100",
			1365 => "0000000110000000000100111100000100",
			1366 => "11111110011010000001011000101101",
			1367 => "0000001111000000000010010100001100",
			1368 => "0000001001000000001011001100000100",
			1369 => "11111111011001110001011000101101",
			1370 => "0000000100000000001010110100000100",
			1371 => "00000000000000000001011000101101",
			1372 => "00000001110010000001011000101101",
			1373 => "0000000001000000000111101000000100",
			1374 => "11111110100000100001011000101101",
			1375 => "0000000001000000000001111000001000",
			1376 => "0000000110000000000101010000000100",
			1377 => "00000001000011010001011000101101",
			1378 => "00000000000000000001011000101101",
			1379 => "0000000110000000000101010000000100",
			1380 => "00000000000000000001011000101101",
			1381 => "11111110111011000001011000101101",
			1382 => "0000000001000000001100011000101000",
			1383 => "0000000001000000000100110100010100",
			1384 => "0000000100000000001000001000001000",
			1385 => "0000000110000000000100111100000100",
			1386 => "00000000000000000001011000101101",
			1387 => "11111111001011000001011000101101",
			1388 => "0000000101000000000011001000001000",
			1389 => "0000001011000000000100010000000100",
			1390 => "00000000000000000001011000101101",
			1391 => "00000001110100010001011000101101",
			1392 => "11111111101000100001011000101101",
			1393 => "0000001000000000000101000100001000",
			1394 => "0000000011000000000001011100000100",
			1395 => "00000000000000000001011000101101",
			1396 => "00000000110110000001011000101101",
			1397 => "0000000000000000000010111100001000",
			1398 => "0000001001000000000010101100000100",
			1399 => "11111110100010100001011000101101",
			1400 => "00000000000000000001011000101101",
			1401 => "00000000000000000001011000101101",
			1402 => "0000000101000000000111111100001000",
			1403 => "0000001110000000001101101100000100",
			1404 => "00000000000110110001011000101101",
			1405 => "11111110100100000001011000101101",
			1406 => "0000001101000000000110111100001000",
			1407 => "0000001110000000000011110000000100",
			1408 => "00000001100100010001011000101101",
			1409 => "00000000000000000001011000101101",
			1410 => "0000000111000000001011011100000100",
			1411 => "11111101111110100001011000101101",
			1412 => "0000000000000000001010101100001000",
			1413 => "0000001001000000000011101000000100",
			1414 => "00000001000111010001011000101101",
			1415 => "11111111000011110001011000101101",
			1416 => "0000001000000000000111000100000100",
			1417 => "00000001010010010001011000101101",
			1418 => "11111111000011100001011000101101",
			1419 => "0000000001000000000001111000001100",
			1420 => "0000000001000000000101011100000100",
			1421 => "11111110011010010001011011100001",
			1422 => "0000000100000000000111011100000100",
			1423 => "11111110101000110001011011100001",
			1424 => "00000000011110000001011011100001",
			1425 => "0000000001000000001101011000111100",
			1426 => "0000001111000000001000011100011100",
			1427 => "0000001101000000001010001000001000",
			1428 => "0000001000000000001011010100000100",
			1429 => "11111110110001100001011011100001",
			1430 => "00000000000000000001011011100001",
			1431 => "0000001100000000000001011000010000",
			1432 => "0000001111000000001111101000001000",
			1433 => "0000001100000000001001110100000100",
			1434 => "11111110101000110001011011100001",
			1435 => "00000000111100110001011011100001",
			1436 => "0000001111000000001000110100000100",
			1437 => "00000001011100010001011011100001",
			1438 => "00000000011110000001011011100001",
			1439 => "11111111010101000001011011100001",
			1440 => "0000000111000000000110110100010100",
			1441 => "0000000100000000000100001100010000",
			1442 => "0000001111000000001000011100001000",
			1443 => "0000000010000000001000110100000100",
			1444 => "11111001100111010001011011100001",
			1445 => "00000000000000000001011011100001",
			1446 => "0000001011000000000010110100000100",
			1447 => "11111101110111110001011011100001",
			1448 => "00000000000000000001011011100001",
			1449 => "00000000011001100001011011100001",
			1450 => "0000000110000000001001111100001000",
			1451 => "0000000001000000000100110100000100",
			1452 => "00000000000000000001011011100001",
			1453 => "00000001011001110001011011100001",
			1454 => "11111110111000010001011011100001",
			1455 => "0000001010000000001000010100001000",
			1456 => "0000000011000000001110100100000100",
			1457 => "00000001010010000001011011100001",
			1458 => "11111110101101000001011011100001",
			1459 => "0000000110000000000100101100001000",
			1460 => "0000001011000000000001001000000100",
			1461 => "00000000000000000001011011100001",
			1462 => "00000001100101100001011011100001",
			1463 => "00000000001011100001011011100001",
			1464 => "0000001001000000000100111100000100",
			1465 => "11111111000010010001011101101101",
			1466 => "0000000100000000000011010100110000",
			1467 => "0000000110000000000100111100001100",
			1468 => "0000001001000000001010100100000100",
			1469 => "00000000000000000001011101101101",
			1470 => "0000001011000000000100010000000100",
			1471 => "00000000000000000001011101101101",
			1472 => "00000000100100010001011101101101",
			1473 => "0000000001000000001100011000001000",
			1474 => "0000001111000000000010010100000100",
			1475 => "00000000000000000001011101101101",
			1476 => "11111111001010110001011101101101",
			1477 => "0000001011000000000110100000010000",
			1478 => "0000001000000000000101000100001000",
			1479 => "0000000111000000001011011100000100",
			1480 => "11111111100111110001011101101101",
			1481 => "00000000000000000001011101101101",
			1482 => "0000000010000000000011110000000100",
			1483 => "00000000110000000001011101101101",
			1484 => "00000000000000000001011101101101",
			1485 => "0000001001000000000011101000000100",
			1486 => "00000000000000000001011101101101",
			1487 => "0000001111000000001000011100000100",
			1488 => "00000000000000000001011101101101",
			1489 => "11111111011011110001011101101101",
			1490 => "0000001010000000000101000100010000",
			1491 => "0000001101000000001001100000000100",
			1492 => "00000001000000110001011101101101",
			1493 => "0000001101000000001010000100000100",
			1494 => "00000000000000000001011101101101",
			1495 => "0000001001000000000011101000000100",
			1496 => "00000000000000000001011101101101",
			1497 => "00000000011000100001011101101101",
			1498 => "00000000000000000001011101101101",
			1499 => "0000001100000000001010111000000100",
			1500 => "11111110100011010001011111110001",
			1501 => "0000000100000000001011001000111000",
			1502 => "0000000110000000000101010000101000",
			1503 => "0000000100000000000011110000011000",
			1504 => "0000001000000000000001010100001100",
			1505 => "0000001011000000001011110100000100",
			1506 => "00000000000000000001011111110001",
			1507 => "0000000100000000000110001100000100",
			1508 => "00000001000101100001011111110001",
			1509 => "00000000000000000001011111110001",
			1510 => "0000000001000000001101011000001000",
			1511 => "0000001100000000001010001100000100",
			1512 => "11111111000100010001011111110001",
			1513 => "00000000000000000001011111110001",
			1514 => "00000000010010100001011111110001",
			1515 => "0000001100000000001000000000000100",
			1516 => "11111111101111000001011111110001",
			1517 => "0000001111000000000011001100001000",
			1518 => "0000000001000000001011111100000100",
			1519 => "00000000000000000001011111110001",
			1520 => "00000001010000000001011111110001",
			1521 => "00000000000000000001011111110001",
			1522 => "0000000001000000001101011000001000",
			1523 => "0000000100000000000011101100000100",
			1524 => "11111110111001110001011111110001",
			1525 => "00000000000000000001011111110001",
			1526 => "0000001000000000001111001000000100",
			1527 => "00000000100101110001011111110001",
			1528 => "11111111101010010001011111110001",
			1529 => "0000001010000000000101000100000100",
			1530 => "00000001101000010001011111110001",
			1531 => "11111111111101000001011111110001",
			1532 => "0000000001000000000100110101000000",
			1533 => "0000000001000000000100110100110000",
			1534 => "0000000001000000000101011100000100",
			1535 => "11111110010101000001100010100101",
			1536 => "0000001100000000001001110100010100",
			1537 => "0000000001000000000101011100001000",
			1538 => "0000000111000000000110100100000100",
			1539 => "00000001101001000001100010100101",
			1540 => "11111110100011100001100010100101",
			1541 => "0000001100000000001000000000000100",
			1542 => "11111110010101110001100010100101",
			1543 => "0000000001000000001110010100000100",
			1544 => "00000000000000000001100010100101",
			1545 => "11111110010110110001100010100101",
			1546 => "0000000111000000000111010000001100",
			1547 => "0000000110000000001000010000000100",
			1548 => "11111110100011010001100010100101",
			1549 => "0000000011000000000110111000000100",
			1550 => "00000011010001010001100010100101",
			1551 => "11111110110100000001100010100101",
			1552 => "0000001100000000000001101000001000",
			1553 => "0000000001000000000111101000000100",
			1554 => "11111110100000100001100010100101",
			1555 => "00000001101001010001100010100101",
			1556 => "11111110010101000001100010100101",
			1557 => "0000000111000000000111010000001000",
			1558 => "0000001100000000001001110100000100",
			1559 => "11111110010110100001100010100101",
			1560 => "00000000000000000001100010100101",
			1561 => "0000000011000000001110000000000100",
			1562 => "00000011100110100001100010100101",
			1563 => "00000000110011110001100010100101",
			1564 => "0000001101000000001100010100000100",
			1565 => "11111110010011000001100010100101",
			1566 => "0000000110000000000100101100010100",
			1567 => "0000000100000000001001000000010000",
			1568 => "0000001000000000000110001000001100",
			1569 => "0000000101000000000111111100000100",
			1570 => "00000001000000010001100010100101",
			1571 => "0000000001000000001100011000000100",
			1572 => "00000010001100110001100010100101",
			1573 => "00000010011001100001100010100101",
			1574 => "11111111000000100001100010100101",
			1575 => "00000100010111000001100010100101",
			1576 => "11111110011010110001100010100101",
			1577 => "0000000010000000001101101100001000",
			1578 => "0000000011000000000001011100000100",
			1579 => "11111110011011010001100101001001",
			1580 => "00000000000000000001100101001001",
			1581 => "0000001111000000001000000100011000",
			1582 => "0000001100000000001010111000000100",
			1583 => "11111111011111010001100101001001",
			1584 => "0000001100000000000001011000010000",
			1585 => "0000001001000000001011001100000100",
			1586 => "00000000000000000001100101001001",
			1587 => "0000000100000000000110111000000100",
			1588 => "00000000000000000001100101001001",
			1589 => "0000000110000000001111000000000100",
			1590 => "00000000000000000001100101001001",
			1591 => "00000001010001110001100101001001",
			1592 => "11111111110011100001100101001001",
			1593 => "0000000001000000001101011000101000",
			1594 => "0000001011000000000110100000011100",
			1595 => "0000000111000000001011011100010000",
			1596 => "0000000101000000000011001000001000",
			1597 => "0000000110000000001001111100000100",
			1598 => "00000000001110000001100101001001",
			1599 => "11111111001000110001100101001001",
			1600 => "0000000001000000001101011000000100",
			1601 => "11111110011100000001100101001001",
			1602 => "00000000000000000001100101001001",
			1603 => "0000000001000000001100011000001000",
			1604 => "0000001100000000001111011100000100",
			1605 => "00000000000000000001100101001001",
			1606 => "11111111011001110001100101001001",
			1607 => "00000001010011110001100101001001",
			1608 => "0000001001000000000011101000001000",
			1609 => "0000000100000000001101001000000100",
			1610 => "00000000110100000001100101001001",
			1611 => "11111110111101110001100101001001",
			1612 => "11111101110010100001100101001001",
			1613 => "0000001010000000000110011100001000",
			1614 => "0000000111000000000000011100000100",
			1615 => "00000000000000000001100101001001",
			1616 => "00000001011100010001100101001001",
			1617 => "00000000000000000001100101001001",
			1618 => "0000000010000000001100111000000100",
			1619 => "11111110100001100001100111010101",
			1620 => "0000000100000000001011001000111000",
			1621 => "0000000110000000000101010000101100",
			1622 => "0000000100000000000011110000011100",
			1623 => "0000000000000000001010101100001100",
			1624 => "0000000111000000000111010000000100",
			1625 => "00000000000000000001100111010101",
			1626 => "0000000001000000000100110100000100",
			1627 => "00000000000000000001100111010101",
			1628 => "00000001001000000001100111010101",
			1629 => "0000000111000000000110110100001000",
			1630 => "0000000001000000001101011000000100",
			1631 => "11111110110100100001100111010101",
			1632 => "00000000000000000001100111010101",
			1633 => "0000000111000000000101110100000100",
			1634 => "00000000101101010001100111010101",
			1635 => "00000000000000000001100111010101",
			1636 => "0000001100000000001000000000000100",
			1637 => "11111111100110110001100111010101",
			1638 => "0000001110000000000110001100001000",
			1639 => "0000000001000000001011111100000100",
			1640 => "00000000000000000001100111010101",
			1641 => "00000001010011100001100111010101",
			1642 => "00000000000000000001100111010101",
			1643 => "0000000001000000001101011000000100",
			1644 => "11111110111001010001100111010101",
			1645 => "0000001000000000001111001000000100",
			1646 => "00000000101011000001100111010101",
			1647 => "11111111100011100001100111010101",
			1648 => "0000001010000000000101000100001000",
			1649 => "0000000110000000001000010000000100",
			1650 => "00000000000000000001100111010101",
			1651 => "00000001110000110001100111010101",
			1652 => "11111111110010110001100111010101",
			1653 => "0000001001000000001010100000010000",
			1654 => "0000001001000000001001111100000100",
			1655 => "11111110011001110001101010100001",
			1656 => "0000000100000000000010100100000100",
			1657 => "11111110100101100001101010100001",
			1658 => "0000000110000000001001111100000100",
			1659 => "00000001100000010001101010100001",
			1660 => "11111111111011100001101010100001",
			1661 => "0000000111000000000001011000100100",
			1662 => "0000001111000000000010111000100000",
			1663 => "0000000100000000000010110000010000",
			1664 => "0000001011000000000000110100001100",
			1665 => "0000001001000000000011101000001000",
			1666 => "0000000110000000001111000000000100",
			1667 => "00000000000000000001101010100001",
			1668 => "11111110011010100001101010100001",
			1669 => "00000000010001000001101010100001",
			1670 => "00000001000011010001101010100001",
			1671 => "0000000110000000001001111100001100",
			1672 => "0000001011000000000100010000000100",
			1673 => "00000000000000000001101010100001",
			1674 => "0000000011000000000110001100000100",
			1675 => "00000001110000100001101010100001",
			1676 => "00000000000000000001101010100001",
			1677 => "11111111110001000001101010100001",
			1678 => "11111110000111100001101010100001",
			1679 => "0000000101000000000110010000001100",
			1680 => "0000001001000000001010100100001000",
			1681 => "0000001001000000001010100100000100",
			1682 => "00000000010010100001101010100001",
			1683 => "11111111111111110001101010100001",
			1684 => "00000001100110010001101010100001",
			1685 => "0000000111000000000110110100010000",
			1686 => "0000000101000000000110010000001000",
			1687 => "0000001010000000001000010100000100",
			1688 => "11111001010000110001101010100001",
			1689 => "00000000000000000001101010100001",
			1690 => "0000000101000000001110110100000100",
			1691 => "00000000110111110001101010100001",
			1692 => "00000000000000000001101010100001",
			1693 => "0000001010000000001010110000010000",
			1694 => "0000000000000000001010101100001000",
			1695 => "0000000011000000000101000000000100",
			1696 => "00000000110110110001101010100001",
			1697 => "11111110010111010001101010100001",
			1698 => "0000001001000000000010101100000100",
			1699 => "00000000000000000001101010100001",
			1700 => "00000001100010100001101010100001",
			1701 => "0000001001000000001000100100000100",
			1702 => "11111110011000110001101010100001",
			1703 => "00000000010110110001101010100001",
			1704 => "0000001001000000000100111100000100",
			1705 => "11111110111000110001101100111101",
			1706 => "0000001101000000000110010000010100",
			1707 => "0000000100000000000111011100010000",
			1708 => "0000001001000000000111101100000100",
			1709 => "11111111110100000001101100111101",
			1710 => "0000001100000000001001110100000100",
			1711 => "00000000000000000001101100111101",
			1712 => "0000001100000000000110100100000100",
			1713 => "00000000011010110001101100111101",
			1714 => "00000000000000000001101100111101",
			1715 => "00000000110101110001101100111101",
			1716 => "0000001011000000000000110100010000",
			1717 => "0000000001000000001010011000001100",
			1718 => "0000000110000000000100111100000100",
			1719 => "00000000000000000001101100111101",
			1720 => "0000001100000000001111011100000100",
			1721 => "11111110110000000001101100111101",
			1722 => "00000000000000000001101100111101",
			1723 => "00000000000000000001101100111101",
			1724 => "0000001101000000000111011000010000",
			1725 => "0000000010000000001101001000001100",
			1726 => "0000000001000000001101111100000100",
			1727 => "00000000000000000001101100111101",
			1728 => "0000001100000000000001011000000100",
			1729 => "00000000100101110001101100111101",
			1730 => "00000000000000000001101100111101",
			1731 => "00000000000000000001101100111101",
			1732 => "0000001000000000000110001000010000",
			1733 => "0000000010000000001000110100001000",
			1734 => "0000000010000000001000000100000100",
			1735 => "00000000000000000001101100111101",
			1736 => "11111111100011110001101100111101",
			1737 => "0000000000000000001010101100000100",
			1738 => "00000000000000000001101100111101",
			1739 => "00000000101001100001101100111101",
			1740 => "0000000001000000000100111100000100",
			1741 => "11111111100000010001101100111101",
			1742 => "00000000000000000001101100111101",
			1743 => "0000001100000000001011000000000100",
			1744 => "11111110011111010001101111110001",
			1745 => "0000001011000000000110100000111000",
			1746 => "0000001001000000000010101100100100",
			1747 => "0000001110000000000110111000010100",
			1748 => "0000001001000000000101010000000100",
			1749 => "11111111100001100001101111110001",
			1750 => "0000000100000000000010110000001000",
			1751 => "0000000111000000000111010000000100",
			1752 => "11111111001101000001101111110001",
			1753 => "00000000100111010001101111110001",
			1754 => "0000000110000000000101010000000100",
			1755 => "00000001010100100001101111110001",
			1756 => "00000000000000000001101111110001",
			1757 => "0000000110000000001000010000000100",
			1758 => "00000000000000000001101111110001",
			1759 => "0000000101000000000110010000001000",
			1760 => "0000000100000000000100001100000100",
			1761 => "11111110100100110001101111110001",
			1762 => "00000000000000000001101111110001",
			1763 => "00000000000000000001101111110001",
			1764 => "0000001100000000000001101000001100",
			1765 => "0000001100000000001001110100000100",
			1766 => "00000000000111100001101111110001",
			1767 => "0000000111000000000001011000000100",
			1768 => "11111111010000110001101111110001",
			1769 => "00000000000000000001101111110001",
			1770 => "0000001001000000001000010100000100",
			1771 => "00000001010110100001101111110001",
			1772 => "00000000000000000001101111110001",
			1773 => "0000001001000000000011101000011000",
			1774 => "0000001000000000000001010100001000",
			1775 => "0000001001000000000011101000000100",
			1776 => "00000000001010010001101111110001",
			1777 => "00000000000000000001101111110001",
			1778 => "0000001100000000001111011100000100",
			1779 => "00000000000000000001101111110001",
			1780 => "0000000110000000001000010000000100",
			1781 => "00000000000000000001101111110001",
			1782 => "0000001101000000000111011000000100",
			1783 => "00000000000000000001101111110001",
			1784 => "11111110101011010001101111110001",
			1785 => "0000001000000000000111000100000100",
			1786 => "00000000101101110001101111110001",
			1787 => "00000000000000000001101111110001",
			1788 => "0000000010000000000011000000001000",
			1789 => "0000001100000000001001110100000100",
			1790 => "11111110011011010001110010111101",
			1791 => "00000000000000000001110010111101",
			1792 => "0000000001000000001101011001001000",
			1793 => "0000001111000000001000000100011100",
			1794 => "0000001001000000001010100100001100",
			1795 => "0000000100000000000011110100000100",
			1796 => "11111111010100100001110010111101",
			1797 => "0000001000000000000001110100000100",
			1798 => "00000000110101010001110010111101",
			1799 => "00000000000000000001110010111101",
			1800 => "0000001111000000000010010100001000",
			1801 => "0000001100000000000001101000000100",
			1802 => "11111111100000000001110010111101",
			1803 => "00000000010110110001110010111101",
			1804 => "0000001100000000001001110100000100",
			1805 => "00000000000000000001110010111101",
			1806 => "00000001011110110001110010111101",
			1807 => "0000000010000000001000110100010000",
			1808 => "0000000101000000000110010000001100",
			1809 => "0000000000000000001010101100000100",
			1810 => "00000000000000000001110010111101",
			1811 => "0000001111000000001000110100000100",
			1812 => "00000000000000000001110010111101",
			1813 => "11111110001110000001110010111101",
			1814 => "00000000000011000001110010111101",
			1815 => "0000001010000000000110011000010000",
			1816 => "0000001001000000000011101000001000",
			1817 => "0000001001000000001010100000000100",
			1818 => "00000000000000000001110010111101",
			1819 => "00000001001011100001110010111101",
			1820 => "0000001010000000001000010100000100",
			1821 => "11111111011011100001110010111101",
			1822 => "00000000000000000001110010111101",
			1823 => "0000001101000000001100010000001000",
			1824 => "0000000001000000000100110100000100",
			1825 => "11111111000100010001110010111101",
			1826 => "00000000100010000001110010111101",
			1827 => "11111110110101110001110010111101",
			1828 => "0000001101000000001010000100001100",
			1829 => "0000000101000000000111111100000100",
			1830 => "00000000000000000001110010111101",
			1831 => "0000001111000000001001001100000100",
			1832 => "00000001011100010001110010111101",
			1833 => "00000000000000000001110010111101",
			1834 => "0000001001000000001000100100000100",
			1835 => "11111111001011110001110010111101",
			1836 => "0000001000000000000001110100000100",
			1837 => "00000001001010100001110010111101",
			1838 => "11111111100111010001110010111101",
			1839 => "0000000010000000001101101100001000",
			1840 => "0000001011000000001010010100000100",
			1841 => "11111110011001110001110110001001",
			1842 => "00000000000000000001110110001001",
			1843 => "0000000001000000001100011000110100",
			1844 => "0000000110000000000101010000101000",
			1845 => "0000000100000000001000001000010100",
			1846 => "0000001011000000000000110100001100",
			1847 => "0000000110000000000100111100001000",
			1848 => "0000000110000000001111000000000100",
			1849 => "00000000000000000001110110001001",
			1850 => "00000000000100110001110110001001",
			1851 => "11111110011000100001110110001001",
			1852 => "0000000001000000000100110100000100",
			1853 => "00000000000000000001110110001001",
			1854 => "00000001000001100001110110001001",
			1855 => "0000001001000000001011001100000100",
			1856 => "11111111001111100001110110001001",
			1857 => "0000000110000000001000010000001000",
			1858 => "0000000110000000000100111100000100",
			1859 => "00000000000000000001110110001001",
			1860 => "00000001111111010001110110001001",
			1861 => "0000000001000000000111101000000100",
			1862 => "11111111010100110001110110001001",
			1863 => "00000001000010010001110110001001",
			1864 => "0000000111000000000111010000001000",
			1865 => "0000000111000000001111011100000100",
			1866 => "11111111010000000001110110001001",
			1867 => "00000000000000000001110110001001",
			1868 => "11111110011011100001110110001001",
			1869 => "0000000101000000000111111100001100",
			1870 => "0000000001000000001010011000001000",
			1871 => "0000000100000000000011001100000100",
			1872 => "00000000000000000001110110001001",
			1873 => "00000000011011010001110110001001",
			1874 => "11111110010101100001110110001001",
			1875 => "0000001101000000000110111100001100",
			1876 => "0000000010000000000010110000000100",
			1877 => "00000001100101110001110110001001",
			1878 => "0000000111000000000101100100000100",
			1879 => "11111111110011000001110110001001",
			1880 => "00000000100001110001110110001001",
			1881 => "0000000111000000001011011100000100",
			1882 => "11111101101111010001110110001001",
			1883 => "0000000001000000001101011000001000",
			1884 => "0000000001000000001101011000000100",
			1885 => "00000000111000000001110110001001",
			1886 => "11111110011101000001110110001001",
			1887 => "0000001000000000000111000100000100",
			1888 => "00000001100010110001110110001001",
			1889 => "11111111001011000001110110001001",
			1890 => "0000000001000000001001011000000100",
			1891 => "11111110011011110001111000100101",
			1892 => "0000000001000000001101011001000100",
			1893 => "0000000011000000001110100100100100",
			1894 => "0000000001000000001100011000011100",
			1895 => "0000000100000000001001001100010000",
			1896 => "0000001100000000001000011000001000",
			1897 => "0000000111000000001011011100000100",
			1898 => "11111110100011100001111000100101",
			1899 => "00000000000000000001111000100101",
			1900 => "0000001010000000001001000100000100",
			1901 => "00000000011111000001111000100101",
			1902 => "11111111101111110001111000100101",
			1903 => "0000000110000000001001111100001000",
			1904 => "0000000011000000000010010100000100",
			1905 => "00000001001110010001111000100101",
			1906 => "00000000000000000001111000100101",
			1907 => "11111111011101010001111000100101",
			1908 => "0000000101000000000101110000000100",
			1909 => "00000000000000000001111000100101",
			1910 => "00000001011110100001111000100101",
			1911 => "0000000111000000000110110100001100",
			1912 => "0000000001000000001010011000000100",
			1913 => "00000000000000000001111000100101",
			1914 => "0000000001000000001101011000000100",
			1915 => "11111101111011110001111000100101",
			1916 => "00000000000000000001111000100101",
			1917 => "0000001010000000001001000100001000",
			1918 => "0000000001000000001101011000000100",
			1919 => "00000001000110110001111000100101",
			1920 => "11111111101101100001111000100101",
			1921 => "0000001011000000000010110100000100",
			1922 => "00000000000000000001111000100101",
			1923 => "0000001100000000000111010000000100",
			1924 => "00000000000000000001111000100101",
			1925 => "11111110110111100001111000100101",
			1926 => "0000001000000000000111000100000100",
			1927 => "00000001011100000001111000100101",
			1928 => "00000000000000000001111000100101",
			1929 => "0000000010000000001101101100001000",
			1930 => "0000001011000000001010010100000100",
			1931 => "11111110011010100001111011110011",
			1932 => "00000000000000000001111011110011",
			1933 => "0000000001000000001010011001001100",
			1934 => "0000001110000000000110111000101100",
			1935 => "0000000101000000000111111100011000",
			1936 => "0000000000000000001111000100001100",
			1937 => "0000001111000000001000110100001000",
			1938 => "0000001000000000000101000100000100",
			1939 => "00000000000000000001111011110011",
			1940 => "11111110011010000001111011110011",
			1941 => "00000000000000000001111011110011",
			1942 => "0000001100000000000100011000000100",
			1943 => "11111111010111100001111011110011",
			1944 => "0000001001000000001011001100000100",
			1945 => "00000000000000000001111011110011",
			1946 => "00000001001011110001111011110011",
			1947 => "0000001001000000001010100100010000",
			1948 => "0000001011000000000000110100001000",
			1949 => "0000001100000000001000011000000100",
			1950 => "00000000000000000001111011110011",
			1951 => "00000000101010100001111011110011",
			1952 => "0000000010000000000110111000000100",
			1953 => "00000000000000000001111011110011",
			1954 => "11111110111111000001111011110011",
			1955 => "00000001011010110001111011110011",
			1956 => "0000000111000000001011011100010100",
			1957 => "0000000100000000000100001100010000",
			1958 => "0000001011000000001110101100001000",
			1959 => "0000001111000000001000110100000100",
			1960 => "00000000000000000001111011110011",
			1961 => "11111101111100000001111011110011",
			1962 => "0000000000000000001000101100000100",
			1963 => "00000000001010100001111011110011",
			1964 => "00000000000000000001111011110011",
			1965 => "00000000000000000001111011110011",
			1966 => "0000001000000000001100000100000100",
			1967 => "00000001010100000001111011110011",
			1968 => "0000001011000000001110101100000100",
			1969 => "00000000000000000001111011110011",
			1970 => "11111110110000100001111011110011",
			1971 => "0000001110000000001000000100000100",
			1972 => "00000001100001100001111011110011",
			1973 => "0000000000000000000111000000000100",
			1974 => "11111110100011000001111011110011",
			1975 => "0000001000000000000111000100001000",
			1976 => "0000001100000000000001101000000100",
			1977 => "11111111110110100001111011110011",
			1978 => "00000001100100100001111011110011",
			1979 => "11111111001010010001111011110011",
			1980 => "00000000000000000001111011110101",
			1981 => "0000001011000000000010011100000100",
			1982 => "00000000000000000001111100000001",
			1983 => "11111100111110000001111100000001",
			1984 => "0000000101000000001111010100000100",
			1985 => "00000000000000000001111100001101",
			1986 => "11111110111000110001111100001101",
			1987 => "0000000100000000000101010100000100",
			1988 => "00000000000000000001111100100001",
			1989 => "0000000100000000000001100100000100",
			1990 => "00000000001010010001111100100001",
			1991 => "00000000000000000001111100100001",
			1992 => "0000001100000000000111010000001000",
			1993 => "0000001100000000001010111000000100",
			1994 => "00000000000000000001111100110101",
			1995 => "00000000001001110001111100110101",
			1996 => "11111111111110100001111100110101",
			1997 => "0000000101000000001111100100000100",
			1998 => "00000000000000000001111101001001",
			1999 => "0000001101000000001000101000000100",
			2000 => "11110010001011010001111101001001",
			2001 => "00000000000000000001111101001001",
			2002 => "0000000100000000000111011100001000",
			2003 => "0000001000000000000110001000000100",
			2004 => "00000000000000000001111101011101",
			2005 => "11111111011001110001111101011101",
			2006 => "00000000000000000001111101011101",
			2007 => "0000001101000000001100111000001100",
			2008 => "0000000100000000000000010100000100",
			2009 => "11111111111111000001111101111001",
			2010 => "0000000100000000000001100100000100",
			2011 => "00000000000110100001111101111001",
			2012 => "00000000000000000001111101111001",
			2013 => "11111111100011000001111101111001",
			2014 => "0000000100000000000101010100001000",
			2015 => "0000000100000000001110100100000100",
			2016 => "00000000000000000001111110011101",
			2017 => "11111111111101110001111110011101",
			2018 => "0000000100000000000001100100001000",
			2019 => "0000000100000000000011010100000100",
			2020 => "00000000000000000001111110011101",
			2021 => "00000000001011100001111110011101",
			2022 => "00000000000000000001111110011101",
			2023 => "0000001010000000000110011000001100",
			2024 => "0000001010000000001000010100000100",
			2025 => "00000000000000000001111111000001",
			2026 => "0000000110000000001111000000000100",
			2027 => "00000000000000000001111111000001",
			2028 => "00000000010010100001111111000001",
			2029 => "0000000110000000001000010000000100",
			2030 => "00000000000000000001111111000001",
			2031 => "11111111111001100001111111000001",
			2032 => "0000000001000000001100011000001100",
			2033 => "0000001010000000000110011100001000",
			2034 => "0000001010000000001000010100000100",
			2035 => "00000000000000000001111111100101",
			2036 => "11111111111000010001111111100101",
			2037 => "00000000000000000001111111100101",
			2038 => "0000001010000000001010110000000100",
			2039 => "00000000001011010001111111100101",
			2040 => "00000000000000000001111111100101",
			2041 => "0000001100000000001011011100001100",
			2042 => "0000000100000000000100001100000100",
			2043 => "00000000000000000010000000001001",
			2044 => "0000000100000000000001100100000100",
			2045 => "00000000000111000010000000001001",
			2046 => "00000000000000000010000000001001",
			2047 => "0000000111000000001011110100000100",
			2048 => "00000000000000000010000000001001",
			2049 => "11111111011010010010000000001001",
			2050 => "0000001010000000000110011000001100",
			2051 => "0000001010000000001000010100000100",
			2052 => "00000000000000000010000000110101",
			2053 => "0000000110000000001111000000000100",
			2054 => "00000000000000000010000000110101",
			2055 => "00000000010100110010000000110101",
			2056 => "0000000110000000001000010000000100",
			2057 => "00000000000000000010000000110101",
			2058 => "0000000000000000001000110000000100",
			2059 => "00000000000000000010000000110101",
			2060 => "11111111110111100010000000110101",
			2061 => "0000001000000000001011010100001100",
			2062 => "0000000000000000000111000000000100",
			2063 => "00000000000000000010000001100001",
			2064 => "0000000000000000000011111100000100",
			2065 => "00000000000010100010000001100001",
			2066 => "00000000000000000010000001100001",
			2067 => "0000000001000000001001100100001000",
			2068 => "0000000000000000001011000100000100",
			2069 => "11111111101001010010000001100001",
			2070 => "00000000000000000010000001100001",
			2071 => "00000000000000000010000001100001",
			2072 => "0000000100000000000111011100010000",
			2073 => "0000001000000000000110001000001100",
			2074 => "0000000100000000000101010100001000",
			2075 => "0000000100000000001110000000000100",
			2076 => "00000000000000000010000010000101",
			2077 => "11111111111111000010000010000101",
			2078 => "00000000000000000010000010000101",
			2079 => "11111111010110100010000010000101",
			2080 => "00000000000000000010000010000101",
			2081 => "0000000111000000000001001000010000",
			2082 => "0000000111000000000001011000000100",
			2083 => "00000000000000000010000010101001",
			2084 => "0000001011000000000000110100000100",
			2085 => "00000000000000000010000010101001",
			2086 => "0000001101000000001001100000000100",
			2087 => "00000000000000000010000010101001",
			2088 => "00000000001001110010000010101001",
			2089 => "11111111111111000010000010101001",
			2090 => "0000000010000000001000000100000100",
			2091 => "00000000000000000010000011001101",
			2092 => "0000000001000000001111000000001100",
			2093 => "0000000100000000001001000000001000",
			2094 => "0000001000000000001001101000000100",
			2095 => "00000000000000000010000011001101",
			2096 => "11111111100100010010000011001101",
			2097 => "00000000000000000010000011001101",
			2098 => "00000000000000000010000011001101",
			2099 => "0000001001000000001010100100010000",
			2100 => "0000000111000000001000011000001000",
			2101 => "0000001100000000001010111000000100",
			2102 => "00000000000000000010000100000001",
			2103 => "00000000000001010010000100000001",
			2104 => "0000000101000000000001000000000100",
			2105 => "00000000000000000010000100000001",
			2106 => "11111111101111110010000100000001",
			2107 => "0000001100000000000001101000000100",
			2108 => "00000000000000000010000100000001",
			2109 => "0000000111000000001011110100000100",
			2110 => "00000000011000000010000100000001",
			2111 => "00000000000000000010000100000001",
			2112 => "0000000100000000000100001100010000",
			2113 => "0000000100000000001100001100000100",
			2114 => "00000000000000000010000100110101",
			2115 => "0000000010000000001000110100001000",
			2116 => "0000001001000000000011101000000100",
			2117 => "11111111110100110010000100110101",
			2118 => "00000000000000000010000100110101",
			2119 => "00000000000000000010000100110101",
			2120 => "0000001001000000001001111100000100",
			2121 => "00000000000000000010000100110101",
			2122 => "0000000110000000000100101100000100",
			2123 => "00000000010100100010000100110101",
			2124 => "00000000000000000010000100110101",
			2125 => "0000001100000000001011011100010100",
			2126 => "0000000001000000001100011000001000",
			2127 => "0000001111000000001111101000000100",
			2128 => "00000000000000000010000101101001",
			2129 => "11111111111101110010000101101001",
			2130 => "0000000111000000001011011100000100",
			2131 => "00000000000000000010000101101001",
			2132 => "0000000001000000000100111100000100",
			2133 => "00000000001101010010000101101001",
			2134 => "00000000000000000010000101101001",
			2135 => "0000001011000000001111010000000100",
			2136 => "00000000000000000010000101101001",
			2137 => "11111101100111010010000101101001",
			2138 => "0000001100000000001011011100010100",
			2139 => "0000001001000000000010101100000100",
			2140 => "00000000000000000010000110011101",
			2141 => "0000000110000000001000010000000100",
			2142 => "00000000000000000010000110011101",
			2143 => "0000001001000000001001000100001000",
			2144 => "0000000101000000000101110000000100",
			2145 => "00000000000000000010000110011101",
			2146 => "00000000001111100010000110011101",
			2147 => "00000000000000000010000110011101",
			2148 => "0000001011000000001111010000000100",
			2149 => "00000000000000000010000110011101",
			2150 => "11111101111110110010000110011101",
			2151 => "0000001000000000001111001000010100",
			2152 => "0000001100000000001001110100000100",
			2153 => "00000000000000000010000111010001",
			2154 => "0000000000000000000010101000000100",
			2155 => "00000000000000000010000111010001",
			2156 => "0000001101000000000111111100000100",
			2157 => "00000000000000000010000111010001",
			2158 => "0000001100000000001011011100000100",
			2159 => "00000000000110110010000111010001",
			2160 => "00000000000000000010000111010001",
			2161 => "0000000000000000001011000100000100",
			2162 => "11111111101011000010000111010001",
			2163 => "00000000000000000010000111010001",
			2164 => "0000000101000000000000010000010100",
			2165 => "0000001011000000000000110100000100",
			2166 => "00000000000000000010000111111101",
			2167 => "0000000101000000001110010000000100",
			2168 => "00000000000000000010000111111101",
			2169 => "0000001100000000000001101000000100",
			2170 => "00000000000000000010000111111101",
			2171 => "0000001100000000001011011100000100",
			2172 => "00000000001011110010000111111101",
			2173 => "00000000000000000010000111111101",
			2174 => "11111111111110110010000111111101",
			2175 => "0000000111000000001011110100010100",
			2176 => "0000001001000000001001111100000100",
			2177 => "00000000000000000010001000111001",
			2178 => "0000000010000000000110111000000100",
			2179 => "00000000000000000010001000111001",
			2180 => "0000001000000000000111000100001000",
			2181 => "0000000111000000000001101000000100",
			2182 => "00000000000000000010001000111001",
			2183 => "00000000010011000010001000111001",
			2184 => "00000000000000000010001000111001",
			2185 => "0000000110000000001000010000000100",
			2186 => "00000000000000000010001000111001",
			2187 => "0000001011000000001101000100000100",
			2188 => "00000000000000000010001000111001",
			2189 => "11111111000111000010001000111001",
			2190 => "0000000100000000000000100000011000",
			2191 => "0000000001000000001101011000010000",
			2192 => "0000000000000000001010101100000100",
			2193 => "00000000000000000010001001111101",
			2194 => "0000000100000000001001000000001000",
			2195 => "0000001010000000001000010100000100",
			2196 => "00000000000000000010001001111101",
			2197 => "11111111101111000010001001111101",
			2198 => "00000000000000000010001001111101",
			2199 => "0000000110000000000100101100000100",
			2200 => "00000000010010000010001001111101",
			2201 => "00000000000000000010001001111101",
			2202 => "0000001010000000000101000100001000",
			2203 => "0000000001000000001001011000000100",
			2204 => "00000000000000000010001001111101",
			2205 => "00000001010111010010001001111101",
			2206 => "00000000000000000010001001111101",
			2207 => "0000000100000000000000010100010100",
			2208 => "0000000111000000001011011100010000",
			2209 => "0000001100000000001111011100001100",
			2210 => "0000000001000000001011001100001000",
			2211 => "0000001000000000000101000100000100",
			2212 => "00000000000000000010001011000001",
			2213 => "11111111101111110010001011000001",
			2214 => "00000000000000000010001011000001",
			2215 => "00000000000000000010001011000001",
			2216 => "00000000000000000010001011000001",
			2217 => "0000001000000000001111001000001100",
			2218 => "0000000001000000001011111100000100",
			2219 => "00000000000000000010001011000001",
			2220 => "0000000000000000000010011000000100",
			2221 => "00000000000000000010001011000001",
			2222 => "00000000101100000010001011000001",
			2223 => "00000000000000000010001011000001",
			2224 => "0000000100000000000000010100010100",
			2225 => "0000000000000000001010101100000100",
			2226 => "00000000000000000010001100000101",
			2227 => "0000001001000000001000100100001100",
			2228 => "0000000111000000000111110000001000",
			2229 => "0000001000000000000001010100000100",
			2230 => "00000000000000000010001100000101",
			2231 => "11111111101100100010001100000101",
			2232 => "00000000000000000010001100000101",
			2233 => "00000000000000000010001100000101",
			2234 => "0000001000000000000111000100001100",
			2235 => "0000000001000000001011111100000100",
			2236 => "00000000000000000010001100000101",
			2237 => "0000000000000000000010011000000100",
			2238 => "00000000000000000010001100000101",
			2239 => "00000000010001000010001100000101",
			2240 => "00000000000000000010001100000101",
			2241 => "0000000100000000000000100000011100",
			2242 => "0000000001000000001101011000010000",
			2243 => "0000001000000000000101000100000100",
			2244 => "00000000000000000010001101010001",
			2245 => "0000000100000000001001000000001000",
			2246 => "0000000000000000000001110100000100",
			2247 => "00000000000000000010001101010001",
			2248 => "11111111101101000010001101010001",
			2249 => "00000000000000000010001101010001",
			2250 => "0000001000000000001111001000001000",
			2251 => "0000001101000000001110110100000100",
			2252 => "00000000000000000010001101010001",
			2253 => "00000000011011010010001101010001",
			2254 => "00000000000000000010001101010001",
			2255 => "0000001010000000000101000100001000",
			2256 => "0000000001000000001001011000000100",
			2257 => "00000000000000000010001101010001",
			2258 => "00000001011011110010001101010001",
			2259 => "00000000000000000010001101010001",
			2260 => "0000000100000000000000010100011100",
			2261 => "0000001011000000000000110100010000",
			2262 => "0000000000000000000001110100000100",
			2263 => "00000000000000000010001110100101",
			2264 => "0000001001000000000011101000001000",
			2265 => "0000000111000000000110110100000100",
			2266 => "11111111101000100010001110100101",
			2267 => "00000000000000000010001110100101",
			2268 => "00000000000000000010001110100101",
			2269 => "0000001010000000000001010000001000",
			2270 => "0000000110000000001111000000000100",
			2271 => "00000000000000000010001110100101",
			2272 => "00000000000010100010001110100101",
			2273 => "00000000000000000010001110100101",
			2274 => "0000001010000000000101000100001100",
			2275 => "0000001001000000001011001100000100",
			2276 => "00000000000000000010001110100101",
			2277 => "0000000111000000001111011100000100",
			2278 => "00000000111000010010001110100101",
			2279 => "00000000000000000010001110100101",
			2280 => "00000000000000000010001110100101",
			2281 => "0000001100000000001011011100011000",
			2282 => "0000001010000000001000010100000100",
			2283 => "00000000000000000010001111100001",
			2284 => "0000001001000000001011001100000100",
			2285 => "00000000000000000010001111100001",
			2286 => "0000001010000000000101000100001100",
			2287 => "0000001001000000001000010100001000",
			2288 => "0000001100000000001010111000000100",
			2289 => "00000000000000000010001111100001",
			2290 => "00000000001110000010001111100001",
			2291 => "00000000000000000010001111100001",
			2292 => "00000000000000000010001111100001",
			2293 => "0000001000000000000110001000000100",
			2294 => "00000000000000000010001111100001",
			2295 => "11111110011101100010001111100001",
			2296 => "0000000100000000000011011000011100",
			2297 => "0000001001000000001010100100000100",
			2298 => "11111111101101100010010000101101",
			2299 => "0000000011000000001110100100001100",
			2300 => "0000001011000000001101000100001000",
			2301 => "0000001101000000001100010100000100",
			2302 => "00000000000000000010010000101101",
			2303 => "00000000011101110010010000101101",
			2304 => "00000000000000000010010000101101",
			2305 => "0000001001000000001000100100001000",
			2306 => "0000001000000000001001101000000100",
			2307 => "00000000000000000010010000101101",
			2308 => "11111111101101100010010000101101",
			2309 => "00000000000000000010010000101101",
			2310 => "0000001010000000000101000100001000",
			2311 => "0000000110000000001000010000000100",
			2312 => "00000000000000000010010000101101",
			2313 => "00000001100001000010010000101101",
			2314 => "00000000000000000010010000101101",
			2315 => "0000000111000000000001001000011000",
			2316 => "0000001100000000001000011000000100",
			2317 => "00000000000000000010010001100001",
			2318 => "0000000110000000000100101100010000",
			2319 => "0000001110000000000001011100000100",
			2320 => "00000000000000000010010001100001",
			2321 => "0000000010000000001000110100000100",
			2322 => "00000000000000000010010001100001",
			2323 => "0000001010000000000101000100000100",
			2324 => "00000000001111010010010001100001",
			2325 => "00000000000000000010010001100001",
			2326 => "00000000000000000010010001100001",
			2327 => "11111111101110110010010001100001",
			2328 => "0000001111000000001111101000010000",
			2329 => "0000000001000000001001011000000100",
			2330 => "00000000000000000010010010101101",
			2331 => "0000000010000000001100111000000100",
			2332 => "00000000000000000010010010101101",
			2333 => "0000000001000000001010011000000100",
			2334 => "00000000110100110010010010101101",
			2335 => "00000000000000000010010010101101",
			2336 => "0000001000000000000001010100000100",
			2337 => "00000000000000000010010010101101",
			2338 => "0000000011000000001011110000000100",
			2339 => "00000000000000000010010010101101",
			2340 => "0000000110000000000100111100000100",
			2341 => "00000000000000000010010010101101",
			2342 => "0000000100000000001110100100000100",
			2343 => "00000000000000000010010010101101",
			2344 => "0000001010000000001000010100000100",
			2345 => "00000000000000000010010010101101",
			2346 => "11111111101011000010010010101101",
			2347 => "0000001010000000000110011000011000",
			2348 => "0000001010000000001000010100000100",
			2349 => "00000000000000000010010100000001",
			2350 => "0000001100000000001001110100000100",
			2351 => "00000000000000000010010100000001",
			2352 => "0000000101000000001100010000001100",
			2353 => "0000000100000000001000011100000100",
			2354 => "00000000000000000010010100000001",
			2355 => "0000000001000000001110010100000100",
			2356 => "00000000000000000010010100000001",
			2357 => "00000001001011010010010100000001",
			2358 => "00000000000000000010010100000001",
			2359 => "0000000100000000001011001000001000",
			2360 => "0000001000000000000110001000000100",
			2361 => "00000000000000000010010100000001",
			2362 => "11111111101011100010010100000001",
			2363 => "0000001010000000000101000100001000",
			2364 => "0000001010000000001100011100000100",
			2365 => "00000000000000000010010100000001",
			2366 => "00000000001001100010010100000001",
			2367 => "00000000000000000010010100000001",
			2368 => "0000000100000000001001000000100000",
			2369 => "0000001000000000000001010100010000",
			2370 => "0000001011000000001011110100000100",
			2371 => "00000000000000000010010101011101",
			2372 => "0000000011000000001100001100001000",
			2373 => "0000000001000000000100110100000100",
			2374 => "00000000000000000010010101011101",
			2375 => "00000000100000100010010101011101",
			2376 => "00000000000000000010010101011101",
			2377 => "0000000001000000001101011000001100",
			2378 => "0000000100000000000011101100001000",
			2379 => "0000000000000000001010101100000100",
			2380 => "00000000000000000010010101011101",
			2381 => "11111111011001110010010101011101",
			2382 => "00000000000000000010010101011101",
			2383 => "00000000000000000010010101011101",
			2384 => "0000001000000000000001110100001100",
			2385 => "0000000000000000000011010000000100",
			2386 => "00000000000000000010010101011101",
			2387 => "0000000001000000000101011100000100",
			2388 => "00000000000000000010010101011101",
			2389 => "00000000111101110010010101011101",
			2390 => "11111111110101000010010101011101",
			2391 => "0000000100000000000000010100100000",
			2392 => "0000001011000000000000110100010100",
			2393 => "0000001000000000000101000100000100",
			2394 => "00000000000000000010010110111001",
			2395 => "0000000001000000001010011000001100",
			2396 => "0000000111000000000110110100001000",
			2397 => "0000001010000000001000100100000100",
			2398 => "00000000000000000010010110111001",
			2399 => "11111111101001110010010110111001",
			2400 => "00000000000000000010010110111001",
			2401 => "00000000000000000010010110111001",
			2402 => "0000001010000000000001010000001000",
			2403 => "0000000110000000001111000000000100",
			2404 => "00000000000000000010010110111001",
			2405 => "00000000000010010010010110111001",
			2406 => "00000000000000000010010110111001",
			2407 => "0000001000000000001111001000001100",
			2408 => "0000001100000000001000000000000100",
			2409 => "00000000000000000010010110111001",
			2410 => "0000000000000000000010011000000100",
			2411 => "00000000000000000010010110111001",
			2412 => "00000000110101110010010110111001",
			2413 => "00000000000000000010010110111001",
			2414 => "0000001011000000000101110100010100",
			2415 => "0000001100000000001010111000000100",
			2416 => "00000000000000000010011000010101",
			2417 => "0000000000000000000010011000000100",
			2418 => "00000000000000000010011000010101",
			2419 => "0000000110000000000101010000001000",
			2420 => "0000001001000000001011001100000100",
			2421 => "00000000000000000010011000010101",
			2422 => "00000000111100000010011000010101",
			2423 => "00000000000000000010011000010101",
			2424 => "0000000001000000001010011000010100",
			2425 => "0000001000000000000101000100000100",
			2426 => "00000000000000000010011000010101",
			2427 => "0000000011000000000101000000001100",
			2428 => "0000001001000000000011101000001000",
			2429 => "0000000101000000001001010000000100",
			2430 => "00000000000000000010011000010101",
			2431 => "11111111100100110010011000010101",
			2432 => "00000000000000000010011000010101",
			2433 => "00000000000000000010011000010101",
			2434 => "0000001000000000000111000100000100",
			2435 => "00000000001000110010011000010101",
			2436 => "00000000000000000010011000010101",
			2437 => "0000000110000000001001111100011100",
			2438 => "0000001001000000000100111100000100",
			2439 => "11111111110010010010011001100001",
			2440 => "0000001100000000001011011100010100",
			2441 => "0000000110000000001000010000000100",
			2442 => "00000000000000000010011001100001",
			2443 => "0000000010000000000011110000001100",
			2444 => "0000001101000000001010000100001000",
			2445 => "0000000110000000000101010000000100",
			2446 => "00000000110011100010011001100001",
			2447 => "00000000000000000010011001100001",
			2448 => "00000000000000000010011001100001",
			2449 => "00000000000000000010011001100001",
			2450 => "00000000000000000010011001100001",
			2451 => "0000001000000000000110001000000100",
			2452 => "00000000000000000010011001100001",
			2453 => "0000001111000000001000011100000100",
			2454 => "00000000000000000010011001100001",
			2455 => "11111111100100000010011001100001",
			2456 => "0000001000000000000110001000011100",
			2457 => "0000001101000000001010000100011000",
			2458 => "0000000010000000000010010100000100",
			2459 => "00000000000000000010011010101101",
			2460 => "0000001100000000000100000100010000",
			2461 => "0000001001000000001001111100000100",
			2462 => "00000000000000000010011010101101",
			2463 => "0000001110000000000010111000001000",
			2464 => "0000001100000000001001110100000100",
			2465 => "00000000000000000010011010101101",
			2466 => "00000000100001100010011010101101",
			2467 => "00000000000000000010011010101101",
			2468 => "00000000000000000010011010101101",
			2469 => "00000000000000000010011010101101",
			2470 => "0000000010000000000110111000000100",
			2471 => "00000000000000000010011010101101",
			2472 => "0000001110000000000011010100000100",
			2473 => "11111111110110110010011010101101",
			2474 => "00000000000000000010011010101101",
			2475 => "0000001000000000001100000100011100",
			2476 => "0000001011000000001110101100010000",
			2477 => "0000000001000000001010011000001100",
			2478 => "0000000000000000001010101100000100",
			2479 => "00000000000000000010011100100001",
			2480 => "0000000000000000001000110000000100",
			2481 => "11111111101001000010011100100001",
			2482 => "00000000000000000010011100100001",
			2483 => "00000000000000000010011100100001",
			2484 => "0000000001000000001101011000001000",
			2485 => "0000001001000000001010100100000100",
			2486 => "00000000000000000010011100100001",
			2487 => "00000000110101000010011100100001",
			2488 => "00000000000000000010011100100001",
			2489 => "0000000100000000000000010100001100",
			2490 => "0000001001000000001000100100001000",
			2491 => "0000001000000000001001101000000100",
			2492 => "00000000000000000010011100100001",
			2493 => "11111111011001000010011100100001",
			2494 => "00000000000000000010011100100001",
			2495 => "0000001000000000000001110100010000",
			2496 => "0000000110000000000100101100001100",
			2497 => "0000001011000000001111011100000100",
			2498 => "00000000000000000010011100100001",
			2499 => "0000000000000000000010011000000100",
			2500 => "00000000000000000010011100100001",
			2501 => "00000000010110000010011100100001",
			2502 => "00000000000000000010011100100001",
			2503 => "11111111111001110010011100100001",
			2504 => "0000001110000000000110111100001100",
			2505 => "0000000001000000001001011000000100",
			2506 => "00000000000000000010011101111101",
			2507 => "0000000100000000001111100000000100",
			2508 => "00000000000000000010011101111101",
			2509 => "00000010000000100010011101111101",
			2510 => "0000000110000000001000010000001100",
			2511 => "0000000111000000001111011100000100",
			2512 => "00000000000000000010011101111101",
			2513 => "0000001001000000001010100000000100",
			2514 => "00000000000000000010011101111101",
			2515 => "00000000000101000010011101111101",
			2516 => "0000001111000000001110000000000100",
			2517 => "00000000000000000010011101111101",
			2518 => "0000000001000000001101011000010000",
			2519 => "0000001110000000001000000100001100",
			2520 => "0000001011000000001011110100000100",
			2521 => "00000000000000000010011101111101",
			2522 => "0000001000000000000001010100000100",
			2523 => "00000000000000000010011101111101",
			2524 => "11111111011101110010011101111101",
			2525 => "00000000000000000010011101111101",
			2526 => "00000000000000000010011101111101",
			2527 => "0000001111000000001111101000010000",
			2528 => "0000001101000000001110101100000100",
			2529 => "00000000000000000010011111010001",
			2530 => "0000000010000000001101101100000100",
			2531 => "00000000000000000010011111010001",
			2532 => "0000000110000000001111000000000100",
			2533 => "00000000000000000010011111010001",
			2534 => "00000000000111110010011111010001",
			2535 => "0000001010000000001000010100000100",
			2536 => "00000000000000000010011111010001",
			2537 => "0000001110000000000011010100010100",
			2538 => "0000001011000000000101110100000100",
			2539 => "00000000000000000010011111010001",
			2540 => "0000000100000000001110100100000100",
			2541 => "00000000000000000010011111010001",
			2542 => "0000000000000000001010101100000100",
			2543 => "00000000000000000010011111010001",
			2544 => "0000000011000000000011101100000100",
			2545 => "11111111110001110010011111010001",
			2546 => "00000000000000000010011111010001",
			2547 => "00000000000000000010011111010001",
			2548 => "0000001110000000000110111100001100",
			2549 => "0000000001000000001001011000000100",
			2550 => "00000000000000000010100000110101",
			2551 => "0000000100000000001111100000000100",
			2552 => "00000000000000000010100000110101",
			2553 => "00000010010101010010100000110101",
			2554 => "0000001000000000000111000100100000",
			2555 => "0000000010000000001000110100010000",
			2556 => "0000000000000000001010101100000100",
			2557 => "00000000000000000010100000110101",
			2558 => "0000001111000000001000000100000100",
			2559 => "00000000000000000010100000110101",
			2560 => "0000000100000000001110100100000100",
			2561 => "00000000000000000010100000110101",
			2562 => "11111111101000000010100000110101",
			2563 => "0000001100000000001001110100000100",
			2564 => "00000000000000000010100000110101",
			2565 => "0000000100000000001100001100000100",
			2566 => "00000000000000000010100000110101",
			2567 => "0000001100000000001011011100000100",
			2568 => "00000000100001000010100000110101",
			2569 => "00000000000000000010100000110101",
			2570 => "0000001011000000000010001000000100",
			2571 => "00000000000000000010100000110101",
			2572 => "11111111100100110010100000110101",
			2573 => "0000000001000000000100110100010100",
			2574 => "0000000100000000000111011100000100",
			2575 => "11111111000011000010100010101001",
			2576 => "0000001000000000000001110100001100",
			2577 => "0000000000000000000000111000000100",
			2578 => "00000000000000000010100010101001",
			2579 => "0000000001000000001001011000000100",
			2580 => "00000000000000000010100010101001",
			2581 => "00000000100010000010100010101001",
			2582 => "00000000000000000010100010101001",
			2583 => "0000000011000000000110001100001100",
			2584 => "0000001100000000000100000100001000",
			2585 => "0000000111000000000111010000000100",
			2586 => "00000000000000000010100010101001",
			2587 => "00000000111001110010100010101001",
			2588 => "00000000000000000010100010101001",
			2589 => "0000001100000000000111010000010000",
			2590 => "0000001111000000000110001100000100",
			2591 => "00000000000000000010100010101001",
			2592 => "0000001010000000001001000100000100",
			2593 => "00000000000000000010100010101001",
			2594 => "0000000001000000001011001100000100",
			2595 => "11111111011000010010100010101001",
			2596 => "00000000000000000010100010101001",
			2597 => "0000000001000000000100111100001000",
			2598 => "0000001001000000000010101100000100",
			2599 => "00000000000000000010100010101001",
			2600 => "00000000010110110010100010101001",
			2601 => "00000000000000000010100010101001",
			2602 => "0000000100000000000011011000101000",
			2603 => "0000000001000000001010011000011000",
			2604 => "0000000111000000001011011100010100",
			2605 => "0000000100000000000000010100010000",
			2606 => "0000001000000000000101000100000100",
			2607 => "00000000000000000010100100001101",
			2608 => "0000001011000000001110101100001000",
			2609 => "0000001010000000001000100100000100",
			2610 => "00000000000000000010100100001101",
			2611 => "11111111010010100010100100001101",
			2612 => "00000000000000000010100100001101",
			2613 => "00000000000000000010100100001101",
			2614 => "00000000000000000010100100001101",
			2615 => "0000000111000000001011110100001100",
			2616 => "0000000111000000000111010000000100",
			2617 => "00000000000000000010100100001101",
			2618 => "0000001000000000000110001000000100",
			2619 => "00000000010001000010100100001101",
			2620 => "00000000000000000010100100001101",
			2621 => "00000000000000000010100100001101",
			2622 => "0000001010000000000101000100001000",
			2623 => "0000000110000000001000010000000100",
			2624 => "00000000000000000010100100001101",
			2625 => "00000001001111010010100100001101",
			2626 => "00000000000000000010100100001101",
			2627 => "0000001100000000001001110100001000",
			2628 => "0000001010000000000110011100000100",
			2629 => "11111111100010000010100101101001",
			2630 => "00000000000000000010100101101001",
			2631 => "0000001101000000000111011000010000",
			2632 => "0000000101000000000101110000000100",
			2633 => "00000000000000000010100101101001",
			2634 => "0000001100000000000001011000001000",
			2635 => "0000000001000000000111101000000100",
			2636 => "00000000000000000010100101101001",
			2637 => "00000000011111100010100101101001",
			2638 => "00000000000000000010100101101001",
			2639 => "0000000111000000000100010000010100",
			2640 => "0000000001000000001010011000000100",
			2641 => "00000000000000000010100101101001",
			2642 => "0000001100000000000111010000001100",
			2643 => "0000000101000000000110010000000100",
			2644 => "00000000000000000010100101101001",
			2645 => "0000001101000000000110111100000100",
			2646 => "00000000000000000010100101101001",
			2647 => "11111111100000010010100101101001",
			2648 => "00000000000000000010100101101001",
			2649 => "00000000000000000010100101101001",
			2650 => "0000000101000000001110000100010000",
			2651 => "0000001100000000001010111000000100",
			2652 => "00000000000000000010100111010101",
			2653 => "0000000100000000001111100000000100",
			2654 => "00000000000000000010100111010101",
			2655 => "0000001000000000001101010000000100",
			2656 => "00000001110110010010100111010101",
			2657 => "00000000000000000010100111010101",
			2658 => "0000000001000000001010011000011000",
			2659 => "0000000110000000000100111100000100",
			2660 => "00000000000000000010100111010101",
			2661 => "0000000111000000001111011100000100",
			2662 => "00000000000000000010100111010101",
			2663 => "0000001001000000000011101000001100",
			2664 => "0000000101000000001110110100001000",
			2665 => "0000001000000000000101000100000100",
			2666 => "00000000000000000010100111010101",
			2667 => "11111111011101110010100111010101",
			2668 => "00000000000000000010100111010101",
			2669 => "00000000000000000010100111010101",
			2670 => "0000000110000000000100101100001100",
			2671 => "0000000111000000000111010000000100",
			2672 => "00000000000000000010100111010101",
			2673 => "0000001010000000001000010100000100",
			2674 => "00000000000000000010100111010101",
			2675 => "00000000010011010010100111010101",
			2676 => "00000000000000000010100111010101",
			2677 => "0000000001000000001100011000101100",
			2678 => "0000001001000000001010100100011100",
			2679 => "0000000001000000000101011100000100",
			2680 => "11111110010010000010101001010001",
			2681 => "0000000111000000001000011000001000",
			2682 => "0000001001000000001000010000000100",
			2683 => "11111111110110010010101001010001",
			2684 => "11111110010100010010101001010001",
			2685 => "0000001110000000001111101000001100",
			2686 => "0000000110000000001000010000000100",
			2687 => "11111110010101110010101001010001",
			2688 => "0000001100000000001000011000000100",
			2689 => "00000111001001010010101001010001",
			2690 => "00000000001101100010101001010001",
			2691 => "11111110010111010010101001010001",
			2692 => "0000000111000000000111010000001000",
			2693 => "0000001100000000001001110100000100",
			2694 => "11111110010001010010101001010001",
			2695 => "00000000000000000010101001010001",
			2696 => "0000000110000000000101010000000100",
			2697 => "00000101011000010010101001010001",
			2698 => "00000000010010110010101001010001",
			2699 => "0000001011000000001011110100000100",
			2700 => "11111110010011010010101001010001",
			2701 => "0000001000000000000111000100001100",
			2702 => "0000000111000000000111010000000100",
			2703 => "00000001001000000010101001010001",
			2704 => "0000001100000000001011011100000100",
			2705 => "00000011100000110010101001010001",
			2706 => "00000010001110110010101001010001",
			2707 => "11111110010111010010101001010001",
			2708 => "0000000011000000001111100100010000",
			2709 => "0000001001000000001011001100000100",
			2710 => "00000000000000000010101011000101",
			2711 => "0000000100000000001111100000000100",
			2712 => "00000000000000000010101011000101",
			2713 => "0000001100000000000001111100000100",
			2714 => "00000000000000000010101011000101",
			2715 => "00000010001010110010101011000101",
			2716 => "0000000110000000001000010000010100",
			2717 => "0000001100000000001001110100000100",
			2718 => "00000000000000000010101011000101",
			2719 => "0000001100000000000100000100001100",
			2720 => "0000001011000000001011110100000100",
			2721 => "00000000000000000010101011000101",
			2722 => "0000001001000000001010100100000100",
			2723 => "00000000000000000010101011000101",
			2724 => "00000000011011100010101011000101",
			2725 => "00000000000000000010101011000101",
			2726 => "0000001111000000001110000000000100",
			2727 => "00000000000000000010101011000101",
			2728 => "0000001001000000000111110100010000",
			2729 => "0000001011000000001011110100000100",
			2730 => "00000000000000000010101011000101",
			2731 => "0000001000000000000001010100000100",
			2732 => "00000000000000000010101011000101",
			2733 => "0000000100000000001110100100000100",
			2734 => "00000000000000000010101011000101",
			2735 => "11111111100100110010101011000101",
			2736 => "00000000000000000010101011000101",
			2737 => "0000001111000000001111101000011000",
			2738 => "0000000001000000001001011000000100",
			2739 => "00000000000000000010101100101001",
			2740 => "0000000010000000001101101100000100",
			2741 => "00000000000000000010101100101001",
			2742 => "0000000110000000000101010000001100",
			2743 => "0000000110000000001111000000000100",
			2744 => "00000000000000000010101100101001",
			2745 => "0000001001000000000010101100000100",
			2746 => "00000000001010000010101100101001",
			2747 => "00000000000000000010101100101001",
			2748 => "00000000000000000010101100101001",
			2749 => "0000001000000000000001010100000100",
			2750 => "00000000000000000010101100101001",
			2751 => "0000001110000000000011010100010100",
			2752 => "0000001011000000000101110100000100",
			2753 => "00000000000000000010101100101001",
			2754 => "0000001010000000001000010100000100",
			2755 => "00000000000000000010101100101001",
			2756 => "0000000100000000001000011100000100",
			2757 => "00000000000000000010101100101001",
			2758 => "0000000000000000001010101100000100",
			2759 => "00000000000000000010101100101001",
			2760 => "11111111101101100010101100101001",
			2761 => "00000000000000000010101100101001",
			2762 => "0000001110000000001101101100011000",
			2763 => "0000001100000000001010111000000100",
			2764 => "00000000000000000010101110100101",
			2765 => "0000000110000000001001111100010000",
			2766 => "0000000010000000001101101100000100",
			2767 => "00000000000000000010101110100101",
			2768 => "0000000110000000001001100100000100",
			2769 => "00000000000000000010101110100101",
			2770 => "0000001100000000001000011000000100",
			2771 => "00000001000001010010101110100101",
			2772 => "00000000000000000010101110100101",
			2773 => "00000000000000000010101110100101",
			2774 => "0000000001000000001010011000011000",
			2775 => "0000000011000000000101000000010100",
			2776 => "0000001010000000001000100100000100",
			2777 => "00000000000000000010101110100101",
			2778 => "0000001001000000000011101000001100",
			2779 => "0000001000000000000101000100000100",
			2780 => "00000000000000000010101110100101",
			2781 => "0000000110000000000100111100000100",
			2782 => "00000000000000000010101110100101",
			2783 => "11111111100000100010101110100101",
			2784 => "00000000000000000010101110100101",
			2785 => "00000000000000000010101110100101",
			2786 => "0000001000000000000111000100001100",
			2787 => "0000000000000000001010101100000100",
			2788 => "00000000000000000010101110100101",
			2789 => "0000001011000000001010010100000100",
			2790 => "00000000000000000010101110100101",
			2791 => "00000000010000000010101110100101",
			2792 => "00000000000000000010101110100101",
			2793 => "0000000001000000001100011000110100",
			2794 => "0000001001000000001010100100100100",
			2795 => "0000000001000000000101011100000100",
			2796 => "11111110010011010010110000110001",
			2797 => "0000001100000000001001110100010000",
			2798 => "0000001001000000001000010000000100",
			2799 => "11111111110110000010110000110001",
			2800 => "0000001100000000001000000000000100",
			2801 => "11111110010100010010110000110001",
			2802 => "0000001100000000001000000000000100",
			2803 => "11111111100000010010110000110001",
			2804 => "11111110011110010010110000110001",
			2805 => "0000001110000000001111101000001100",
			2806 => "0000001001000000000100101100000100",
			2807 => "11111110010101000010110000110001",
			2808 => "0000000010000000001000000100000100",
			2809 => "11111110100101100010110000110001",
			2810 => "00000100100011110010110000110001",
			2811 => "11111110011000000010110000110001",
			2812 => "0000001011000000001011110100001000",
			2813 => "0000001100000000001001110100000100",
			2814 => "11111110010010100010110000110001",
			2815 => "00000000010011110010110000110001",
			2816 => "0000000110000000000101010000000100",
			2817 => "00000011111100100010110000110001",
			2818 => "00000000010011100010110000110001",
			2819 => "0000001011000000001011110100000100",
			2820 => "11111110010100100010110000110001",
			2821 => "0000001000000000000111000100001100",
			2822 => "0000001100000000001001110100000100",
			2823 => "00000001000000010010110000110001",
			2824 => "0000001100000000001011011100000100",
			2825 => "00000010111110100010110000110001",
			2826 => "00000001110010100010110000110001",
			2827 => "11111110011001110010110000110001",
			2828 => "0000001001000000001010100000010000",
			2829 => "0000000010000000000110111000000100",
			2830 => "11111110011011110010110011001101",
			2831 => "0000000010000000001110100100001000",
			2832 => "0000000100000000000100001100000100",
			2833 => "11111111110000010010110011001101",
			2834 => "00000000110101100010110011001101",
			2835 => "11111110110010000010110011001101",
			2836 => "0000000100000000000011110000101000",
			2837 => "0000001011000000000000110100010000",
			2838 => "0000001010000000001000100100000100",
			2839 => "00000000000000000010110011001101",
			2840 => "0000000001000000001010011000001000",
			2841 => "0000000001000000000100110100000100",
			2842 => "00000000000000000010110011001101",
			2843 => "11111110010001110010110011001101",
			2844 => "00000000000000000010110011001101",
			2845 => "0000000011000000001110100100000100",
			2846 => "00000001011100110010110011001101",
			2847 => "0000001110000000001110000000001000",
			2848 => "0000001110000000001110000000000100",
			2849 => "00000000000000000010110011001101",
			2850 => "11111101101111110010110011001101",
			2851 => "0000000111000000001011011100000100",
			2852 => "11111111001110100010110011001101",
			2853 => "0000000100000000001100001100000100",
			2854 => "11111111110011100010110011001101",
			2855 => "00000001000110100010110011001101",
			2856 => "0000001010000000001010110000001100",
			2857 => "0000001011000000000100010000000100",
			2858 => "00000000000000000010110011001101",
			2859 => "0000001011000000001100100100000100",
			2860 => "00000001011100110010110011001101",
			2861 => "00000000000000000010110011001101",
			2862 => "0000000100000000000011010100000100",
			2863 => "11111110110111100010110011001101",
			2864 => "0000001000000000000111000100000100",
			2865 => "00000001010010000010110011001101",
			2866 => "11111111010000000010110011001101",
			2867 => "0000001001000000000100111100000100",
			2868 => "11111111011010000010110101001001",
			2869 => "0000001111000000001100001100100000",
			2870 => "0000001011000000000110100000010100",
			2871 => "0000000110000000001001111100010000",
			2872 => "0000001000000000000001010100000100",
			2873 => "00000000000000000010110101001001",
			2874 => "0000000010000000000010010100000100",
			2875 => "00000000000000000010110101001001",
			2876 => "0000001100000000001010111000000100",
			2877 => "00000000000000000010110101001001",
			2878 => "00000000110001000010110101001001",
			2879 => "00000000000000000010110101001001",
			2880 => "0000000110000000001000010000000100",
			2881 => "00000000000000000010110101001001",
			2882 => "0000001000000000000001010100000100",
			2883 => "11111111110110100010110101001001",
			2884 => "00000000000000000010110101001001",
			2885 => "0000001001000000001000100100010000",
			2886 => "0000000111000000000111110000001100",
			2887 => "0000001110000000001000011100000100",
			2888 => "00000000000000000010110101001001",
			2889 => "0000000110000000000100111100000100",
			2890 => "00000000000000000010110101001001",
			2891 => "11111111010000000010110101001001",
			2892 => "00000000000000000010110101001001",
			2893 => "0000000110000000000100101100001000",
			2894 => "0000001100000000001010011100000100",
			2895 => "00000000000000000010110101001001",
			2896 => "00000000100010010010110101001001",
			2897 => "00000000000000000010110101001001",
			2898 => "0000001001000000001010100100100000",
			2899 => "0000000110000000000100111100001000",
			2900 => "0000001001000000001010100100000100",
			2901 => "11111110011001000010111000000101",
			2902 => "00000000000000000010111000000101",
			2903 => "0000001110000000001111101000010100",
			2904 => "0000000100000000001110111000000100",
			2905 => "11111110100100000010111000000101",
			2906 => "0000000110000000001000010000001000",
			2907 => "0000001100000000000100011000000100",
			2908 => "11111111001010010010111000000101",
			2909 => "00000010011100110010111000000101",
			2910 => "0000001001000000000111101100000100",
			2911 => "11111110100010010010111000000101",
			2912 => "00000000100111110010111000000101",
			2913 => "11111110011011010010111000000101",
			2914 => "0000001011000000000001001000011100",
			2915 => "0000000100000000000011110000010000",
			2916 => "0000000110000000000100111100001000",
			2917 => "0000000101000000000101110000000100",
			2918 => "11111110110110110010111000000101",
			2919 => "00000001011011000010111000000101",
			2920 => "0000000001000000001010011000000100",
			2921 => "11111110000100010010111000000101",
			2922 => "11111111100000000010111000000101",
			2923 => "0000001110000000000110111000000100",
			2924 => "00000010101000010010111000000101",
			2925 => "0000001001000000000011101000000100",
			2926 => "11111110110000110010111000000101",
			2927 => "00000000000010100010111000000101",
			2928 => "0000001011000000000110100000010000",
			2929 => "0000000110000000001001111100001100",
			2930 => "0000001100000000000100000100000100",
			2931 => "00000001101001010010111000000101",
			2932 => "0000001100000000000100000100000100",
			2933 => "00000000000000000010111000000101",
			2934 => "00000001011101100010111000000101",
			2935 => "11111111101011100010111000000101",
			2936 => "0000000000000000001010101100001000",
			2937 => "0000001111000000001000011100000100",
			2938 => "00000001010101010010111000000101",
			2939 => "11111110000000100010111000000101",
			2940 => "0000001110000000001011110000000100",
			2941 => "11111110111001010010111000000101",
			2942 => "0000000110000000000100101100000100",
			2943 => "00000001100111110010111000000101",
			2944 => "11111110110000010010111000000101",
			2945 => "0000001001000000000100101100000100",
			2946 => "11111111000001000010111010001001",
			2947 => "0000001111000000001110100100100000",
			2948 => "0000000010000000001011110000010000",
			2949 => "0000000111000000000001011000001100",
			2950 => "0000001000000000000101000100000100",
			2951 => "00000000000000000010111010001001",
			2952 => "0000000000000000001111000100000100",
			2953 => "11111111100001100010111010001001",
			2954 => "00000000000000000010111010001001",
			2955 => "00000000000000000010111010001001",
			2956 => "0000000111000000001011011100001100",
			2957 => "0000000110000000001001111100001000",
			2958 => "0000001101000000001010001000000100",
			2959 => "00000000000000000010111010001001",
			2960 => "00000000110101010010111010001001",
			2961 => "00000000000000000010111010001001",
			2962 => "00000000000000000010111010001001",
			2963 => "0000000111000000001011011100010000",
			2964 => "0000001001000000000111110100001100",
			2965 => "0000000100000000000100001100001000",
			2966 => "0000000001000000001011001100000100",
			2967 => "11111111000111100010111010001001",
			2968 => "00000000000000000010111010001001",
			2969 => "00000000000000000010111010001001",
			2970 => "00000000000000000010111010001001",
			2971 => "0000001000000000000111000100001100",
			2972 => "0000000100000000001100001100000100",
			2973 => "00000000000000000010111010001001",
			2974 => "0000000001000000000100110100000100",
			2975 => "00000000000000000010111010001001",
			2976 => "00000000110001000010111010001001",
			2977 => "00000000000000000010111010001001",
			2978 => "0000001001000000001010100000010100",
			2979 => "0000000110000000000100111100000100",
			2980 => "11111110011100000010111100110101",
			2981 => "0000001111000000000110111000001100",
			2982 => "0000001100000000001010111000000100",
			2983 => "00000000000000000010111100110101",
			2984 => "0000000100000000001001001100000100",
			2985 => "00000000000000000010111100110101",
			2986 => "00000000101110100010111100110101",
			2987 => "11111110110011010010111100110101",
			2988 => "0000000100000000000011110000101000",
			2989 => "0000001011000000000000110100010000",
			2990 => "0000000110000000000100111100001000",
			2991 => "0000000101000000000101110000000100",
			2992 => "00000000000000000010111100110101",
			2993 => "00000000100100010010111100110101",
			2994 => "0000000001000000001010011000000100",
			2995 => "11111110010011010010111100110101",
			2996 => "00000000000000000010111100110101",
			2997 => "0000001111000000001000011100000100",
			2998 => "00000001011011100010111100110101",
			2999 => "0000001001000000000011101000001000",
			3000 => "0000001100000000000100000100000100",
			3001 => "00000000111110010010111100110101",
			3002 => "11111111111100000010111100110101",
			3003 => "0000001000000000000001010100001000",
			3004 => "0000001101000000000110111100000100",
			3005 => "00000000000000000010111100110101",
			3006 => "11111101111110010010111100110101",
			3007 => "00000000010101100010111100110101",
			3008 => "0000000110000000001001111100001100",
			3009 => "0000001011000000000100010000000100",
			3010 => "00000000000000000010111100110101",
			3011 => "0000001111000000001010110100000100",
			3012 => "00000001011010100010111100110101",
			3013 => "00000000000000000010111100110101",
			3014 => "0000001001000000000011101000000100",
			3015 => "11111110111001000010111100110101",
			3016 => "0000000110000000000100101100001000",
			3017 => "0000001100000000001000011000000100",
			3018 => "00000000000000000010111100110101",
			3019 => "00000001011000000010111100110101",
			3020 => "11111111001011100010111100110101",
			3021 => "0000000000000000001011000101000000",
			3022 => "0000000100000000000111011100110000",
			3023 => "0000000111000000000001011000010000",
			3024 => "0000001000000000000101000100000100",
			3025 => "00000000000000000010111111001001",
			3026 => "0000001001000000000111110100001000",
			3027 => "0000001100000000001111011100000100",
			3028 => "11111111100000110010111111001001",
			3029 => "00000000000000000010111111001001",
			3030 => "00000000000000000010111111001001",
			3031 => "0000001100000000000111010000010000",
			3032 => "0000001001000000000000001000000100",
			3033 => "00000000000000000010111111001001",
			3034 => "0000000111000000000101110100001000",
			3035 => "0000000111000000000101100100000100",
			3036 => "00000000000000000010111111001001",
			3037 => "00000000011111000010111111001001",
			3038 => "00000000000000000010111111001001",
			3039 => "0000001010000000001001000100000100",
			3040 => "00000000000000000010111111001001",
			3041 => "0000000100000000000011110000000100",
			3042 => "00000000000000000010111111001001",
			3043 => "0000000010000000000101010100000100",
			3044 => "11111111110000110010111111001001",
			3045 => "00000000000000000010111111001001",
			3046 => "0000001000000000000001110100001100",
			3047 => "0000000000000000000011010000000100",
			3048 => "00000000000000000010111111001001",
			3049 => "0000001001000000000100111100000100",
			3050 => "00000000000000000010111111001001",
			3051 => "00000000101101010010111111001001",
			3052 => "00000000000000000010111111001001",
			3053 => "0000000000000000000000101000001000",
			3054 => "0000000100000000001001000000000100",
			3055 => "00000000000000000010111111001001",
			3056 => "00000011011000010010111111001001",
			3057 => "00000000000000000010111111001001",
			3058 => "0000000001000000001100011000110100",
			3059 => "0000001001000000001010100100101100",
			3060 => "0000001001000000001010100100100000",
			3061 => "0000000001000000000101011100000100",
			3062 => "11111110010000110011000001101101",
			3063 => "0000001100000000001001110100001100",
			3064 => "0000001001000000001000010000000100",
			3065 => "11111111101110100011000001101101",
			3066 => "0000001001000000001001111100000100",
			3067 => "11111110100101100011000001101101",
			3068 => "11111110010010000011000001101101",
			3069 => "0000001110000000001011101100001000",
			3070 => "0000001001000000000100101100000100",
			3071 => "11111110010101100011000001101101",
			3072 => "00000011101100010011000001101101",
			3073 => "0000001001000000001010100000000100",
			3074 => "11111110010110100011000001101101",
			3075 => "11111111011011010011000001101101",
			3076 => "0000001100000000000001101000001000",
			3077 => "0000000101000000001001010000000100",
			3078 => "11111110010010010011000001101101",
			3079 => "00000000011001100011000001101101",
			3080 => "00000011100000010011000001101101",
			3081 => "0000000110000000001000010000000100",
			3082 => "00000100011110010011000001101101",
			3083 => "11111110011011100011000001101101",
			3084 => "0000001101000000001100010100001000",
			3085 => "0000000100000000001101001000000100",
			3086 => "11111110010001110011000001101101",
			3087 => "00000000000000000011000001101101",
			3088 => "0000001010000000000110011100010000",
			3089 => "0000001100000000001001110100000100",
			3090 => "00000010000110100011000001101101",
			3091 => "0000000111000000000111010000000100",
			3092 => "00000010110111110011000001101101",
			3093 => "0000001100000000001011011100000100",
			3094 => "00000100011010100011000001101101",
			3095 => "00000011001000010011000001101101",
			3096 => "0000000111000000000101110100000100",
			3097 => "11111110011011000011000001101101",
			3098 => "00000000111010000011000001101101",
			3099 => "0000000001000000001100011000101100",
			3100 => "0000000001000000000101011100001100",
			3101 => "0000000001000000001001011000000100",
			3102 => "11111110011000000011000100110001",
			3103 => "0000000001000000001001011000000100",
			3104 => "00000000100000110011000100110001",
			3105 => "11111110011011110011000100110001",
			3106 => "0000000100000000000100001100010100",
			3107 => "0000000111000000000000011100001000",
			3108 => "0000000101000000001110010000000100",
			3109 => "11111110010111010011000100110001",
			3110 => "11111111111010110011000100110001",
			3111 => "0000000110000000001000010000001000",
			3112 => "0000000001000000001101111100000100",
			3113 => "11111110111010010011000100110001",
			3114 => "00000001110011000011000100110001",
			3115 => "11111110011101100011000100110001",
			3116 => "0000000010000000000110001100000100",
			3117 => "00000010111011000011000100110001",
			3118 => "0000000110000000000101010000000100",
			3119 => "00000001000100000011000100110001",
			3120 => "11111110011101010011000100110001",
			3121 => "0000001100000000001001110100001100",
			3122 => "0000000110000000000101010000001000",
			3123 => "0000001111000000001011110000000100",
			3124 => "11111110000010100011000100110001",
			3125 => "00000000111111100011000100110001",
			3126 => "11111110001110000011000100110001",
			3127 => "0000000110000000000100101100100100",
			3128 => "0000001011000000000001001000001100",
			3129 => "0000001100000000001000011000001000",
			3130 => "0000001000000000000001110000000100",
			3131 => "00000001100110110011000100110001",
			3132 => "11111110100010000011000100110001",
			3133 => "00000010000010010011000100110001",
			3134 => "0000000110000000001001111100010000",
			3135 => "0000001101000000001010000100001000",
			3136 => "0000001011000000000000110100000100",
			3137 => "00000001001110000011000100110001",
			3138 => "00000001101101100011000100110001",
			3139 => "0000001101000000001010000100000100",
			3140 => "00000000000000000011000100110001",
			3141 => "00000001101101010011000100110001",
			3142 => "0000000001000000001011001100000100",
			3143 => "11111111001111110011000100110001",
			3144 => "00000001110100000011000100110001",
			3145 => "0000000000000000000000110000000100",
			3146 => "11111110111101000011000100110001",
			3147 => "00000000010000110011000100110001",
			3148 => "0000000100000000001001000000111100",
			3149 => "0000001000000000000110001000110100",
			3150 => "0000000100000000000011110000100000",
			3151 => "0000001000000000000001010100010000",
			3152 => "0000000111000000000111010000000100",
			3153 => "00000000000000000011000111000101",
			3154 => "0000000011000000001100001100001000",
			3155 => "0000000001000000000100110100000100",
			3156 => "00000000000000000011000111000101",
			3157 => "00000000011110010011000111000101",
			3158 => "00000000000000000011000111000101",
			3159 => "0000001100000000000111010000001100",
			3160 => "0000000111000000000101110100001000",
			3161 => "0000001001000000000011101000000100",
			3162 => "11111111011001100011000111000101",
			3163 => "00000000000000000011000111000101",
			3164 => "00000000000000000011000111000101",
			3165 => "00000000000000000011000111000101",
			3166 => "0000001100000000001001110100000100",
			3167 => "00000000000000000011000111000101",
			3168 => "0000001100000000001011011100001100",
			3169 => "0000001110000000001101001000001000",
			3170 => "0000000001000000000111101000000100",
			3171 => "00000000000000000011000111000101",
			3172 => "00000000100101110011000111000101",
			3173 => "00000000000000000011000111000101",
			3174 => "00000000000000000011000111000101",
			3175 => "0000000010000000000101010100000100",
			3176 => "11111111001000010011000111000101",
			3177 => "00000000000000000011000111000101",
			3178 => "0000001000000000000001110100001100",
			3179 => "0000000000000000000011010000000100",
			3180 => "00000000000000000011000111000101",
			3181 => "0000000001000000000101011100000100",
			3182 => "00000000000000000011000111000101",
			3183 => "00000000111011100011000111000101",
			3184 => "11111111110110010011000111000101",
			3185 => "0000000010000000000010010100001100",
			3186 => "0000001000000000000101000100000100",
			3187 => "00000000000000000011001001111001",
			3188 => "0000000101000000000111111100000100",
			3189 => "11111110110101100011001001111001",
			3190 => "00000000000000000011001001111001",
			3191 => "0000001110000000000110111000100000",
			3192 => "0000000001000000000111101000010000",
			3193 => "0000000010000000001110000000001100",
			3194 => "0000000100000000000111011100000100",
			3195 => "00000000000000000011001001111001",
			3196 => "0000000110000000001111000000000100",
			3197 => "00000000000000000011001001111001",
			3198 => "00000000011010100011001001111001",
			3199 => "11111111011110000011001001111001",
			3200 => "0000001100000000000111010000001100",
			3201 => "0000001101000000001001011100000100",
			3202 => "00000000000000000011001001111001",
			3203 => "0000001100000000001001110100000100",
			3204 => "00000000000000000011001001111001",
			3205 => "00000000111000000011001001111001",
			3206 => "00000000000000000011001001111001",
			3207 => "0000000111000000000110110100010100",
			3208 => "0000000001000000001101011000001100",
			3209 => "0000001011000000001110101100001000",
			3210 => "0000000000000000001010101100000100",
			3211 => "00000000000000000011001001111001",
			3212 => "11111110110101100011001001111001",
			3213 => "00000000000000000011001001111001",
			3214 => "0000001000000000001011010100000100",
			3215 => "00000000000011000011001001111001",
			3216 => "00000000000000000011001001111001",
			3217 => "0000000011000000000011110000001100",
			3218 => "0000000100000000001110100100000100",
			3219 => "00000000000000000011001001111001",
			3220 => "0000000001000000000100110100000100",
			3221 => "00000000000000000011001001111001",
			3222 => "00000000101011000011001001111001",
			3223 => "0000000001000000001001100100001100",
			3224 => "0000001010000000001001000100000100",
			3225 => "00000000000000000011001001111001",
			3226 => "0000001100000000000111010000000100",
			3227 => "00000000000000000011001001111001",
			3228 => "11111111011111100011001001111001",
			3229 => "00000000000000000011001001111001",
			3230 => "0000000001000000001100011000101000",
			3231 => "0000000001000000000101011100000100",
			3232 => "11111110011000010011001100100101",
			3233 => "0000000100000000000100001100010100",
			3234 => "0000000111000000000000011100001000",
			3235 => "0000000101000000001110010000000100",
			3236 => "11111110010110110011001100100101",
			3237 => "11111111110111110011001100100101",
			3238 => "0000001001000000001010100000000100",
			3239 => "11111110100000100011001100100101",
			3240 => "0000000101000000000011001000000100",
			3241 => "00000001110111110011001100100101",
			3242 => "00000000000000000011001100100101",
			3243 => "0000000101000000001100010100001100",
			3244 => "0000001000000000000001110100001000",
			3245 => "0000001011000000000101110100000100",
			3246 => "00000011101001110011001100100101",
			3247 => "00000001111011110011001100100101",
			3248 => "00000000000000000011001100100101",
			3249 => "11111110011110110011001100100101",
			3250 => "0000001100000000001001110100001100",
			3251 => "0000001010000000001001000100001000",
			3252 => "0000000100000000001100001100000100",
			3253 => "11111110000001100011001100100101",
			3254 => "00000001000101010011001100100101",
			3255 => "11111110001011010011001100100101",
			3256 => "0000001000000000000001110100100000",
			3257 => "0000000001000000001100011000001100",
			3258 => "0000001010000000001000010100000100",
			3259 => "00000001110000100011001100100101",
			3260 => "0000001110000000000110111000000100",
			3261 => "00000001100001000011001100100101",
			3262 => "11111101101111010011001100100101",
			3263 => "0000001101000000000110111100000100",
			3264 => "00000001110001000011001100100101",
			3265 => "0000000000000000000111000000001000",
			3266 => "0000001111000000001000011100000100",
			3267 => "00000001100110110011001100100101",
			3268 => "11111110100100010011001100100101",
			3269 => "0000001010000000001010110000000100",
			3270 => "00000001110001100011001100100101",
			3271 => "00000000100011110011001100100101",
			3272 => "11111110101010010011001100100101",
			3273 => "0000000001000000000101011100000100",
			3274 => "11111110110000100011001110101001",
			3275 => "0000000010000000000011110000110100",
			3276 => "0000000101000000000110010000011100",
			3277 => "0000001001000000001010100100010100",
			3278 => "0000000100000000000100001100001100",
			3279 => "0000001000000000000001010100000100",
			3280 => "00000000000000000011001110101001",
			3281 => "0000000111000000001011011100000100",
			3282 => "11111111010001100011001110101001",
			3283 => "00000000000000000011001110101001",
			3284 => "0000000111000000000111010000000100",
			3285 => "00000000110110000011001110101001",
			3286 => "00000000000000000011001110101001",
			3287 => "0000001101000000001100010100000100",
			3288 => "00000000000000000011001110101001",
			3289 => "00000001001010000011001110101001",
			3290 => "0000001100000000001010001100010000",
			3291 => "0000001001000000000011101000000100",
			3292 => "00000000000000000011001110101001",
			3293 => "0000001010000000001000010100001000",
			3294 => "0000001101000000000110111100000100",
			3295 => "00000000000000000011001110101001",
			3296 => "11111110110101010011001110101001",
			3297 => "00000000000000000011001110101001",
			3298 => "0000000000000000001000110000000100",
			3299 => "00000000101010010011001110101001",
			3300 => "00000000000000000011001110101001",
			3301 => "0000001000000000001100000100000100",
			3302 => "00000000000000000011001110101001",
			3303 => "0000000001000000001011001100000100",
			3304 => "11111111010000110011001110101001",
			3305 => "00000000000000000011001110101001",
			3306 => "0000000010000000001100111000000100",
			3307 => "11111110100010010011010000100101",
			3308 => "0000000100000000001011001000110000",
			3309 => "0000001010000000001100011100100100",
			3310 => "0000000001000000001101011000011100",
			3311 => "0000000000000000001010101100001100",
			3312 => "0000000111000000000111010000000100",
			3313 => "00000000000000000011010000100101",
			3314 => "0000000001000000000100110100000100",
			3315 => "00000000000000000011010000100101",
			3316 => "00000001000011100011010000100101",
			3317 => "0000000100000000000011110000001000",
			3318 => "0000000111000000000110110100000100",
			3319 => "11111111000001110011010000100101",
			3320 => "00000000000000000011010000100101",
			3321 => "0000001010000000000110011000000100",
			3322 => "00000000101100010011010000100101",
			3323 => "00000000000000000011010000100101",
			3324 => "0000001101000000001001100000000100",
			3325 => "00000000000000000011010000100101",
			3326 => "00000001001011000011010000100101",
			3327 => "0000000010000000000010010100000100",
			3328 => "00000000000000000011010000100101",
			3329 => "0000001000000000000110001000000100",
			3330 => "00000000000000000011010000100101",
			3331 => "11111111000000010011010000100101",
			3332 => "0000001010000000000101000100001000",
			3333 => "0000000011000000001110010000000100",
			3334 => "00000000000000000011010000100101",
			3335 => "00000001101100100011010000100101",
			3336 => "11111111110011110011010000100101",
			3337 => "0000001001000000001010100100100100",
			3338 => "0000000110000000000100111100000100",
			3339 => "11111110011001000011010100000001",
			3340 => "0000000110000000001000010000001100",
			3341 => "0000000100000000001110111000000100",
			3342 => "11111110101101000011010100000001",
			3343 => "0000001100000000001010111000000100",
			3344 => "11111111010100000011010100000001",
			3345 => "00000010010011110011010100000001",
			3346 => "0000001001000000000100101100000100",
			3347 => "11111110011000000011010100000001",
			3348 => "0000000100000000000011101100001100",
			3349 => "0000001001000000000111101100001000",
			3350 => "0000001001000000000111101100000100",
			3351 => "11111111110011000011010100000001",
			3352 => "00000000000000000011010100000001",
			3353 => "11111110011101010011010100000001",
			3354 => "00000001001011000011010100000001",
			3355 => "0000001011000000000000110100100100",
			3356 => "0000001110000000000110111000010100",
			3357 => "0000000100000000001000001000010000",
			3358 => "0000000101000000000111111100001000",
			3359 => "0000000110000000000100111100000100",
			3360 => "00000000000111100011010100000001",
			3361 => "11111110010001100011010100000001",
			3362 => "0000001001000000001010100100000100",
			3363 => "00000000000000000011010100000001",
			3364 => "00000001011110010011010100000001",
			3365 => "00000010100101100011010100000001",
			3366 => "0000001110000000000110111000000100",
			3367 => "11110100010011010011010100000001",
			3368 => "0000001100000000001000011000001000",
			3369 => "0000001001000000000011101000000100",
			3370 => "11111110000001000011010100000001",
			3371 => "11111111011011110011010100000001",
			3372 => "00000001100110100011010100000001",
			3373 => "0000001101000000000110111100010000",
			3374 => "0000001100000000000001011000001000",
			3375 => "0000001110000000000011110000000100",
			3376 => "00000001101000010011010100000001",
			3377 => "00000000000000000011010100000001",
			3378 => "0000001011000000000110100000000100",
			3379 => "00000000111111010011010100000001",
			3380 => "11111111100100110011010100000001",
			3381 => "0000000111000000000110110100001000",
			3382 => "0000001010000000001000010100000100",
			3383 => "11111001001011100011010100000001",
			3384 => "00000000010111110011010100000001",
			3385 => "0000000110000000000100101100001100",
			3386 => "0000001110000000001000000100001000",
			3387 => "0000000111000000000101110100000100",
			3388 => "00000001100011000011010100000001",
			3389 => "11111110111000000011010100000001",
			3390 => "00000001101000110011010100000001",
			3391 => "11111110111011110011010100000001",
			3392 => "0000001100000000001000000000001100",
			3393 => "0000000010000000000110111000000100",
			3394 => "11111110011010010011010110111101",
			3395 => "0000000010000000000110111000000100",
			3396 => "00000000100101100011010110111101",
			3397 => "11111110101110000011010110111101",
			3398 => "0000000001000000001101011001000000",
			3399 => "0000000011000000001110100100100100",
			3400 => "0000001001000000001001111100001100",
			3401 => "0000001100000000001000000000001000",
			3402 => "0000000001000000000101011100000100",
			3403 => "00000000000000000011010110111101",
			3404 => "00000000010100000011010110111101",
			3405 => "11111110110000010011010110111101",
			3406 => "0000000110000000000100111100001000",
			3407 => "0000001111000000001000101000000100",
			3408 => "00000000000000000011010110111101",
			3409 => "00000001100101000011010110111101",
			3410 => "0000000100000000001010110100001000",
			3411 => "0000000001000000001100011000000100",
			3412 => "11111110101001110011010110111101",
			3413 => "00000000100011000011010110111101",
			3414 => "0000000110000000001001111100000100",
			3415 => "00000001011010010011010110111101",
			3416 => "00000000000000000011010110111101",
			3417 => "0000000111000000000110110100010000",
			3418 => "0000001001000000000010101100001000",
			3419 => "0000000110000000000101010000000100",
			3420 => "00000000001010100011010110111101",
			3421 => "00000000000000000011010110111101",
			3422 => "0000001001000000000011101000000100",
			3423 => "11111110100100010011010110111101",
			3424 => "11111100011111010011010110111101",
			3425 => "0000001010000000001010110000001000",
			3426 => "0000000001000000000100110100000100",
			3427 => "00000000000000000011010110111101",
			3428 => "00000001010111100011010110111101",
			3429 => "11111110101101010011010110111101",
			3430 => "0000001010000000001000010100001000",
			3431 => "0000001001000000000011101000000100",
			3432 => "00000001010000100011010110111101",
			3433 => "11111110101000000011010110111101",
			3434 => "0000000110000000000100101100001000",
			3435 => "0000001101000000001110110100000100",
			3436 => "00000000000000000011010110111101",
			3437 => "00000001100100100011010110111101",
			3438 => "00000000001010110011010110111101",
			3439 => "0000001001000000000100111100000100",
			3440 => "11111110011101010011011001011001",
			3441 => "0000000110000000000101010000110000",
			3442 => "0000000100000000000011110000100000",
			3443 => "0000000101000000000111111100000100",
			3444 => "11111110111001000011011001011001",
			3445 => "0000001111000000001000110100001100",
			3446 => "0000000001000000000100110100000100",
			3447 => "00000000000000000011011001011001",
			3448 => "0000001000000000000001110000000100",
			3449 => "00000001010110100011011001011001",
			3450 => "00000000000000000011011001011001",
			3451 => "0000001010000000001000010100001000",
			3452 => "0000000110000000001000010000000100",
			3453 => "00000000000000000011011001011001",
			3454 => "11111110101010010011011001011001",
			3455 => "0000000101000000000011001000000100",
			3456 => "00000000000000000011011001011001",
			3457 => "00000000101110000011011001011001",
			3458 => "0000000010000000000010110000001000",
			3459 => "0000000010000000000110111000000100",
			3460 => "00000000000000000011011001011001",
			3461 => "00000001010001100011011001011001",
			3462 => "0000000001000000001011001100000100",
			3463 => "11111111101110110011011001011001",
			3464 => "00000000000000000011011001011001",
			3465 => "0000000100000000000100001100001100",
			3466 => "0000001001000000001000100100001000",
			3467 => "0000001010000000000110011000000100",
			3468 => "00000000000000000011011001011001",
			3469 => "11111110101001000011011001011001",
			3470 => "00000000000000000011011001011001",
			3471 => "0000001000000000000111000100001000",
			3472 => "0000000001000000000100110100000100",
			3473 => "00000000000000000011011001011001",
			3474 => "00000000111111010011011001011001",
			3475 => "0000000110000000001001111100000100",
			3476 => "00000000001011100011011001011001",
			3477 => "11111110111000100011011001011001",
			3478 => "0000001100000000001010111000000100",
			3479 => "11111111000110110011011011100101",
			3480 => "0000000100000000000011010100110000",
			3481 => "0000000110000000000100111100001100",
			3482 => "0000000001000000000100110100000100",
			3483 => "00000000000000000011011011100101",
			3484 => "0000001011000000000100010000000100",
			3485 => "00000000000000000011011011100101",
			3486 => "00000000100010010011011011100101",
			3487 => "0000000001000000001100011000001000",
			3488 => "0000001111000000000010010100000100",
			3489 => "00000000000000000011011011100101",
			3490 => "11111111001110110011011011100101",
			3491 => "0000001000000000000001010100010000",
			3492 => "0000001011000000000110100000001000",
			3493 => "0000001000000000000101000100000100",
			3494 => "11111111110110010011011011100101",
			3495 => "00000000010010110011011011100101",
			3496 => "0000001000000000000001010100000100",
			3497 => "00000000000000000011011011100101",
			3498 => "11111111100110000011011011100101",
			3499 => "0000000010000000000010110000001000",
			3500 => "0000000101000000000111111100000100",
			3501 => "00000000000000000011011011100101",
			3502 => "00000000011111110011011011100101",
			3503 => "00000000000000000011011011100101",
			3504 => "0000001010000000000101000100010000",
			3505 => "0000000001000000000101011100000100",
			3506 => "00000000000000000011011011100101",
			3507 => "0000001101000000001001100000000100",
			3508 => "00000000110111110011011011100101",
			3509 => "0000001101000000001010000100000100",
			3510 => "00000000000000000011011011100101",
			3511 => "00000000010010010011011011100101",
			3512 => "00000000000000000011011011100101",
			3513 => "0000001001000000001010100100101000",
			3514 => "0000000010000000001101101100000100",
			3515 => "11111110011000010011011110100001",
			3516 => "0000000110000000000101010000100000",
			3517 => "0000000100000000001110111000001100",
			3518 => "0000001100000000001000011000000100",
			3519 => "11111110010111110011011110100001",
			3520 => "0000000111000000000001011000000100",
			3521 => "00000000101100110011011110100001",
			3522 => "11111110111101110011011110100001",
			3523 => "0000001001000000001011001100000100",
			3524 => "11111110100100110011011110100001",
			3525 => "0000000010000000000101000000001000",
			3526 => "0000000111000000001011000000000100",
			3527 => "11111111100100010011011110100001",
			3528 => "00000011011100000011011110100001",
			3529 => "0000000001000000000111101000000100",
			3530 => "11111110011011110011011110100001",
			3531 => "00000010000000010011011110100001",
			3532 => "11111110011000110011011110100001",
			3533 => "0000001100000000001001110100001000",
			3534 => "0000000101000000000111111100000100",
			3535 => "11111110010001000011011110100001",
			3536 => "00000000110000110011011110100001",
			3537 => "0000001000000000001001101000011100",
			3538 => "0000001101000000001010000100010100",
			3539 => "0000001011000000000001001000001000",
			3540 => "0000000001000000001100011000000100",
			3541 => "11111111010110100011011110100001",
			3542 => "00000001101101010011011110100001",
			3543 => "0000001101000000000110111100000100",
			3544 => "00000001101100000011011110100001",
			3545 => "0000001011000000001110101100000100",
			3546 => "11111111010000000011011110100001",
			3547 => "00000001011111010011011110100001",
			3548 => "0000000100000000000010110000000100",
			3549 => "11111110101011110011011110100001",
			3550 => "00000001100111100011011110100001",
			3551 => "0000000100000000000000010100001000",
			3552 => "0000000001000000001011001100000100",
			3553 => "11111101101110010011011110100001",
			3554 => "00000000110111000011011110100001",
			3555 => "0000001000000000000111000100001000",
			3556 => "0000001000000000001011010100000100",
			3557 => "00000000001101010011011110100001",
			3558 => "00000001111000010011011110100001",
			3559 => "11111110110001100011011110100001",
			3560 => "0000001001000000001010100100100100",
			3561 => "0000000010000000001101101100000100",
			3562 => "11111110011000010011100001010101",
			3563 => "0000000110000000000101010000011100",
			3564 => "0000000100000000001110111000001100",
			3565 => "0000001100000000001000011000000100",
			3566 => "11111110010111000011100001010101",
			3567 => "0000000111000000000001011000000100",
			3568 => "00000000110001100011100001010101",
			3569 => "11111110111011000011100001010101",
			3570 => "0000001001000000001011001100000100",
			3571 => "11111110100010110011100001010101",
			3572 => "0000000011000000001100010100000100",
			3573 => "00001010001001100011100001010101",
			3574 => "0000000010000000000011110000000100",
			3575 => "00000010101011010011100001010101",
			3576 => "00000000010111100011100001010101",
			3577 => "11111110011000100011100001010101",
			3578 => "0000000101000000000111111100001000",
			3579 => "0000001100000000001001110100000100",
			3580 => "11111110010000110011100001010101",
			3581 => "00000000111100010011100001010101",
			3582 => "0000000110000000001001111100100100",
			3583 => "0000001111000000000010111000011100",
			3584 => "0000001011000000000110100000001100",
			3585 => "0000000100000000001110111000001000",
			3586 => "0000001001000000001010100100000100",
			3587 => "00000000111010000011100001010101",
			3588 => "00000001101011100011100001010101",
			3589 => "00000010011110010011100001010101",
			3590 => "0000000000000000000111000000001000",
			3591 => "0000001001000000000011101000000100",
			3592 => "00000001101000010011100001010101",
			3593 => "11111110001111100011100001010101",
			3594 => "0000001101000000000111011000000100",
			3595 => "00000000000000000011100001010101",
			3596 => "00000001101100100011100001010101",
			3597 => "0000000101000000000110010000000100",
			3598 => "11111110011111010011100001010101",
			3599 => "00000001100110010011100001010101",
			3600 => "0000000001000000001001100100000100",
			3601 => "11111101011101110011100001010101",
			3602 => "0000000110000000000100101100000100",
			3603 => "00000001101111100011100001010101",
			3604 => "00000000000000000011100001010101",
			3605 => "0000001100000000001000000000001100",
			3606 => "0000000100000000001100111100000100",
			3607 => "11111110011101010011100100101001",
			3608 => "0000000100000000000000101100000100",
			3609 => "00000000000000000011100100101001",
			3610 => "11111111011101110011100100101001",
			3611 => "0000001011000000000110100000111100",
			3612 => "0000001100000000001000011000100100",
			3613 => "0000000111000000001111011100001100",
			3614 => "0000000100000000001000001000000100",
			3615 => "00000000000000000011100100101001",
			3616 => "0000001111000000001000011100000100",
			3617 => "00000001010101000011100100101001",
			3618 => "00000000000000000011100100101001",
			3619 => "0000000111000000000101100100001100",
			3620 => "0000001100000000001000000000000100",
			3621 => "00000000000000000011100100101001",
			3622 => "0000001000000000000101000100000100",
			3623 => "00000000000000000011100100101001",
			3624 => "11111110111001110011100100101001",
			3625 => "0000001011000000000001001000000100",
			3626 => "00000000000000000011100100101001",
			3627 => "0000000110000000000101010000000100",
			3628 => "00000000011111100011100100101001",
			3629 => "00000000000000000011100100101001",
			3630 => "0000001001000000001010100100001000",
			3631 => "0000001100000000001000011000000100",
			3632 => "00000000000000000011100100101001",
			3633 => "11111111100100100011100100101001",
			3634 => "0000001110000000001000011100000100",
			3635 => "00000001011010100011100100101001",
			3636 => "0000000011000000000110001100000100",
			3637 => "11111111100101010011100100101001",
			3638 => "0000001111000000001010110100000100",
			3639 => "00000000011110010011100100101001",
			3640 => "00000000000000000011100100101001",
			3641 => "0000001100000000000111010000010000",
			3642 => "0000000011000000001100001100000100",
			3643 => "00000000000000000011100100101001",
			3644 => "0000001011000000001101000100001000",
			3645 => "0000000010000000001100001100000100",
			3646 => "11111110001001000011100100101001",
			3647 => "00000000000000000011100100101001",
			3648 => "00000000000000000011100100101001",
			3649 => "0000001110000000001110000000001000",
			3650 => "0000000111000000000100010000000100",
			3651 => "00000000000000000011100100101001",
			3652 => "11111110111101010011100100101001",
			3653 => "0000000110000000000100101100001000",
			3654 => "0000001001000000000010101100000100",
			3655 => "00000000000000000011100100101001",
			3656 => "00000001010101100011100100101001",
			3657 => "11111111010100100011100100101001",
			3658 => "0000000001000000000100110100011100",
			3659 => "0000000110000000000100111100000100",
			3660 => "11111110011001010011100111010101",
			3661 => "0000000011000000000010010100010000",
			3662 => "0000000100000000000100001100000100",
			3663 => "11111110100100010011100111010101",
			3664 => "0000000111000000000111010000001000",
			3665 => "0000001100000000001010111000000100",
			3666 => "11111110111110000011100111010101",
			3667 => "00000010000101010011100111010101",
			3668 => "11111111100010000011100111010101",
			3669 => "0000000110000000001000010000000100",
			3670 => "11111111111111000011100111010101",
			3671 => "11111110011010110011100111010101",
			3672 => "0000001100000000001001110100000100",
			3673 => "11111110100101000011100111010101",
			3674 => "0000000110000000000100111100001000",
			3675 => "0000000000000000001000101100000100",
			3676 => "00000001100110100011100111010101",
			3677 => "00000100001011010011100111010101",
			3678 => "0000000001000000001010011000011000",
			3679 => "0000000111000000001011011100010000",
			3680 => "0000000100000000000011110000001000",
			3681 => "0000001011000000000000110100000100",
			3682 => "11111101010110010011100111010101",
			3683 => "00000000000000000011100111010101",
			3684 => "0000001110000000001000110100000100",
			3685 => "00000001011110100011100111010101",
			3686 => "11111110101011110011100111010101",
			3687 => "0000000110000000001000010000000100",
			3688 => "00000001100011000011100111010101",
			3689 => "11111110110110100011100111010101",
			3690 => "0000001011000000000110100000001100",
			3691 => "0000001110000000000010111000001000",
			3692 => "0000001101000000001001100000000100",
			3693 => "00000000010100010011100111010101",
			3694 => "00000001100111100011100111010101",
			3695 => "11111111011100000011100111010101",
			3696 => "0000001010000000001000010100000100",
			3697 => "11111101001100000011100111010101",
			3698 => "0000000110000000000100101100000100",
			3699 => "00000001010101010011100111010101",
			3700 => "11111111000001010011100111010101",
			3701 => "0000000010000000000011000000001000",
			3702 => "0000000101000000001110010000000100",
			3703 => "11111110100011100011101010100001",
			3704 => "00000000000000000011101010100001",
			3705 => "0000000011000000001100001100111000",
			3706 => "0000000001000000001100011000100100",
			3707 => "0000001111000000001011110000010100",
			3708 => "0000000111000000001111011100001100",
			3709 => "0000000100000000001000001000000100",
			3710 => "00000000000000000011101010100001",
			3711 => "0000000001000000000101011100000100",
			3712 => "00000000000000000011101010100001",
			3713 => "00000000111110000011101010100001",
			3714 => "0000000101000000000111111100000100",
			3715 => "11111111101011000011101010100001",
			3716 => "00000000000000000011101010100001",
			3717 => "0000000011000000001000000100001100",
			3718 => "0000000100000000001011100000001000",
			3719 => "0000000010000000000110111000000100",
			3720 => "00000000000000000011101010100001",
			3721 => "11111111000010010011101010100001",
			3722 => "00000000000000000011101010100001",
			3723 => "00000000000000000011101010100001",
			3724 => "0000000111000000000101110100001100",
			3725 => "0000001111000000000110001100001000",
			3726 => "0000001101000000001100010100000100",
			3727 => "00000000000000000011101010100001",
			3728 => "00000001010100010011101010100001",
			3729 => "00000000000000000011101010100001",
			3730 => "0000000101000000000010000000000100",
			3731 => "00000000000000000011101010100001",
			3732 => "11111111111101110011101010100001",
			3733 => "0000000000000000000111000000001100",
			3734 => "0000001001000000000010101100000100",
			3735 => "00000000000000000011101010100001",
			3736 => "0000001101000000000110111100000100",
			3737 => "00000000000000000011101010100001",
			3738 => "11111110101011100011101010100001",
			3739 => "0000000100000000001001001100001000",
			3740 => "0000000001000000001100011000000100",
			3741 => "00000000000000000011101010100001",
			3742 => "00000000111001000011101010100001",
			3743 => "0000001001000000001000100100001000",
			3744 => "0000001110000000001110100100000100",
			3745 => "00000000000000000011101010100001",
			3746 => "11111110111100010011101010100001",
			3747 => "0000001000000000000111000100001000",
			3748 => "0000001100000000001111011100000100",
			3749 => "00000000000000000011101010100001",
			3750 => "00000000111001010011101010100001",
			3751 => "11111111111011110011101010100001",
			3752 => "0000001100000000001000000000010000",
			3753 => "0000000100000000001100111100000100",
			3754 => "11111110011110010011101101110101",
			3755 => "0000000100000000000000101100001000",
			3756 => "0000000110000000001001100100000100",
			3757 => "00000000000000000011101101110101",
			3758 => "00000000001010100011101101110101",
			3759 => "11111111101000000011101101110101",
			3760 => "0000001011000000000110100001000000",
			3761 => "0000001100000000001000011000100100",
			3762 => "0000000010000000000010110000100000",
			3763 => "0000000100000000000011110000010000",
			3764 => "0000000101000000000111111100001000",
			3765 => "0000000110000000001111000000000100",
			3766 => "00000000000000000011101101110101",
			3767 => "11111110110010010011101101110101",
			3768 => "0000001010000000001001000100000100",
			3769 => "00000000010111100011101101110101",
			3770 => "11111111111011110011101101110101",
			3771 => "0000000110000000001000010000001000",
			3772 => "0000000010000000001100001100000100",
			3773 => "00000001001111010011101101110101",
			3774 => "00000000000000000011101101110101",
			3775 => "0000000001000000001101111100000100",
			3776 => "11111111101001100011101101110101",
			3777 => "00000000001011100011101101110101",
			3778 => "11111110110110100011101101110101",
			3779 => "0000000001000000001101111100001000",
			3780 => "0000001100000000001000011000000100",
			3781 => "00000000000000000011101101110101",
			3782 => "11111111101100010011101101110101",
			3783 => "0000001110000000001000011100001000",
			3784 => "0000001101000000001111010100000100",
			3785 => "00000001011000010011101101110101",
			3786 => "00000000000000000011101101110101",
			3787 => "0000000011000000000110001100000100",
			3788 => "11111111101001100011101101110101",
			3789 => "0000001111000000001010110100000100",
			3790 => "00000000011000010011101101110101",
			3791 => "00000000000000000011101101110101",
			3792 => "0000000001000000001101011000010000",
			3793 => "0000000110000000001000010000000100",
			3794 => "00000000000000000011101101110101",
			3795 => "0000001110000000001110100100001000",
			3796 => "0000000101000000000010000100000100",
			3797 => "11111110011100110011101101110101",
			3798 => "00000000000000000011101101110101",
			3799 => "00000000000000000011101101110101",
			3800 => "0000000110000000000100101100001000",
			3801 => "0000001100000000001010001100000100",
			3802 => "00000000000000000011101101110101",
			3803 => "00000001001101000011101101110101",
			3804 => "11111111010111110011101101110101",
			3805 => "0000001001000000001010100000101000",
			3806 => "0000000110000000000100111100000100",
			3807 => "11111110011001100011110001101001",
			3808 => "0000001111000000000110111000011000",
			3809 => "0000001100000000001010111000000100",
			3810 => "11111110111101010011110001101001",
			3811 => "0000001111000000001111101000001000",
			3812 => "0000001010000000000110011000000100",
			3813 => "00000000000000000011110001101001",
			3814 => "00000001101111110011110001101001",
			3815 => "0000001111000000000110111000001000",
			3816 => "0000000110000000001000010000000100",
			3817 => "00000000000000000011110001101001",
			3818 => "11111111010010010011110001101001",
			3819 => "00000000101100110011110001101001",
			3820 => "0000001101000000001100010100001000",
			3821 => "0000001101000000001010001000000100",
			3822 => "11111110111101100011110001101001",
			3823 => "00000000000000000011110001101001",
			3824 => "11111110011100010011110001101001",
			3825 => "0000000001000000001100011000101100",
			3826 => "0000001110000000000010010100011000",
			3827 => "0000000011000000000001011100001000",
			3828 => "0000001000000000001001101000000100",
			3829 => "11111110101101000011110001101001",
			3830 => "00000000000000000011110001101001",
			3831 => "0000000111000000000100010000001100",
			3832 => "0000000010000000001011110000001000",
			3833 => "0000000111000000000111010000000100",
			3834 => "11111110101010010011110001101001",
			3835 => "00000001011011000011110001101001",
			3836 => "00000001111101110011110001101001",
			3837 => "11111111011010100011110001101001",
			3838 => "0000001010000000001000010100000100",
			3839 => "00000001000111100011110001101001",
			3840 => "0000001001000000001010100100001100",
			3841 => "0000001001000000001010100100000100",
			3842 => "11111110110110100011110001101001",
			3843 => "0000000010000000000110001100000100",
			3844 => "00000000000000000011110001101001",
			3845 => "00000000000001000011110001101001",
			3846 => "11111101110000010011110001101001",
			3847 => "0000001000000000000110001000100000",
			3848 => "0000001101000000001010000100011000",
			3849 => "0000000111000000000111010000001100",
			3850 => "0000001110000000000110111000001000",
			3851 => "0000000010000000001011110000000100",
			3852 => "00000000000000000011110001101001",
			3853 => "00000001000011010011110001101001",
			3854 => "11111110111011000011110001101001",
			3855 => "0000000111000000000111110000001000",
			3856 => "0000001100000000000100000100000100",
			3857 => "00000001100110110011110001101001",
			3858 => "00000000110011110011110001101001",
			3859 => "00000000000000000011110001101001",
			3860 => "0000000010000000000101000000000100",
			3861 => "11111110101111000011110001101001",
			3862 => "00000001100000010011110001101001",
			3863 => "0000000111000000000010001000000100",
			3864 => "11111110101001110011110001101001",
			3865 => "00000000000000000011110001101001",
			3866 => "0000001100000000000100011000000100",
			3867 => "11111110011011000011110100001101",
			3868 => "0000000001000000001010011000111100",
			3869 => "0000000100000000000000010100101100",
			3870 => "0000001011000000000000110100011000",
			3871 => "0000001110000000000110111000010000",
			3872 => "0000001100000000000001101000001000",
			3873 => "0000000100000000000011001100000100",
			3874 => "11111110100010010011110100001101",
			3875 => "00000000000000000011110100001101",
			3876 => "0000001101000000001100010100000100",
			3877 => "00000000000000000011110100001101",
			3878 => "00000000111000010011110100001101",
			3879 => "0000001100000000001111011100000100",
			3880 => "11111110000100010011110100001101",
			3881 => "00000000000000000011110100001101",
			3882 => "0000001100000000000100000100001000",
			3883 => "0000001001000000001010100100000100",
			3884 => "00000000000000000011110100001101",
			3885 => "00000001011001100011110100001101",
			3886 => "0000001110000000001000110100001000",
			3887 => "0000000100000000000110001100000100",
			3888 => "00000000000000000011110100001101",
			3889 => "11111110101010110011110100001101",
			3890 => "00000000000000000011110100001101",
			3891 => "0000000110000000001001111100001100",
			3892 => "0000001101000000001100010000001000",
			3893 => "0000001001000000001011001100000100",
			3894 => "00000000000000000011110100001101",
			3895 => "00000001011010010011110100001101",
			3896 => "00000000000000000011110100001101",
			3897 => "11111110111101000011110100001101",
			3898 => "0000000011000000000101000000000100",
			3899 => "00000001100000000011110100001101",
			3900 => "0000000000000000000111000000000100",
			3901 => "11111110011101100011110100001101",
			3902 => "0000001000000000000111000100001000",
			3903 => "0000001100000000000001101000000100",
			3904 => "11111111110011100011110100001101",
			3905 => "00000001100001110011110100001101",
			3906 => "11111111001011010011110100001101",
			3907 => "0000001001000000000100111100000100",
			3908 => "11111110011100110011110111001001",
			3909 => "0000000011000000001110100100101100",
			3910 => "0000000010000000000011000000001000",
			3911 => "0000001011000000000001001000000100",
			3912 => "11111110111101010011110111001001",
			3913 => "00000000000000000011110111001001",
			3914 => "0000000001000000001100011000011100",
			3915 => "0000001110000000001000101000010000",
			3916 => "0000000001000000000111101000001000",
			3917 => "0000001111000000001111101000000100",
			3918 => "00000000101000010011110111001001",
			3919 => "11111111001110000011110111001001",
			3920 => "0000000111000000000110110100000100",
			3921 => "00000001010100010011110111001001",
			3922 => "00000000000000000011110111001001",
			3923 => "0000000100000000001110111000001000",
			3924 => "0000000110000000000100111100000100",
			3925 => "00000000000000000011110111001001",
			3926 => "11111110100100010011110111001001",
			3927 => "00000000001100010011110111001001",
			3928 => "0000001100000000001001110100000100",
			3929 => "00000000000000000011110111001001",
			3930 => "00000001011010110011110111001001",
			3931 => "0000000111000000000110110100010100",
			3932 => "0000000001000000001101011000001000",
			3933 => "0000001001000000000010101100000100",
			3934 => "00000000000000000011110111001001",
			3935 => "11111110011101100011110111001001",
			3936 => "0000001110000000000110001100000100",
			3937 => "00000000101011000011110111001001",
			3938 => "0000001000000000001001101000000100",
			3939 => "00000000000000000011110111001001",
			3940 => "11111111011110110011110111001001",
			3941 => "0000000111000000001011110100010100",
			3942 => "0000001001000000000010101100001100",
			3943 => "0000000110000000001001111100001000",
			3944 => "0000001001000000001010100100000100",
			3945 => "00000000000000000011110111001001",
			3946 => "00000000010010000011110111001001",
			3947 => "11111111010111110011110111001001",
			3948 => "0000000100000000001100001100000100",
			3949 => "00000000000000000011110111001001",
			3950 => "00000001001110000011110111001001",
			3951 => "0000001100000000000100000100000100",
			3952 => "00000000000000000011110111001001",
			3953 => "11111111001001110011110111001001",
			3954 => "0000001100000000001000000000000100",
			3955 => "11111110100011010011111010010101",
			3956 => "0000001011000000000110100001000100",
			3957 => "0000001100000000001000011000101000",
			3958 => "0000000111000000001111011100010000",
			3959 => "0000000111000000001000011000000100",
			3960 => "00000000000000000011111010010101",
			3961 => "0000000000000000001000110000000100",
			3962 => "00000000000000000011111010010101",
			3963 => "0000001111000000001000110100000100",
			3964 => "00000001001111110011111010010101",
			3965 => "00000000000000000011111010010101",
			3966 => "0000000110000000000101010000010000",
			3967 => "0000001011000000000001001000001000",
			3968 => "0000000010000000001000000100000100",
			3969 => "11111111001011010011111010010101",
			3970 => "00000000000000000011111010010101",
			3971 => "0000000001000000001101111100000100",
			3972 => "00000000000000000011111010010101",
			3973 => "00000000111001110011111010010101",
			3974 => "0000000010000000001110100100000100",
			3975 => "00000000000000000011111010010101",
			3976 => "11111110101110100011111010010101",
			3977 => "0000000001000000001101111100001000",
			3978 => "0000001100000000001000011000000100",
			3979 => "00000000000000000011111010010101",
			3980 => "11111111101010110011111010010101",
			3981 => "0000001110000000001000011100001000",
			3982 => "0000001111000000000011110000000100",
			3983 => "00000001011010000011111010010101",
			3984 => "00000000000000000011111010010101",
			3985 => "0000000011000000000110001100000100",
			3986 => "11111111100111100011111010010101",
			3987 => "0000001111000000001010110100000100",
			3988 => "00000000011010000011111010010101",
			3989 => "00000000000000000011111010010101",
			3990 => "0000000001000000001101011000010000",
			3991 => "0000000110000000001000010000000100",
			3992 => "00000000000000000011111010010101",
			3993 => "0000001110000000001110100100001000",
			3994 => "0000000101000000000010000100000100",
			3995 => "11111110010111100011111010010101",
			3996 => "00000000000000000011111010010101",
			3997 => "00000000000000000011111010010101",
			3998 => "0000000110000000000100101100001100",
			3999 => "0000000111000000000100010000001000",
			4000 => "0000001100000000001010001100000100",
			4001 => "11111111111100000011111010010101",
			4002 => "00000000000000000011111010010101",
			4003 => "00000001010001000011111010010101",
			4004 => "11111111010101110011111010010101",
			4005 => "0000001001000000000100111100000100",
			4006 => "11111110011100100011111101100011",
			4007 => "0000000110000000000101010001001100",
			4008 => "0000000000000000000111000000101000",
			4009 => "0000000110000000001000010000010100",
			4010 => "0000000111000000001011011100001100",
			4011 => "0000000001000000001010011000001000",
			4012 => "0000001011000000001110101100000100",
			4013 => "11111111000101110011111101100011",
			4014 => "00000000000000000011111101100011",
			4015 => "00000000100000110011111101100011",
			4016 => "0000000001000000000100110100000100",
			4017 => "00000000000000000011111101100011",
			4018 => "00000001010111100011111101100011",
			4019 => "0000001011000000000110100000001100",
			4020 => "0000000001000000001100011000000100",
			4021 => "11111110110011110011111101100011",
			4022 => "0000000011000000001110000000000100",
			4023 => "00000000000000000011111101100011",
			4024 => "00000000110010110011111101100011",
			4025 => "0000001111000000001000011100000100",
			4026 => "00000000000000000011111101100011",
			4027 => "11111110001111110011111101100011",
			4028 => "0000000010000000000010110000011100",
			4029 => "0000001100000000001011000000001100",
			4030 => "0000001110000000000010000000001000",
			4031 => "0000000011000000000110010000000100",
			4032 => "00000000000000000011111101100011",
			4033 => "00000000001011000011111101100011",
			4034 => "11111111011111000011111101100011",
			4035 => "0000000010000000001110000000001000",
			4036 => "0000000001000000001100011000000100",
			4037 => "11111111111011010011111101100011",
			4038 => "00000000000000000011111101100011",
			4039 => "0000000111000000000001101000000100",
			4040 => "00000000000000000011111101100011",
			4041 => "00000001011011100011111101100011",
			4042 => "0000000001000000001011001100000100",
			4043 => "11111111101001000011111101100011",
			4044 => "00000000000000000011111101100011",
			4045 => "0000000001000000001101011000001100",
			4046 => "0000000000000000000000110000001000",
			4047 => "0000000111000000000111110000000100",
			4048 => "11111110101101010011111101100011",
			4049 => "00000000000000000011111101100011",
			4050 => "00000000000000000011111101100011",
			4051 => "0000001000000000001111001000001000",
			4052 => "0000000010000000000101000000000100",
			4053 => "00000000000000000011111101100011",
			4054 => "00000000111111010011111101100011",
			4055 => "11111111011110110011111101100011",
			4056 => "00000000000000000011111101100101",
			4057 => "0000000101000000001111010100000100",
			4058 => "00000000000000000011111101110001",
			4059 => "11111110101111110011111101110001",
			4060 => "0000001100000000001011011100000100",
			4061 => "00000000000000000011111101111101",
			4062 => "11111111100110100011111101111101",
			4063 => "0000000100000000000011010100000100",
			4064 => "11111111111110100011111110010001",
			4065 => "0000000100000000000001100100000100",
			4066 => "00000000000011000011111110010001",
			4067 => "00000000000000000011111110010001",
			4068 => "0000001000000000000110001000001000",
			4069 => "0000001000000000000001010100000100",
			4070 => "00000000000000000011111110100101",
			4071 => "00000000000100110011111110100101",
			4072 => "00000000000000000011111110100101",
			4073 => "0000000101000000001111100100000100",
			4074 => "00000000000000000011111110111001",
			4075 => "0000001101000000001000101000000100",
			4076 => "11111011010001100011111110111001",
			4077 => "00000000000000000011111110111001",
			4078 => "0000000111000000000001001000001100",
			4079 => "0000000100000000000100001100000100",
			4080 => "00000000000000000011111111010101",
			4081 => "0000000100000000000001100100000100",
			4082 => "00000000001100110011111111010101",
			4083 => "00000000000000000011111111010101",
			4084 => "11111111011011000011111111010101",
			4085 => "0000000111000000000001001000001100",
			4086 => "0000000100000000000000010100000100",
			4087 => "00000000000000000011111111110001",
			4088 => "0000000100000000000001100100000100",
			4089 => "00000000000110100011111111110001",
			4090 => "00000000000000000011111111110001",
			4091 => "11111111100101010011111111110001",
			4092 => "0000000100000000000100001100001100",
			4093 => "0000000100000000001110100100000100",
			4094 => "00000000000000000100000000010101",
			4095 => "0000000100000000000000010100000100",
			4096 => "11111111111100010100000000010101",
			4097 => "00000000000000000100000000010101",
			4098 => "0000000100000000000001100100000100",
			4099 => "00000000000111010100000000010101",
			4100 => "00000000000000000100000000010101",
			4101 => "0000000001000000001100011000001100",
			4102 => "0000001010000000000110011100001000",
			4103 => "0000001010000000001000010100000100",
			4104 => "00000000000000000100000000111001",
			4105 => "11111111110110100100000000111001",
			4106 => "00000000000000000100000000111001",
			4107 => "0000001010000000001010110000000100",
			4108 => "00000000001111000100000000111001",
			4109 => "00000000000000000100000000111001",
			4110 => "0000001100000000000111010000001100",
			4111 => "0000001100000000001010111000000100",
			4112 => "00000000000000000100000001011101",
			4113 => "0000001011000000000110100000000100",
			4114 => "00000000010000010100000001011101",
			4115 => "00000000000000000100000001011101",
			4116 => "0000000111000000001011011100000100",
			4117 => "00000000000000000100000001011101",
			4118 => "11111111111101010100000001011101",
			4119 => "0000000100000000000100001100001100",
			4120 => "0000000100000000001100001100000100",
			4121 => "00000000000000000100000010001001",
			4122 => "0000001001000000001000100100000100",
			4123 => "11111111111011010100000010001001",
			4124 => "00000000000000000100000010001001",
			4125 => "0000001001000000001001111100000100",
			4126 => "00000000000000000100000010001001",
			4127 => "0000000110000000000100101100000100",
			4128 => "00000000010010110100000010001001",
			4129 => "00000000000000000100000010001001",
			4130 => "0000001001000000001010100100001100",
			4131 => "0000000111000000001000011000001000",
			4132 => "0000001100000000001010111000000100",
			4133 => "00000000000000000100000010110101",
			4134 => "00000000000001000100000010110101",
			4135 => "11111111110001110100000010110101",
			4136 => "0000001100000000000001101000000100",
			4137 => "00000000000000000100000010110101",
			4138 => "0000000111000000001011110100000100",
			4139 => "00000000010101110100000010110101",
			4140 => "00000000000000000100000010110101",
			4141 => "0000001100000000000111010000010000",
			4142 => "0000001100000000001010111000000100",
			4143 => "00000000000000000100000011011001",
			4144 => "0000001101000000001010000100001000",
			4145 => "0000001101000000001110101100000100",
			4146 => "00000000000000000100000011011001",
			4147 => "00000000001111010100000011011001",
			4148 => "00000000000000000100000011011001",
			4149 => "11111111111110010100000011011001",
			4150 => "0000001101000000001100111000010000",
			4151 => "0000001100000000000100011000000100",
			4152 => "00000000000000000100000011111101",
			4153 => "0000000110000000000100101100001000",
			4154 => "0000000110000000001001100100000100",
			4155 => "00000000000000000100000011111101",
			4156 => "00000000000101110100000011111101",
			4157 => "00000000000000000100000011111101",
			4158 => "11111111110100110100000011111101",
			4159 => "0000001111000000001110100100000100",
			4160 => "00000000000000000100000100100001",
			4161 => "0000000001000000001111000000001100",
			4162 => "0000001010000000001000010100000100",
			4163 => "00000000000000000100000100100001",
			4164 => "0000000011000000000011101100000100",
			4165 => "11111111100001010100000100100001",
			4166 => "00000000000000000100000100100001",
			4167 => "00000000000000000100000100100001",
			4168 => "0000001001000000001010100100001000",
			4169 => "0000001011000000000101110100000100",
			4170 => "00000000000000000100000101001101",
			4171 => "11111111101111010100000101001101",
			4172 => "0000001100000000000001101000000100",
			4173 => "00000000000000000100000101001101",
			4174 => "0000001000000000000111000100001000",
			4175 => "0000000000000000000111000000000100",
			4176 => "00000000000000000100000101001101",
			4177 => "00000000100011100100000101001101",
			4178 => "00000000000000000100000101001101",
			4179 => "0000000111000000000001001000010100",
			4180 => "0000000100000000000000010100001000",
			4181 => "0000000001000000001101011000000100",
			4182 => "11111111111110010100000101111001",
			4183 => "00000000000000000100000101111001",
			4184 => "0000001001000000001001111100000100",
			4185 => "00000000000000000100000101111001",
			4186 => "0000000110000000000100101100000100",
			4187 => "00000000010100010100000101111001",
			4188 => "00000000000000000100000101111001",
			4189 => "11111110111101000100000101111001",
			4190 => "0000000100000000000000010100001100",
			4191 => "0000000100000000001110100100000100",
			4192 => "00000000000000000100000110101101",
			4193 => "0000001111000000001010110100000100",
			4194 => "11111111111010000100000110101101",
			4195 => "00000000000000000100000110101101",
			4196 => "0000000100000000000001100100001100",
			4197 => "0000000010000000001101101100000100",
			4198 => "00000000000000000100000110101101",
			4199 => "0000000010000000001110100100000100",
			4200 => "00000000001110000100000110101101",
			4201 => "00000000000000000100000110101101",
			4202 => "00000000000000000100000110101101",
			4203 => "0000001000000000001111001000010000",
			4204 => "0000000100000000000000010100000100",
			4205 => "00000000000000000100000111100001",
			4206 => "0000000111000000000001101000000100",
			4207 => "00000000000000000100000111100001",
			4208 => "0000000000000000000010011000000100",
			4209 => "00000000000000000100000111100001",
			4210 => "00000000001011000100000111100001",
			4211 => "0000000100000000000000101100001000",
			4212 => "0000001010000000001100011100000100",
			4213 => "00000000000000000100000111100001",
			4214 => "11111111100011110100000111100001",
			4215 => "00000000000000000100000111100001",
			4216 => "0000001000000000000110001000010100",
			4217 => "0000000100000000001110100100000100",
			4218 => "00000000000000000100001000010101",
			4219 => "0000001100000000001001110100000100",
			4220 => "00000000000000000100001000010101",
			4221 => "0000000111000000001011110100001000",
			4222 => "0000000001000000001110010100000100",
			4223 => "00000000000000000100001000010101",
			4224 => "00000000010100000100001000010101",
			4225 => "00000000000000000100001000010101",
			4226 => "0000000100000000001001000000000100",
			4227 => "11111111010011100100001000010101",
			4228 => "00000000000000000100001000010101",
			4229 => "0000001011000000000110100000010100",
			4230 => "0000001011000000001010011100000100",
			4231 => "00000000000000000100001001000001",
			4232 => "0000000010000000000010110000001100",
			4233 => "0000000010000000001100111000000100",
			4234 => "00000000000000000100001001000001",
			4235 => "0000000011000000000101000000000100",
			4236 => "00000000010011110100001001000001",
			4237 => "00000000000000000100001001000001",
			4238 => "00000000000000000100001001000001",
			4239 => "00000000000000000100001001000001",
			4240 => "0000001011000000000101110100010000",
			4241 => "0000001100000000000100011000000100",
			4242 => "00000000000000000100001010000101",
			4243 => "0000000100000000000100001100000100",
			4244 => "00000000000000000100001010000101",
			4245 => "0000001000000000000111000000000100",
			4246 => "00000001001100100100001010000101",
			4247 => "00000000000000000100001010000101",
			4248 => "0000001000000000000110001000001100",
			4249 => "0000001100000000000001101000000100",
			4250 => "00000000000000000100001010000101",
			4251 => "0000001100000000000100000100000100",
			4252 => "00000000001000000100001010000101",
			4253 => "00000000000000000100001010000101",
			4254 => "0000001110000000000011010100000100",
			4255 => "11111111100001010100001010000101",
			4256 => "00000000000000000100001010000101",
			4257 => "0000000111000000001011110100010100",
			4258 => "0000001001000000001001111100000100",
			4259 => "00000000000000000100001011000001",
			4260 => "0000000010000000000110111000000100",
			4261 => "00000000000000000100001011000001",
			4262 => "0000001000000000000111000100001000",
			4263 => "0000001100000000001001110100000100",
			4264 => "00000000000000000100001011000001",
			4265 => "00000000010011110100001011000001",
			4266 => "00000000000000000100001011000001",
			4267 => "0000000110000000001000010000000100",
			4268 => "00000000000000000100001011000001",
			4269 => "0000001011000000001101000100000100",
			4270 => "00000000000000000100001011000001",
			4271 => "11111111001010000100001011000001",
			4272 => "0000000100000000000100001100010100",
			4273 => "0000000001000000001101011000010000",
			4274 => "0000001000000000000101000100000100",
			4275 => "00000000000000000100001100000101",
			4276 => "0000000101000000001110110100001000",
			4277 => "0000000110000000000100111100000100",
			4278 => "00000000000000000100001100000101",
			4279 => "11111111100010000100001100000101",
			4280 => "00000000000000000100001100000101",
			4281 => "00000000000000000100001100000101",
			4282 => "0000001000000000000111000100001100",
			4283 => "0000000001000000001011111100000100",
			4284 => "00000000000000000100001100000101",
			4285 => "0000001010000000000001010000000100",
			4286 => "00000000000000000100001100000101",
			4287 => "00000000011010000100001100000101",
			4288 => "00000000000000000100001100000101",
			4289 => "0000000100000000000000010100010100",
			4290 => "0000001011000000000000110100010000",
			4291 => "0000000111000000001011011100001100",
			4292 => "0000000001000000001011001100001000",
			4293 => "0000001000000000000101000100000100",
			4294 => "00000000000000000100001101001001",
			4295 => "11111111110010000100001101001001",
			4296 => "00000000000000000100001101001001",
			4297 => "00000000000000000100001101001001",
			4298 => "00000000000000000100001101001001",
			4299 => "0000001000000000001111001000001100",
			4300 => "0000000001000000001011111100000100",
			4301 => "00000000000000000100001101001001",
			4302 => "0000001000000000001001101000000100",
			4303 => "00000000000000000100001101001001",
			4304 => "00000000101001010100001101001001",
			4305 => "00000000000000000100001101001001",
			4306 => "0000001100000000001011011100011100",
			4307 => "0000001001000000000010101100001100",
			4308 => "0000001111000000001111101000000100",
			4309 => "00000000000000000100001110001101",
			4310 => "0000000110000000000100111100000100",
			4311 => "00000000000000000100001110001101",
			4312 => "11111111111100010100001110001101",
			4313 => "0000000110000000001000010000000100",
			4314 => "00000000000000000100001110001101",
			4315 => "0000001001000000001001000100001000",
			4316 => "0000001100000000001001110100000100",
			4317 => "00000000000000000100001110001101",
			4318 => "00000000001101110100001110001101",
			4319 => "00000000000000000100001110001101",
			4320 => "0000001011000000001111010000000100",
			4321 => "00000000000000000100001110001101",
			4322 => "11111110010000000100001110001101",
			4323 => "0000000111000000001000011000010100",
			4324 => "0000001100000000000100011000000100",
			4325 => "00000000000000000100001111100001",
			4326 => "0000000100000000001000001000000100",
			4327 => "00000000000000000100001111100001",
			4328 => "0000001000000000000111000000001000",
			4329 => "0000001111000000001000011100000100",
			4330 => "00000001010111100100001111100001",
			4331 => "00000000000000000100001111100001",
			4332 => "00000000000000000100001111100001",
			4333 => "0000001000000000000110001000001100",
			4334 => "0000001100000000001001110100000100",
			4335 => "00000000000000000100001111100001",
			4336 => "0000001100000000000100000100000100",
			4337 => "00000000001000000100001111100001",
			4338 => "00000000000000000100001111100001",
			4339 => "0000000110000000001000010000000100",
			4340 => "00000000000000000100001111100001",
			4341 => "0000000001000000001001100100000100",
			4342 => "11111111011101010100001111100001",
			4343 => "00000000000000000100001111100001",
			4344 => "0000000110000000001000010000011000",
			4345 => "0000000010000000001101101100000100",
			4346 => "00000000000000000100010000011101",
			4347 => "0000001010000000001000010100000100",
			4348 => "00000000000000000100010000011101",
			4349 => "0000001001000000001011001100000100",
			4350 => "00000000000000000100010000011101",
			4351 => "0000001100000000000001011000001000",
			4352 => "0000001100000000001010111000000100",
			4353 => "00000000000000000100010000011101",
			4354 => "00000001001010000100010000011101",
			4355 => "00000000000000000100010000011101",
			4356 => "0000001000000000001111001000000100",
			4357 => "00000000000000000100010000011101",
			4358 => "11111111110000010100010000011101",
			4359 => "0000001100000000001011011100011000",
			4360 => "0000000100000000001100001100000100",
			4361 => "00000000000000000100010001011001",
			4362 => "0000001001000000001011001100000100",
			4363 => "00000000000000000100010001011001",
			4364 => "0000000010000000000011110000001100",
			4365 => "0000000100000000000011110000000100",
			4366 => "00000000000000000100010001011001",
			4367 => "0000001100000000001010111000000100",
			4368 => "00000000000000000100010001011001",
			4369 => "00000000010111000100010001011001",
			4370 => "00000000000000000100010001011001",
			4371 => "0000001000000000000110001000000100",
			4372 => "00000000000000000100010001011001",
			4373 => "11111110101010000100010001011001",
			4374 => "0000000010000000001000000100010100",
			4375 => "0000000010000000001101101100000100",
			4376 => "00000000000000000100010010100101",
			4377 => "0000000110000000000101010000001100",
			4378 => "0000000001000000001001011000000100",
			4379 => "00000000000000000100010010100101",
			4380 => "0000000110000000001111000000000100",
			4381 => "00000000000000000100010010100101",
			4382 => "00000000000100010100010010100101",
			4383 => "00000000000000000100010010100101",
			4384 => "0000000001000000001101011000010000",
			4385 => "0000000000000000001010101100000100",
			4386 => "00000000000000000100010010100101",
			4387 => "0000000110000000000100111100000100",
			4388 => "00000000000000000100010010100101",
			4389 => "0000001010000000001000010100000100",
			4390 => "00000000000000000100010010100101",
			4391 => "11111111101100110100010010100101",
			4392 => "00000000000000000100010010100101",
			4393 => "0000001101000000001100111000011000",
			4394 => "0000001100000000000100011000000100",
			4395 => "00000000000000000100010011011001",
			4396 => "0000000110000000000100101100010000",
			4397 => "0000000010000000001101101100000100",
			4398 => "00000000000000000100010011011001",
			4399 => "0000000110000000001111000000000100",
			4400 => "00000000000000000100010011011001",
			4401 => "0000001011000000000110100000000100",
			4402 => "00000000001000100100010011011001",
			4403 => "00000000000000000100010011011001",
			4404 => "00000000000000000100010011011001",
			4405 => "11111111110011110100010011011001",
			4406 => "0000000010000000001000000100011000",
			4407 => "0000000110000000001001100100000100",
			4408 => "00000000000000000100010100100101",
			4409 => "0000001111000000001000110100010000",
			4410 => "0000000110000000000101010000001100",
			4411 => "0000001101000000001110101100000100",
			4412 => "00000000000000000100010100100101",
			4413 => "0000000010000000001100111000000100",
			4414 => "00000000000000000100010100100101",
			4415 => "00000000101101110100010100100101",
			4416 => "00000000000000000100010100100101",
			4417 => "00000000000000000100010100100101",
			4418 => "0000001100000000000111010000000100",
			4419 => "00000000000000000100010100100101",
			4420 => "0000000100000000000110001100000100",
			4421 => "00000000000000000100010100100101",
			4422 => "0000000110000000001000010000000100",
			4423 => "00000000000000000100010100100101",
			4424 => "11111111101001000100010100100101",
			4425 => "0000000100000000000100001100011100",
			4426 => "0000001011000000000000110100010100",
			4427 => "0000001000000000000101000100000100",
			4428 => "00000000000000000100010101111001",
			4429 => "0000001001000000000011101000001100",
			4430 => "0000001100000000001111011100001000",
			4431 => "0000000111000000000110110100000100",
			4432 => "11111111100010110100010101111001",
			4433 => "00000000000000000100010101111001",
			4434 => "00000000000000000100010101111001",
			4435 => "00000000000000000100010101111001",
			4436 => "0000001101000000001010000100000100",
			4437 => "00000000000110100100010101111001",
			4438 => "00000000000000000100010101111001",
			4439 => "0000001000000000001111001000001100",
			4440 => "0000001001000000000101010000000100",
			4441 => "00000000000000000100010101111001",
			4442 => "0000001100000000000101100100000100",
			4443 => "00000000111110100100010101111001",
			4444 => "00000000000000000100010101111001",
			4445 => "00000000000000000100010101111001",
			4446 => "0000000000000000001011000100100100",
			4447 => "0000000110000000000101010000011000",
			4448 => "0000001011000000000110100000001100",
			4449 => "0000001011000000000000110100000100",
			4450 => "00000000000000000100010111010101",
			4451 => "0000000110000000000101010000000100",
			4452 => "00000000100010100100010111010101",
			4453 => "00000000000000000100010111010101",
			4454 => "0000000110000000001000010000000100",
			4455 => "00000000000000000100010111010101",
			4456 => "0000000110000000001000010000000100",
			4457 => "11111111111000110100010111010101",
			4458 => "00000000000000000100010111010101",
			4459 => "0000001011000000001111010000001000",
			4460 => "0000001011000000000010001000000100",
			4461 => "00000000000000000100010111010101",
			4462 => "11111111110110100100010111010101",
			4463 => "00000000000000000100010111010101",
			4464 => "0000000000000000000000101000001000",
			4465 => "0000000010000000000110111100000100",
			4466 => "00000000000000000100010111010101",
			4467 => "00000010000010010100010111010101",
			4468 => "00000000000000000100010111010101",
			4469 => "0000000100000000000000010100100000",
			4470 => "0000001011000000000000110100010100",
			4471 => "0000001000000000000101000100000100",
			4472 => "00000000000000000100011000110001",
			4473 => "0000000001000000001010011000001100",
			4474 => "0000000111000000000110110100001000",
			4475 => "0000001010000000001000100100000100",
			4476 => "00000000000000000100011000110001",
			4477 => "11111111101100000100011000110001",
			4478 => "00000000000000000100011000110001",
			4479 => "00000000000000000100011000110001",
			4480 => "0000001010000000000001010000001000",
			4481 => "0000001010000000001000100100000100",
			4482 => "00000000000000000100011000110001",
			4483 => "00000000000001000100011000110001",
			4484 => "00000000000000000100011000110001",
			4485 => "0000001000000000001111001000001100",
			4486 => "0000000001000000001011111100000100",
			4487 => "00000000000000000100011000110001",
			4488 => "0000001000000000001001101000000100",
			4489 => "00000000000000000100011000110001",
			4490 => "00000000101111010100011000110001",
			4491 => "00000000000000000100011000110001",
			4492 => "0000000100000000000000010100010100",
			4493 => "0000000000000000001010101100000100",
			4494 => "00000000000000000100011010000101",
			4495 => "0000001001000000001000100100001100",
			4496 => "0000000111000000000111110000001000",
			4497 => "0000001010000000001000010100000100",
			4498 => "00000000000000000100011010000101",
			4499 => "11111111101000110100011010000101",
			4500 => "00000000000000000100011010000101",
			4501 => "00000000000000000100011010000101",
			4502 => "0000001010000000000101000100010100",
			4503 => "0000001001000000001011001100000100",
			4504 => "00000000000000000100011010000101",
			4505 => "0000000000000000000010011000000100",
			4506 => "00000000000000000100011010000101",
			4507 => "0000000110000000000100101100001000",
			4508 => "0000000111000000001011000000000100",
			4509 => "00000000000000000100011010000101",
			4510 => "00000000010110000100011010000101",
			4511 => "00000000000000000100011010000101",
			4512 => "00000000000000000100011010000101",
			4513 => "0000001101000000001010000100100000",
			4514 => "0000001100000000001001110100001000",
			4515 => "0000000100000000000000101100000100",
			4516 => "11111111111011110100011011010001",
			4517 => "00000000000000000100011011010001",
			4518 => "0000000100000000001110100100000100",
			4519 => "00000000000000000100011011010001",
			4520 => "0000001000000000000111000100010000",
			4521 => "0000001110000000001000011100001100",
			4522 => "0000001100000000000001011000001000",
			4523 => "0000000001000000001110010100000100",
			4524 => "00000000000000000100011011010001",
			4525 => "00000000110110000100011011010001",
			4526 => "00000000000000000100011011010001",
			4527 => "00000000000000000100011011010001",
			4528 => "00000000000000000100011011010001",
			4529 => "0000000001000000001101011000000100",
			4530 => "00000000000000000100011011010001",
			4531 => "11111111110100110100011011010001",
			4532 => "0000001101000000001010000100011100",
			4533 => "0000001001000000001001111100000100",
			4534 => "00000000000000000100011100011101",
			4535 => "0000000110000000001001111100010100",
			4536 => "0000000010000000000110111000000100",
			4537 => "00000000000000000100011100011101",
			4538 => "0000001100000000000100000100001100",
			4539 => "0000000010000000001010110100001000",
			4540 => "0000001100000000001001110100000100",
			4541 => "00000000000000000100011100011101",
			4542 => "00000000100010000100011100011101",
			4543 => "00000000000000000100011100011101",
			4544 => "00000000000000000100011100011101",
			4545 => "00000000000000000100011100011101",
			4546 => "0000001110000000000011010100001000",
			4547 => "0000000110000000001000010000000100",
			4548 => "00000000000000000100011100011101",
			4549 => "11111111111010110100011100011101",
			4550 => "00000000000000000100011100011101",
			4551 => "0000000100000000000011011000100100",
			4552 => "0000001000000000000110001000011000",
			4553 => "0000001001000000000111101100000100",
			4554 => "00000000000000000100011101111001",
			4555 => "0000001011000000000110100000010000",
			4556 => "0000001110000000001000011100001100",
			4557 => "0000000011000000000001011100000100",
			4558 => "00000000000000000100011101111001",
			4559 => "0000001011000000000100010000000100",
			4560 => "00000000000000000100011101111001",
			4561 => "00000000101100110100011101111001",
			4562 => "00000000000000000100011101111001",
			4563 => "00000000000000000100011101111001",
			4564 => "0000000100000000001001000000001000",
			4565 => "0000000011000000001110111000000100",
			4566 => "11111111011111110100011101111001",
			4567 => "00000000000000000100011101111001",
			4568 => "00000000000000000100011101111001",
			4569 => "0000001010000000000101000100001000",
			4570 => "0000000110000000001000010000000100",
			4571 => "00000000000000000100011101111001",
			4572 => "00000001101101100100011101111001",
			4573 => "00000000000000000100011101111001",
			4574 => "0000000100000000000100001100011100",
			4575 => "0000001000000000000101000100000100",
			4576 => "00000000000000000100011111001101",
			4577 => "0000000101000000001110110100010100",
			4578 => "0000001001000000000111110100010000",
			4579 => "0000000110000000000100111100000100",
			4580 => "00000000000000000100011111001101",
			4581 => "0000001011000000001101000100001000",
			4582 => "0000000000000000000001110100000100",
			4583 => "00000000000000000100011111001101",
			4584 => "11111111011100100100011111001101",
			4585 => "00000000000000000100011111001101",
			4586 => "00000000000000000100011111001101",
			4587 => "00000000000000000100011111001101",
			4588 => "0000001000000000000111000100001100",
			4589 => "0000001001000000000101010000000100",
			4590 => "00000000000000000100011111001101",
			4591 => "0000001010000000000001010000000100",
			4592 => "00000000000000000100011111001101",
			4593 => "00000000011011110100011111001101",
			4594 => "00000000000000000100011111001101",
			4595 => "0000001100000000001011011100100100",
			4596 => "0000000100000000000100001100001100",
			4597 => "0000000111000000001011011100001000",
			4598 => "0000001011000000001110101100000100",
			4599 => "11111111110100010100100000100001",
			4600 => "00000000000000000100100000100001",
			4601 => "00000000000000000100100000100001",
			4602 => "0000001010000000000101000100010100",
			4603 => "0000001001000000001011001100000100",
			4604 => "00000000000000000100100000100001",
			4605 => "0000000010000000001010110100001100",
			4606 => "0000001101000000001100000000001000",
			4607 => "0000000111000000001011000000000100",
			4608 => "00000000000000000100100000100001",
			4609 => "00000000010111010100100000100001",
			4610 => "00000000000000000100100000100001",
			4611 => "00000000000000000100100000100001",
			4612 => "00000000000000000100100000100001",
			4613 => "0000001000000000000110001000000100",
			4614 => "00000000000000000100100000100001",
			4615 => "11111110100100010100100000100001",
			4616 => "0000001111000000001111101000011000",
			4617 => "0000000001000000001001011000000100",
			4618 => "00000000000000000100100001111101",
			4619 => "0000000010000000001101101100000100",
			4620 => "00000000000000000100100001111101",
			4621 => "0000000110000000000101010000001100",
			4622 => "0000001100000000001010111000000100",
			4623 => "00000000000000000100100001111101",
			4624 => "0000000001000000001010011000000100",
			4625 => "00000000001010100100100001111101",
			4626 => "00000000000000000100100001111101",
			4627 => "00000000000000000100100001111101",
			4628 => "0000001000000000000001010100000100",
			4629 => "00000000000000000100100001111101",
			4630 => "0000001110000000000011010100010000",
			4631 => "0000001010000000001000010100000100",
			4632 => "00000000000000000100100001111101",
			4633 => "0000000000000000001010101100000100",
			4634 => "00000000000000000100100001111101",
			4635 => "0000000011000000000011101100000100",
			4636 => "11111111101100100100100001111101",
			4637 => "00000000000000000100100001111101",
			4638 => "00000000000000000100100001111101",
			4639 => "0000000010000000001011110000011000",
			4640 => "0000000010000000001101101100000100",
			4641 => "00000000000000000100100011110001",
			4642 => "0000000110000000001000010000010000",
			4643 => "0000000110000000001111000000000100",
			4644 => "00000000000000000100100011110001",
			4645 => "0000001100000000001010111000000100",
			4646 => "00000000000000000100100011110001",
			4647 => "0000000000000000000001110100000100",
			4648 => "00000000000000000100100011110001",
			4649 => "00000001011001000100100011110001",
			4650 => "00000000000000000100100011110001",
			4651 => "0000001000000000001111001000011000",
			4652 => "0000000000000000000111000000001100",
			4653 => "0000000000000000001010101100000100",
			4654 => "00000000000000000100100011110001",
			4655 => "0000000000000000000111000000000100",
			4656 => "11111111111101000100100011110001",
			4657 => "00000000000000000100100011110001",
			4658 => "0000001011000000000100010000000100",
			4659 => "00000000000000000100100011110001",
			4660 => "0000001011000000000111100000000100",
			4661 => "00000000000110000100100011110001",
			4662 => "00000000000000000100100011110001",
			4663 => "0000001110000000000011010100001000",
			4664 => "0000000011000000000011101100000100",
			4665 => "11111111110001110100100011110001",
			4666 => "00000000000000000100100011110001",
			4667 => "00000000000000000100100011110001",
			4668 => "0000000100000000000011011000101000",
			4669 => "0000000001000000001010011000011000",
			4670 => "0000001000000000000101000100000100",
			4671 => "00000000000000000100100101010101",
			4672 => "0000000100000000000111011100010000",
			4673 => "0000001011000000000110100000001100",
			4674 => "0000000101000000000110010000001000",
			4675 => "0000001001000000000011101000000100",
			4676 => "11111111100000000100100101010101",
			4677 => "00000000000000000100100101010101",
			4678 => "00000000000000000100100101010101",
			4679 => "00000000000000000100100101010101",
			4680 => "00000000000000000100100101010101",
			4681 => "0000001011000000001110101000001100",
			4682 => "0000001000000000000110001000001000",
			4683 => "0000001011000000001010010100000100",
			4684 => "00000000000000000100100101010101",
			4685 => "00000000001100110100100101010101",
			4686 => "00000000000000000100100101010101",
			4687 => "00000000000000000100100101010101",
			4688 => "0000001010000000000101000100001000",
			4689 => "0000000001000000001001011000000100",
			4690 => "00000000000000000100100101010101",
			4691 => "00000001001010000100100101010101",
			4692 => "00000000000000000100100101010101",
			4693 => "0000001001000000001010100000001000",
			4694 => "0000001111000000001110100100000100",
			4695 => "11111111100010010100100110110001",
			4696 => "00000000000000000100100110110001",
			4697 => "0000001110000000001000011100011000",
			4698 => "0000000110000000001001111100010100",
			4699 => "0000001011000000000100010000000100",
			4700 => "00000000000000000100100110110001",
			4701 => "0000000011000000001100001100001100",
			4702 => "0000001011000000000110100000001000",
			4703 => "0000000101000000001001010000000100",
			4704 => "00000000000000000100100110110001",
			4705 => "00000000110111100100100110110001",
			4706 => "00000000000000000100100110110001",
			4707 => "00000000000000000100100110110001",
			4708 => "00000000000000000100100110110001",
			4709 => "0000001001000000001000100100001100",
			4710 => "0000000111000000000111110000001000",
			4711 => "0000000100000000000100001100000100",
			4712 => "11111111101101100100100110110001",
			4713 => "00000000000000000100100110110001",
			4714 => "00000000000000000100100110110001",
			4715 => "00000000000000000100100110110001",
			4716 => "0000000101000000001110000100010000",
			4717 => "0000001100000000001010111000000100",
			4718 => "00000000000000000100101000011101",
			4719 => "0000000100000000001111100000000100",
			4720 => "00000000000000000100101000011101",
			4721 => "0000001000000000001101010000000100",
			4722 => "00000001101111000100101000011101",
			4723 => "00000000000000000100101000011101",
			4724 => "0000000001000000001010011000011000",
			4725 => "0000000110000000000100111100000100",
			4726 => "00000000000000000100101000011101",
			4727 => "0000000111000000001111011100000100",
			4728 => "00000000000000000100101000011101",
			4729 => "0000001001000000000011101000001100",
			4730 => "0000000101000000001110110100001000",
			4731 => "0000001000000000000101000100000100",
			4732 => "00000000000000000100101000011101",
			4733 => "11111111100000010100101000011101",
			4734 => "00000000000000000100101000011101",
			4735 => "00000000000000000100101000011101",
			4736 => "0000000110000000000100101100001100",
			4737 => "0000000111000000000111010000000100",
			4738 => "00000000000000000100101000011101",
			4739 => "0000000000000000001010101100000100",
			4740 => "00000000000000000100101000011101",
			4741 => "00000000010101110100101000011101",
			4742 => "00000000000000000100101000011101",
			4743 => "0000000000000000001011000100110000",
			4744 => "0000001100000000000111010000100000",
			4745 => "0000000101000000000111111100001100",
			4746 => "0000000010000000000110111000001000",
			4747 => "0000000000000000000001110100000100",
			4748 => "00000000000000000100101010001001",
			4749 => "11111111110001110100101010001001",
			4750 => "00000000000000000100101010001001",
			4751 => "0000000110000000000100101100010000",
			4752 => "0000001101000000001111010100001100",
			4753 => "0000000001000000001101111100000100",
			4754 => "00000000000000000100101010001001",
			4755 => "0000000011000000000010111000000100",
			4756 => "00000000101000000100101010001001",
			4757 => "00000000000000000100101010001001",
			4758 => "00000000000000000100101010001001",
			4759 => "00000000000000000100101010001001",
			4760 => "0000000010000000001000000100000100",
			4761 => "00000000000000000100101010001001",
			4762 => "0000001001000000001000100100001000",
			4763 => "0000000110000000001000010000000100",
			4764 => "00000000000000000100101010001001",
			4765 => "11111111101000110100101010001001",
			4766 => "00000000000000000100101010001001",
			4767 => "0000000000000000000000101000000100",
			4768 => "00000001001110010100101010001001",
			4769 => "00000000000000000100101010001001",
			4770 => "0000000010000000001011110000011100",
			4771 => "0000000010000000001101101100000100",
			4772 => "00000000000000000100101011111101",
			4773 => "0000000110000000001000010000010100",
			4774 => "0000000110000000001111000000000100",
			4775 => "00000000000000000100101011111101",
			4776 => "0000001100000000001010111000000100",
			4777 => "00000000000000000100101011111101",
			4778 => "0000000100000000000110111000000100",
			4779 => "00000000000000000100101011111101",
			4780 => "0000001010000000001000100100000100",
			4781 => "00000000000000000100101011111101",
			4782 => "00000001100010000100101011111101",
			4783 => "00000000000000000100101011111101",
			4784 => "0000001101000000001100000000001100",
			4785 => "0000001001000000000100101100000100",
			4786 => "00000000000000000100101011111101",
			4787 => "0000000001000000000111101000000100",
			4788 => "00000000000000000100101011111101",
			4789 => "00000000000101000100101011111101",
			4790 => "0000001001000000001000100100010000",
			4791 => "0000000110000000001000010000000100",
			4792 => "00000000000000000100101011111101",
			4793 => "0000001000000000000001010100000100",
			4794 => "00000000000000000100101011111101",
			4795 => "0000000100000000001110100100000100",
			4796 => "00000000000000000100101011111101",
			4797 => "11111111100100110100101011111101",
			4798 => "00000000000000000100101011111101",
			4799 => "0000000001000000001100011000100100",
			4800 => "0000001001000000001010100000010000",
			4801 => "0000000001000000001011111100000100",
			4802 => "11111110010111010100101110010001",
			4803 => "0000000010000000001110000000000100",
			4804 => "11111110011000010100101110010001",
			4805 => "0000001110000000001011101100000100",
			4806 => "00000001111000010100101110010001",
			4807 => "11111110011001000100101110010001",
			4808 => "0000000111000000001111011100000100",
			4809 => "11111110010111110100101110010001",
			4810 => "0000001110000000000010010100001000",
			4811 => "0000000001000000000100110100000100",
			4812 => "00000011000001000100101110010001",
			4813 => "00000001010001110100101110010001",
			4814 => "0000001100000000001000011000000100",
			4815 => "11111110010100110100101110010001",
			4816 => "00000000000000000100101110010001",
			4817 => "0000001101000000001100010100001100",
			4818 => "0000001110000000001101101100001000",
			4819 => "0000000111000000001000011000000100",
			4820 => "11111111000110100100101110010001",
			4821 => "00000000100111110100101110010001",
			4822 => "11111110011001100100101110010001",
			4823 => "0000001010000000001100011100010100",
			4824 => "0000000111000000000111010000000100",
			4825 => "00000000011010000100101110010001",
			4826 => "0000001100000000000101100100001100",
			4827 => "0000001011000000001110101000001000",
			4828 => "0000001001000000001010100100000100",
			4829 => "00000001011101110100101110010001",
			4830 => "00000001111000110100101110010001",
			4831 => "00000000111101110100101110010001",
			4832 => "00000000010111110100101110010001",
			4833 => "0000000101000000001100010000000100",
			4834 => "11111110100110010100101110010001",
			4835 => "00000000100110100100101110010001",
			4836 => "0000001001000000001010100100100000",
			4837 => "0000001001000000001010100100010100",
			4838 => "0000001001000000001001111100000100",
			4839 => "11111110010110110100110000010101",
			4840 => "0000000111000000000001101000000100",
			4841 => "11111110010111110100110000010101",
			4842 => "0000001110000000001111101000001000",
			4843 => "0000000010000000001110000000000100",
			4844 => "11111110011011000100110000010101",
			4845 => "00000010011100110100110000010101",
			4846 => "11111110011001010100110000010101",
			4847 => "0000000101000000000101110000000100",
			4848 => "11111110010111110100110000010101",
			4849 => "0000000011000000001011110000000100",
			4850 => "00000010100011010100110000010101",
			4851 => "11111111100011100100110000010101",
			4852 => "0000001011000000000101110100000100",
			4853 => "11111110011000100100110000010101",
			4854 => "0000001000000000000110001000011000",
			4855 => "0000000111000000000111010000001000",
			4856 => "0000000101000000000101110000000100",
			4857 => "11111110100111010100110000010101",
			4858 => "00000000111100000100110000010101",
			4859 => "0000001100000000000101100100001100",
			4860 => "0000001011000000001110101000001000",
			4861 => "0000001001000000001010100100000100",
			4862 => "00000001100001110100110000010101",
			4863 => "00000001111110000100110000010101",
			4864 => "00000001000110110100110000010101",
			4865 => "00000000011110110100110000010101",
			4866 => "0000000100000000000111011100000100",
			4867 => "11111110100111010100110000010101",
			4868 => "00000000110010100100110000010101",
			4869 => "0000000001000000000100110100101100",
			4870 => "0000001001000000001010100100011100",
			4871 => "0000000001000000000101011100000100",
			4872 => "11111110010110010100110010100001",
			4873 => "0000000100000000000011110100010000",
			4874 => "0000000100000000001110111000000100",
			4875 => "11111110010110110100110010100001",
			4876 => "0000000100000000001110111000000100",
			4877 => "00000001100100010100110010100001",
			4878 => "0000001011000000001011110100000100",
			4879 => "00000000000000000100110010100001",
			4880 => "11111110011011110100110010100001",
			4881 => "0000001100000000001000011000000100",
			4882 => "00000011001110000100110010100001",
			4883 => "11111110011111010100110010100001",
			4884 => "0000000111000000000111010000001000",
			4885 => "0000001100000000001001110100000100",
			4886 => "11111110011001000100110010100001",
			4887 => "00000000001101000100110010100001",
			4888 => "0000001110000000001011110000000100",
			4889 => "00000010110110110100110010100001",
			4890 => "00000000001100100100110010100001",
			4891 => "0000001101000000001100010100000100",
			4892 => "11111110010101010100110010100001",
			4893 => "0000000110000000000100101100010100",
			4894 => "0000001100000000001001110100000100",
			4895 => "00000000101110010100110010100001",
			4896 => "0000000110000000000100101100001100",
			4897 => "0000000100000000001111100000001000",
			4898 => "0000000110000000000101010000000100",
			4899 => "00000010000100110100110010100001",
			4900 => "00000001100000010100110010100001",
			4901 => "00000011001001110100110010100001",
			4902 => "00000000100110010100110010100001",
			4903 => "11111110011111100100110010100001",
			4904 => "0000000001000000001100011000110000",
			4905 => "0000001001000000001010100100101000",
			4906 => "0000001001000000001010100100011100",
			4907 => "0000000110000000000100111100000100",
			4908 => "11011011100010000100110100111101",
			4909 => "0000001111000000001110000000010000",
			4910 => "0000000010000000001110000000001000",
			4911 => "0000000111000000001000011000000100",
			4912 => "11011011101001110100110100111101",
			4913 => "11011100111111010100110100111101",
			4914 => "0000000001000000001011111100000100",
			4915 => "11011011110001000100110100111101",
			4916 => "11100101111111000100110100111101",
			4917 => "0000000110000000001000010000000100",
			4918 => "11011100100100100100110100111101",
			4919 => "11011011100010100100110100111101",
			4920 => "0000001100000000000001101000001000",
			4921 => "0000000101000000001001010000000100",
			4922 => "11011011100011000100110100111101",
			4923 => "11011101100001010100110100111101",
			4924 => "11100011101010010100110100111101",
			4925 => "0000000110000000001000010000000100",
			4926 => "11101010011111110100110100111101",
			4927 => "11011011101001100100110100111101",
			4928 => "0000000101000000000111111100001000",
			4929 => "0000000111000000000111010000000100",
			4930 => "11011011100011010100110100111101",
			4931 => "11100011101101000100110100111101",
			4932 => "0000001000000000001111001000010000",
			4933 => "0000000111000000000000011100001000",
			4934 => "0000001010000000001001000100000100",
			4935 => "11101010101000000100110100111101",
			4936 => "11100100011110110100110100111101",
			4937 => "0000001100000000001011011100000100",
			4938 => "11101011010000010100110100111101",
			4939 => "11100111011111010100110100111101",
			4940 => "0000000110000000000100101100000100",
			4941 => "11011111100101100100110100111101",
			4942 => "11011011101101100100110100111101",
			4943 => "0000001100000000001001110100001000",
			4944 => "0000001010000000000110011100000100",
			4945 => "11111111011101100100110111000001",
			4946 => "00000000000000000100110111000001",
			4947 => "0000001101000000000110111100100000",
			4948 => "0000000001000000001100011000011000",
			4949 => "0000001101000000001110110100010000",
			4950 => "0000001101000000001010001000000100",
			4951 => "00000000000000000100110111000001",
			4952 => "0000000000000000001110111100001000",
			4953 => "0000000000000000001111001000000100",
			4954 => "00000000000000000100110111000001",
			4955 => "00000000001101000100110111000001",
			4956 => "00000000000000000100110111000001",
			4957 => "0000000000000000001010101100000100",
			4958 => "00000000000000000100110111000001",
			4959 => "11111111111000110100110111000001",
			4960 => "0000001011000000000001001000000100",
			4961 => "00000000000000000100110111000001",
			4962 => "00000000101011110100110111000001",
			4963 => "0000001001000000000011101000001000",
			4964 => "0000001100000000000100000100000100",
			4965 => "00000000000100100100110111000001",
			4966 => "00000000000000000100110111000001",
			4967 => "0000001100000000000111010000010000",
			4968 => "0000000101000000001110110100001100",
			4969 => "0000000011000000000101000000000100",
			4970 => "00000000000000000100110111000001",
			4971 => "0000000001000000001111000000000100",
			4972 => "11111111010100000100110111000001",
			4973 => "00000000000000000100110111000001",
			4974 => "00000000000000000100110111000001",
			4975 => "00000000000000000100110111000001",
			4976 => "0000001100000000001011000000000100",
			4977 => "11111110110001000100111000110101",
			4978 => "0000000110000000001000010000001100",
			4979 => "0000001111000000000010010100000100",
			4980 => "00000000000000000100111000110101",
			4981 => "0000000001000000000100110100000100",
			4982 => "00000000000000000100111000110101",
			4983 => "00000000110100010100111000110101",
			4984 => "0000000000000000001010101100010000",
			4985 => "0000001111000000001000110100000100",
			4986 => "00000000000000000100111000110101",
			4987 => "0000001100000000000111010000001000",
			4988 => "0000000000000000001010101100000100",
			4989 => "00000000000000000100111000110101",
			4990 => "11111111000111000100111000110101",
			4991 => "00000000000000000100111000110101",
			4992 => "0000000110000000000101010000010000",
			4993 => "0000000100000000001100001100000100",
			4994 => "00000000000000000100111000110101",
			4995 => "0000000001000000001011111100000100",
			4996 => "00000000000000000100111000110101",
			4997 => "0000001110000000000110001100000100",
			4998 => "00000000111100010100111000110101",
			4999 => "00000000000000000100111000110101",
			5000 => "0000000001000000001010011000000100",
			5001 => "11111111010011010100111000110101",
			5002 => "0000000110000000000100101100000100",
			5003 => "00000000010011010100111000110101",
			5004 => "11111111100101100100111000110101",
			5005 => "0000000001000000000100110100110100",
			5006 => "0000001001000000001010100100100100",
			5007 => "0000000001000000000101011100000100",
			5008 => "11111110010101110100111011001001",
			5009 => "0000000100000000000011110100010000",
			5010 => "0000000100000000001110111000000100",
			5011 => "11111110010110010100111011001001",
			5012 => "0000000100000000001110111000000100",
			5013 => "00000001101110110100111011001001",
			5014 => "0000001011000000001011110100000100",
			5015 => "00000000000000000100111011001001",
			5016 => "11111110011010010100111011001001",
			5017 => "0000000010000000000110001100000100",
			5018 => "00000100110100110100111011001001",
			5019 => "0000000100000000001011100000001000",
			5020 => "0000000101000000000010000100000100",
			5021 => "00000001010010000100111011001001",
			5022 => "11111111100011110100111011001001",
			5023 => "11111110011101100100111011001001",
			5024 => "0000000111000000000111010000001000",
			5025 => "0000001100000000001001110100000100",
			5026 => "11111110011000000100111011001001",
			5027 => "00000000001001100100111011001001",
			5028 => "0000001110000000001011110000000100",
			5029 => "00000011001010100100111011001001",
			5030 => "00000000001011100100111011001001",
			5031 => "0000001101000000001100010100000100",
			5032 => "11111110010100010100111011001001",
			5033 => "0000001000000000000001110100010000",
			5034 => "0000001100000000001001110100000100",
			5035 => "00000000110111110100111011001001",
			5036 => "0000001000000000001111001000001000",
			5037 => "0000001100000000001011011100000100",
			5038 => "00000010001101010100111011001001",
			5039 => "00000001011101000100111011001001",
			5040 => "00000001010001010100111011001001",
			5041 => "11111110100100000100111011001001",
			5042 => "0000000001000000001100011000100100",
			5043 => "0000000001000000000101011100000100",
			5044 => "11111110011000000100111101110101",
			5045 => "0000000100000000000100001100010100",
			5046 => "0000000111000000000000011100001000",
			5047 => "0000000101000000001110010000000100",
			5048 => "11111110010110100100111101110101",
			5049 => "11111111110100110100111101110101",
			5050 => "0000000110000000001000010000001000",
			5051 => "0000000001000000001101111100000100",
			5052 => "11111110110100010100111101110101",
			5053 => "00000001111010110100111101110101",
			5054 => "11111110011001010100111101110101",
			5055 => "0000000010000000000110001100000100",
			5056 => "00000011100000100100111101110101",
			5057 => "0000000110000000000101010000000100",
			5058 => "00000001011100000100111101110101",
			5059 => "11111110011000010100111101110101",
			5060 => "0000001100000000001001110100001100",
			5061 => "0000001010000000001001000100001000",
			5062 => "0000000100000000001100001100000100",
			5063 => "11111110000010000100111101110101",
			5064 => "00000001001110100100111101110101",
			5065 => "11111110001010000100111101110101",
			5066 => "0000000110000000000100101100100000",
			5067 => "0000001011000000000001001000001100",
			5068 => "0000001110000000000110111000000100",
			5069 => "00000010000010000100111101110101",
			5070 => "0000001001000000000011101000000100",
			5071 => "11111110010011110100111101110101",
			5072 => "00000001101001100100111101110101",
			5073 => "0000000110000000001001111100001100",
			5074 => "0000001011000000000110100000000100",
			5075 => "00000001110010100100111101110101",
			5076 => "0000001011000000001101000100000100",
			5077 => "00000001001000110100111101110101",
			5078 => "00000001101100110100111101110101",
			5079 => "0000000001000000001011001100000100",
			5080 => "11111111001101100100111101110101",
			5081 => "00000001111010010100111101110101",
			5082 => "0000000100000000000011011000000100",
			5083 => "11111110111001010100111101110101",
			5084 => "00000000001101110100111101110101",
			5085 => "0000000001000000000111101000000100",
			5086 => "11111110111011100100111111110001",
			5087 => "0000000100000000000011110000100100",
			5088 => "0000001011000000000000110100010000",
			5089 => "0000001000000000000101000100000100",
			5090 => "00000000000000000100111111110001",
			5091 => "0000000001000000001010011000001000",
			5092 => "0000001100000000001111011100000100",
			5093 => "11111110111100100100111111110001",
			5094 => "00000000000000000100111111110001",
			5095 => "00000000000000000100111111110001",
			5096 => "0000000011000000001100001100001100",
			5097 => "0000001011000000001101000100001000",
			5098 => "0000001010000000001001000100000100",
			5099 => "00000000101101110100111111110001",
			5100 => "00000000000000000100111111110001",
			5101 => "00000000000000000100111111110001",
			5102 => "0000001010000000001000010100000100",
			5103 => "11111111101110010100111111110001",
			5104 => "00000000000000000100111111110001",
			5105 => "0000000110000000000100101100010100",
			5106 => "0000001100000000001011011100010000",
			5107 => "0000001100000000001001110100000100",
			5108 => "00000000000000000100111111110001",
			5109 => "0000001110000000000110001100001000",
			5110 => "0000000001000000000100110100000100",
			5111 => "00000000000000000100111111110001",
			5112 => "00000000111100010100111111110001",
			5113 => "00000000000000000100111111110001",
			5114 => "00000000000000000100111111110001",
			5115 => "11111111110010000100111111110001",
			5116 => "0000000010000000000011000000001000",
			5117 => "0000001011000000000001001000000100",
			5118 => "11111110100110100101000010001101",
			5119 => "00000000000000000101000010001101",
			5120 => "0000000110000000000101010000101100",
			5121 => "0000001101000000001111010100011100",
			5122 => "0000000001000000001010011000011000",
			5123 => "0000001110000000000110111000001100",
			5124 => "0000001001000000000100111100000100",
			5125 => "00000000000000000101000010001101",
			5126 => "0000000100000000001000001000000100",
			5127 => "00000000000000000101000010001101",
			5128 => "00000000111000000101000010001101",
			5129 => "0000000111000000001011011100001000",
			5130 => "0000000000000000000010011000000100",
			5131 => "11111111000010010101000010001101",
			5132 => "00000000000000000101000010001101",
			5133 => "00000000000000000101000010001101",
			5134 => "00000001010000100101000010001101",
			5135 => "0000001001000000000011101000001000",
			5136 => "0000000001000000001100011000000100",
			5137 => "00000000000000000101000010001101",
			5138 => "00000000011111000101000010001101",
			5139 => "0000000000000000000111000000000100",
			5140 => "11111110111010100101000010001101",
			5141 => "00000000000000000101000010001101",
			5142 => "0000001001000000001000100100001100",
			5143 => "0000000100000000000011101100001000",
			5144 => "0000001010000000000110011000000100",
			5145 => "00000000000000000101000010001101",
			5146 => "11111110111000010101000010001101",
			5147 => "00000000000000000101000010001101",
			5148 => "0000001001000000001000010100001000",
			5149 => "0000000001000000001001100100000100",
			5150 => "00000000000000000101000010001101",
			5151 => "00000000101000000101000010001101",
			5152 => "0000001010000000000110011100000100",
			5153 => "00000000000000000101000010001101",
			5154 => "11111111111001100101000010001101",
			5155 => "0000000001000000000101011100000100",
			5156 => "11111110110010010101000100001001",
			5157 => "0000000110000000000101010000101100",
			5158 => "0000001001000000000011101000011000",
			5159 => "0000001001000000001010100100010000",
			5160 => "0000000000000000000010011000001100",
			5161 => "0000000110000000000100111100000100",
			5162 => "00000000000000000101000100001001",
			5163 => "0000000001000000001100011000000100",
			5164 => "11111111100010110101000100001001",
			5165 => "00000000000000000101000100001001",
			5166 => "00000000101100010101000100001001",
			5167 => "0000001101000000001100010100000100",
			5168 => "00000000000000000101000100001001",
			5169 => "00000001000101100101000100001001",
			5170 => "0000001010000000001000010100010000",
			5171 => "0000001110000000001110000000000100",
			5172 => "00000000000000000101000100001001",
			5173 => "0000001100000000001010001100001000",
			5174 => "0000001101000000000111011000000100",
			5175 => "00000000000000000101000100001001",
			5176 => "11111110111000110101000100001001",
			5177 => "00000000000000000101000100001001",
			5178 => "00000000101011100101000100001001",
			5179 => "0000000111000000001111011100000100",
			5180 => "00000000000000000101000100001001",
			5181 => "0000000001000000001101011000000100",
			5182 => "11111111001010000101000100001001",
			5183 => "0000001000000000000111000100000100",
			5184 => "00000000010100000101000100001001",
			5185 => "11111111101101100101000100001001",
			5186 => "0000000010000000000011000000001100",
			5187 => "0000001000000000000101000100000100",
			5188 => "00000000000000000101000110011101",
			5189 => "0000001111000000001111101000000100",
			5190 => "11111111010100100101000110011101",
			5191 => "00000000000000000101000110011101",
			5192 => "0000000101000000000110010000011000",
			5193 => "0000000110000000001001111100010100",
			5194 => "0000001001000000000100111100000100",
			5195 => "00000000000000000101000110011101",
			5196 => "0000001111000000000010111000001100",
			5197 => "0000000100000000001110100100000100",
			5198 => "00000000000000000101000110011101",
			5199 => "0000000110000000000100111100000100",
			5200 => "00000000000000000101000110011101",
			5201 => "00000000101101010101000110011101",
			5202 => "00000000000000000101000110011101",
			5203 => "00000000000000000101000110011101",
			5204 => "0000000111000000000100010000010100",
			5205 => "0000001001000000000011101000000100",
			5206 => "00000000000000000101000110011101",
			5207 => "0000000011000000000101000000000100",
			5208 => "00000000000000000101000110011101",
			5209 => "0000001011000000001101000100001000",
			5210 => "0000001101000000000110111100000100",
			5211 => "00000000000000000101000110011101",
			5212 => "11111111010010010101000110011101",
			5213 => "00000000000000000101000110011101",
			5214 => "0000000110000000000100101100010000",
			5215 => "0000001111000000001000011100000100",
			5216 => "00000000000000000101000110011101",
			5217 => "0000001110000000001011110000000100",
			5218 => "00000000000000000101000110011101",
			5219 => "0000001001000000001010100100000100",
			5220 => "00000000000000000101000110011101",
			5221 => "00000000110100000101000110011101",
			5222 => "11111111111000100101000110011101",
			5223 => "0000001001000000000100101100001000",
			5224 => "0000000100000000001100111100000100",
			5225 => "11111110101000100101001000100001",
			5226 => "00000000000000000101001000100001",
			5227 => "0000000111000000000111010000001000",
			5228 => "0000000000000000000010111100000100",
			5229 => "11111111010000110101001000100001",
			5230 => "00000000000000000101001000100001",
			5231 => "0000001011000000000110100000011000",
			5232 => "0000001100000000000100000100010000",
			5233 => "0000001110000000001000001000001100",
			5234 => "0000000000000000000001110100000100",
			5235 => "00000000000000000101001000100001",
			5236 => "0000001001000000000111101100000100",
			5237 => "00000000000000000101001000100001",
			5238 => "00000001000111100101001000100001",
			5239 => "00000000000000000101001000100001",
			5240 => "0000001001000000000010101100000100",
			5241 => "11111111111111010101001000100001",
			5242 => "00000000000000000101001000100001",
			5243 => "0000001110000000001110000000001000",
			5244 => "0000000100000000001100001100000100",
			5245 => "00000000000000000101001000100001",
			5246 => "11111111010001110101001000100001",
			5247 => "0000000110000000000100101100010000",
			5248 => "0000000111000000000100010000001000",
			5249 => "0000000111000000000010001000000100",
			5250 => "00000000000000000101001000100001",
			5251 => "11111111110111000101001000100001",
			5252 => "0000000001000000001100011000000100",
			5253 => "00000000000000000101001000100001",
			5254 => "00000001000011110101001000100001",
			5255 => "11111111101000000101001000100001",
			5256 => "0000001100000000001011000000000100",
			5257 => "11111111010100110101001010011101",
			5258 => "0000000110000000001001111100110000",
			5259 => "0000000100000000000011110000011100",
			5260 => "0000001011000000000000110100010000",
			5261 => "0000000110000000000100111100000100",
			5262 => "00000000000000000101001010011101",
			5263 => "0000000001000000001010011000001000",
			5264 => "0000001100000000001111011100000100",
			5265 => "11111111001011010101001010011101",
			5266 => "00000000000000000101001010011101",
			5267 => "00000000000000000101001010011101",
			5268 => "0000001011000000000110100000001000",
			5269 => "0000000001000000000100110100000100",
			5270 => "00000000000000000101001010011101",
			5271 => "00000000011100110101001010011101",
			5272 => "00000000000000000101001010011101",
			5273 => "0000001110000000001000001000010000",
			5274 => "0000001001000000000101010000000100",
			5275 => "00000000000000000101001010011101",
			5276 => "0000000111000000000001101000000100",
			5277 => "00000000000000000101001010011101",
			5278 => "0000000001000000001011111100000100",
			5279 => "00000000000000000101001010011101",
			5280 => "00000000101100110101001010011101",
			5281 => "00000000000000000101001010011101",
			5282 => "0000000001000000001001100100000100",
			5283 => "11111111011101000101001010011101",
			5284 => "0000001000000000000111000100000100",
			5285 => "00000000000101110101001010011101",
			5286 => "00000000000000000101001010011101",
			5287 => "0000001100000000001011000000000100",
			5288 => "11111110101111000101001100100001",
			5289 => "0000000110000000001000010000010000",
			5290 => "0000000011000000000001011100000100",
			5291 => "00000000000000000101001100100001",
			5292 => "0000000001000000000100110100000100",
			5293 => "00000000000000000101001100100001",
			5294 => "0000001111000000000010010100000100",
			5295 => "00000000000000000101001100100001",
			5296 => "00000000111000100101001100100001",
			5297 => "0000000000000000001010101100010000",
			5298 => "0000001111000000001000110100000100",
			5299 => "00000000000000000101001100100001",
			5300 => "0000001100000000000111010000001000",
			5301 => "0000001000000000000001010100000100",
			5302 => "00000000000000000101001100100001",
			5303 => "11111111000000110101001100100001",
			5304 => "00000000000000000101001100100001",
			5305 => "0000000110000000000101010000010000",
			5306 => "0000001010000000001000010100000100",
			5307 => "00000000000000000101001100100001",
			5308 => "0000000001000000001011111100000100",
			5309 => "00000000000000000101001100100001",
			5310 => "0000001111000000000011001100000100",
			5311 => "00000000111101100101001100100001",
			5312 => "00000000000000000101001100100001",
			5313 => "0000000001000000001010011000000100",
			5314 => "11111111010000010101001100100001",
			5315 => "0000000110000000000100101100001000",
			5316 => "0000000000000000000011010000000100",
			5317 => "00000000011110000101001100100001",
			5318 => "00000000000000000101001100100001",
			5319 => "11111111100011000101001100100001",
			5320 => "0000001001000000000100111100000100",
			5321 => "11111110100100010101001110110101",
			5322 => "0000000110000000000101010000110000",
			5323 => "0000000000000000000111000000100000",
			5324 => "0000000011000000001100001100011000",
			5325 => "0000000111000000000001011000001100",
			5326 => "0000000100000000001110100100001000",
			5327 => "0000001011000000000000110100000100",
			5328 => "11111110111010110101001110110101",
			5329 => "00000000000000000101001110110101",
			5330 => "00000000000000000101001110110101",
			5331 => "0000000111000000000101110100001000",
			5332 => "0000000001000000000100110100000100",
			5333 => "00000000000000000101001110110101",
			5334 => "00000001001100110101001110110101",
			5335 => "00000000000000000101001110110101",
			5336 => "0000001001000000000011101000000100",
			5337 => "00000000000000000101001110110101",
			5338 => "11111110101010010101001110110101",
			5339 => "0000000100000000000110001100000100",
			5340 => "00000000000000000101001110110101",
			5341 => "0000001111000000001101001000001000",
			5342 => "0000001111000000001111100100000100",
			5343 => "00000000000000000101001110110101",
			5344 => "00000001000000110101001110110101",
			5345 => "00000000000000000101001110110101",
			5346 => "0000001001000000001000100100001100",
			5347 => "0000000100000000000011101100001000",
			5348 => "0000001000000000001100000100000100",
			5349 => "00000000000000000101001110110101",
			5350 => "11111110110101100101001110110101",
			5351 => "00000000000000000101001110110101",
			5352 => "0000001000000000000111000100001000",
			5353 => "0000001100000000001000011000000100",
			5354 => "00000000000000000101001110110101",
			5355 => "00000000111001010101001110110101",
			5356 => "11111111111100100101001110110101",
			5357 => "0000000001000000000100110100101000",
			5358 => "0000000110000000000100111100000100",
			5359 => "11111110011001100101010010010001",
			5360 => "0000001111000000000110111000010000",
			5361 => "0000000100000000000111011100001000",
			5362 => "0000000011000000001100111000000100",
			5363 => "11111110101111100101010010010001",
			5364 => "00000000000000000101010010010001",
			5365 => "0000001001000000001011001100000100",
			5366 => "11111111100100010101010010010001",
			5367 => "00000001111101000101010010010001",
			5368 => "0000000110000000001000010000001000",
			5369 => "0000000110000000001000010000000100",
			5370 => "11111111011110110101010010010001",
			5371 => "00000000100011000101010010010001",
			5372 => "0000000011000000001000101000001000",
			5373 => "0000000011000000000001011100000100",
			5374 => "11111111100111000101010010010001",
			5375 => "00000000000000000101010010010001",
			5376 => "11111110100010000101010010010001",
			5377 => "0000000001000000001100011000100100",
			5378 => "0000000110000000000100111100010000",
			5379 => "0000000011000000000001011100000100",
			5380 => "11111110110100010101010010010001",
			5381 => "0000001111000000000010010100001000",
			5382 => "0000000010000000001111101000000100",
			5383 => "00000001010000010101010010010001",
			5384 => "11111111101100100101010010010001",
			5385 => "00000001111101010101010010010001",
			5386 => "0000000100000000001110111000010000",
			5387 => "0000001110000000001000101000001000",
			5388 => "0000001101000000001110010000000100",
			5389 => "11111111111110100101010010010001",
			5390 => "00000000110001110101010010010001",
			5391 => "0000000100000000001000011100000100",
			5392 => "00000000000000000101010010010001",
			5393 => "11111101111000010101010010010001",
			5394 => "00000000111010100101010010010001",
			5395 => "0000001000000000000110001000011100",
			5396 => "0000001101000000001010000100010100",
			5397 => "0000000101000000000101110000000100",
			5398 => "11111111011001010101010010010001",
			5399 => "0000001100000000000100000100001000",
			5400 => "0000001110000000001000001000000100",
			5401 => "00000001100111000101010010010001",
			5402 => "00000000000000000101010010010001",
			5403 => "0000001101000000000110111100000100",
			5404 => "00000001010110010101010010010001",
			5405 => "00000000000000000101010010010001",
			5406 => "0000001000000000000001010100000100",
			5407 => "11111110100101110101010010010001",
			5408 => "00000001100010010101010010010001",
			5409 => "0000000010000000000101010100000100",
			5410 => "00000000000000000101010010010001",
			5411 => "11111110111000010101010010010001",
			5412 => "0000001100000000001000000000001100",
			5413 => "0000000010000000000110111000000100",
			5414 => "11111110011010100101010101001101",
			5415 => "0000000010000000000110111000000100",
			5416 => "00000000100100010101010101001101",
			5417 => "11111110110000010101010101001101",
			5418 => "0000000001000000001101011001000000",
			5419 => "0000000011000000001110100100100100",
			5420 => "0000001001000000001001111100001100",
			5421 => "0000001100000000001000000000001000",
			5422 => "0000000001000000000101011100000100",
			5423 => "00000000000000000101010101001101",
			5424 => "00000000010100000101010101001101",
			5425 => "11111110110011000101010101001101",
			5426 => "0000000110000000000100111100001000",
			5427 => "0000001111000000001000101000000100",
			5428 => "00000000000000000101010101001101",
			5429 => "00000001100011110101010101001101",
			5430 => "0000000100000000001101001000001000",
			5431 => "0000000001000000001100011000000100",
			5432 => "11111110101101010101010101001101",
			5433 => "00000000011101100101010101001101",
			5434 => "0000000110000000001001111100000100",
			5435 => "00000001010101000101010101001101",
			5436 => "00000000000000000101010101001101",
			5437 => "0000000111000000000110110100010000",
			5438 => "0000001001000000000010101100001000",
			5439 => "0000000110000000000101010000000100",
			5440 => "00000000000111100101010101001101",
			5441 => "00000000000000000101010101001101",
			5442 => "0000001001000000000011101000000100",
			5443 => "11111110101101010101010101001101",
			5444 => "11111100110011010101010101001101",
			5445 => "0000001010000000000110011000000100",
			5446 => "00000001010011100101010101001101",
			5447 => "0000001101000000001100010000000100",
			5448 => "00000000000000000101010101001101",
			5449 => "11111110110000000101010101001101",
			5450 => "0000001010000000001000010100001000",
			5451 => "0000001001000000000011101000000100",
			5452 => "00000001001110000101010101001101",
			5453 => "11111110101101000101010101001101",
			5454 => "0000000110000000000100101100001000",
			5455 => "0000001101000000001110110100000100",
			5456 => "00000000000000000101010101001101",
			5457 => "00000001100011110101010101001101",
			5458 => "00000000001011110101010101001101",
			5459 => "0000001100000000001011000000000100",
			5460 => "11111110110011010101010111110001",
			5461 => "0000000011000000000110001100110100",
			5462 => "0000000100000000001100001100011100",
			5463 => "0000000110000000001000010000001100",
			5464 => "0000001001000000001010100100000100",
			5465 => "00000000000000000101010111110001",
			5466 => "0000000111000000000111010000000100",
			5467 => "00000000000000000101010111110001",
			5468 => "00000000101011110101010111110001",
			5469 => "0000001100000000001010001100001100",
			5470 => "0000001111000000001000110100000100",
			5471 => "00000000000000000101010111110001",
			5472 => "0000001000000000000001010100000100",
			5473 => "11111111000111100101010111110001",
			5474 => "00000000000000000101010111110001",
			5475 => "00000000000000000101010111110001",
			5476 => "0000001001000000000100101100001000",
			5477 => "0000001111000000001111101000000100",
			5478 => "00000000000000000101010111110001",
			5479 => "11111111110011110101010111110001",
			5480 => "0000000110000000001001111100001100",
			5481 => "0000001100000000000001011000001000",
			5482 => "0000001100000000001001110100000100",
			5483 => "00000000000000000101010111110001",
			5484 => "00000001000010000101010111110001",
			5485 => "00000000000000000101010111110001",
			5486 => "00000000000000000101010111110001",
			5487 => "0000001100000000000111010000010000",
			5488 => "0000001010000000001001000100000100",
			5489 => "00000000000000000101010111110001",
			5490 => "0000001111000000000110001100000100",
			5491 => "00000000000000000101010111110001",
			5492 => "0000001110000000001000011100000100",
			5493 => "00000000000000000101010111110001",
			5494 => "11111111010001100101010111110001",
			5495 => "0000000110000000000100101100001000",
			5496 => "0000000001000000001100011000000100",
			5497 => "00000000000000000101010111110001",
			5498 => "00000000101111100101010111110001",
			5499 => "11111111110100110101010111110001",
			5500 => "0000001001000000001010100100100000",
			5501 => "0000000010000000001101101100000100",
			5502 => "11111110011000110101011010110101",
			5503 => "0000001110000000001111101000011000",
			5504 => "0000001100000000000100011000000100",
			5505 => "11111110100000010101011010110101",
			5506 => "0000000100000000001110111000001000",
			5507 => "0000000001000000000100110100000100",
			5508 => "11111110100101100101011010110101",
			5509 => "00000000000000000101011010110101",
			5510 => "0000001100000000001000000000000100",
			5511 => "00000010111001100101011010110101",
			5512 => "0000001001000000000111101100000100",
			5513 => "11111110011100110101011010110101",
			5514 => "00000001000011100101011010110101",
			5515 => "11111110011010000101011010110101",
			5516 => "0000001011000000000001001000011100",
			5517 => "0000000100000000000011110000010000",
			5518 => "0000000110000000000100111100001000",
			5519 => "0000000101000000000101110000000100",
			5520 => "11111110110000010101011010110101",
			5521 => "00000001100001100101011010110101",
			5522 => "0000000001000000001010011000000100",
			5523 => "11111110000010110101011010110101",
			5524 => "11111111101000110101011010110101",
			5525 => "0000001110000000000110111000000100",
			5526 => "00000010111101110101011010110101",
			5527 => "0000000101000000001110010000000100",
			5528 => "11111110101000100101011010110101",
			5529 => "00000000100110110101011010110101",
			5530 => "0000001100000000001011011100100100",
			5531 => "0000000110000000001001111100011000",
			5532 => "0000001101000000001010000100010000",
			5533 => "0000001100000000000100000100001000",
			5534 => "0000000101000000001110110100000100",
			5535 => "00000001101010110101011010110101",
			5536 => "00000001000001100101011010110101",
			5537 => "0000000101000000000010000000000100",
			5538 => "00000000000000000101011010110101",
			5539 => "00000001100110000101011010110101",
			5540 => "0000000010000000000101000000000100",
			5541 => "11111110111010110101011010110101",
			5542 => "00000001100100100101011010110101",
			5543 => "0000000001000000001001100100000100",
			5544 => "11111110111100010101011010110101",
			5545 => "0000001100000000001111011100000100",
			5546 => "11111111111011110101011010110101",
			5547 => "00000001100100010101011010110101",
			5548 => "11111111001110110101011010110101",
			5549 => "0000001001000000001010100100101000",
			5550 => "0000000010000000001101101100000100",
			5551 => "11111110011000100101011101110001",
			5552 => "0000000110000000000101010000100000",
			5553 => "0000000100000000001110111000001100",
			5554 => "0000001100000000001000011000000100",
			5555 => "11111110011000110101011101110001",
			5556 => "0000000111000000000001011000000100",
			5557 => "00000000101000110101011101110001",
			5558 => "11111111000000110101011101110001",
			5559 => "0000001001000000001011001100000100",
			5560 => "11111110100111000101011101110001",
			5561 => "0000000010000000001100001100001000",
			5562 => "0000000111000000001011000000000100",
			5563 => "11111111100110110101011101110001",
			5564 => "00000011000000110101011101110001",
			5565 => "0000001001000000000100101100000100",
			5566 => "11111110100001110101011101110001",
			5567 => "00000001110010000101011101110001",
			5568 => "11111110011001010101011101110001",
			5569 => "0000001100000000001001110100001000",
			5570 => "0000000101000000000111111100000100",
			5571 => "11111110010001010101011101110001",
			5572 => "00000000101010010101011101110001",
			5573 => "0000001010000000000001010000011100",
			5574 => "0000001101000000001010000100010100",
			5575 => "0000001011000000000001001000001000",
			5576 => "0000001110000000000110111000000100",
			5577 => "00000001011110110101011101110001",
			5578 => "11111111111001110101011101110001",
			5579 => "0000001101000000000110111100000100",
			5580 => "00000001101011000101011101110001",
			5581 => "0000001011000000001110101100000100",
			5582 => "11111111001011000101011101110001",
			5583 => "00000001011011110101011101110001",
			5584 => "0000000000000000000111000000000100",
			5585 => "11111110011101010101011101110001",
			5586 => "00000001100101100101011101110001",
			5587 => "0000000100000000000100001100001000",
			5588 => "0000001001000000000111110100000100",
			5589 => "11111101101011110101011101110001",
			5590 => "00000001001011000101011101110001",
			5591 => "0000000110000000000100101100001000",
			5592 => "0000001110000000000010111000000100",
			5593 => "00000001111010110101011101110001",
			5594 => "00000000111100110101011101110001",
			5595 => "11111110110111000101011101110001",
			5596 => "0000000010000000001101101100001000",
			5597 => "0000000011000000000001011100000100",
			5598 => "11111110011011000101100000011101",
			5599 => "00000000000000000101100000011101",
			5600 => "0000001111000000001000000100100000",
			5601 => "0000000110000000000101010000010100",
			5602 => "0000001100000000001010111000000100",
			5603 => "11111111110101100101100000011101",
			5604 => "0000001001000000001011001100000100",
			5605 => "00000000000000000101100000011101",
			5606 => "0000000100000000000110111000000100",
			5607 => "00000000000000000101100000011101",
			5608 => "0000000110000000001111000000000100",
			5609 => "00000000000000000101100000011101",
			5610 => "00000001010110110101100000011101",
			5611 => "0000001111000000001011110000001000",
			5612 => "0000000001000000000001111000000100",
			5613 => "00000000000000000101100000011101",
			5614 => "00000000011010000101100000011101",
			5615 => "11111111010100100101100000011101",
			5616 => "0000000001000000001101011000101000",
			5617 => "0000001011000000000110100000011100",
			5618 => "0000001110000000001000011100010000",
			5619 => "0000001001000000000010101100001000",
			5620 => "0000000010000000001000110100000100",
			5621 => "11111110101101010101100000011101",
			5622 => "00000000000111110101100000011101",
			5623 => "0000000101000000000101110000000100",
			5624 => "00000000000000000101100000011101",
			5625 => "00000001011000000101100000011101",
			5626 => "0000001101000000000110111100001000",
			5627 => "0000001100000000000100000100000100",
			5628 => "11111110011010010101100000011101",
			5629 => "00000000000000000101100000011101",
			5630 => "00000000000000000101100000011101",
			5631 => "0000001001000000000011101000001000",
			5632 => "0000000100000000001101001000000100",
			5633 => "00000000110110110101100000011101",
			5634 => "11111110111010010101100000011101",
			5635 => "11111101100101110101100000011101",
			5636 => "0000001000000000000111000100000100",
			5637 => "00000001011101100101100000011101",
			5638 => "00000000000000000101100000011101",
			5639 => "0000001001000000001010100100100100",
			5640 => "0000000110000000000100111100000100",
			5641 => "11111110011001000101100100010001",
			5642 => "0000000110000000001000010000001100",
			5643 => "0000000100000000001110111000000100",
			5644 => "11111110110000010101100100010001",
			5645 => "0000001001000000001011001100000100",
			5646 => "11111111010111100101100100010001",
			5647 => "00000010001001000101100100010001",
			5648 => "0000001001000000000100101100000100",
			5649 => "11111110011000100101100100010001",
			5650 => "0000000100000000000011101100001100",
			5651 => "0000001001000000000111101100001000",
			5652 => "0000001001000000000111101100000100",
			5653 => "11111111110111110101100100010001",
			5654 => "00000000000000000101100100010001",
			5655 => "11111110011110110101100100010001",
			5656 => "00000001000100110101100100010001",
			5657 => "0000001011000000000000110100101000",
			5658 => "0000001110000000000110111000010100",
			5659 => "0000000100000000001000001000010000",
			5660 => "0000000101000000000111111100001000",
			5661 => "0000001000000000000101000100000100",
			5662 => "00000000001010110101100100010001",
			5663 => "11111110010100100101100100010001",
			5664 => "0000000110000000001000010000000100",
			5665 => "00000001011011000101100100010001",
			5666 => "00000000000000000101100100010001",
			5667 => "00000010100001000101100100010001",
			5668 => "0000001100000000001000011000010000",
			5669 => "0000000100000000000110001100000100",
			5670 => "11111100011110100101100100010001",
			5671 => "0000001010000000000110011000000100",
			5672 => "00000000011001110101100100010001",
			5673 => "0000000000000000000011111100000100",
			5674 => "11111110010010110101100100010001",
			5675 => "00000000000000000101100100010001",
			5676 => "00000001011111000101100100010001",
			5677 => "0000001101000000000110111100010000",
			5678 => "0000001100000000000001011000001000",
			5679 => "0000001110000000000011110000000100",
			5680 => "00000001100111100101100100010001",
			5681 => "00000000000000000101100100010001",
			5682 => "0000001011000000000110100000000100",
			5683 => "00000000111001100101100100010001",
			5684 => "11111111100100110101100100010001",
			5685 => "0000000010000000001000110100010000",
			5686 => "0000000011000000000101000000001000",
			5687 => "0000000100000000001100001100000100",
			5688 => "00000001100000110101100100010001",
			5689 => "00000000000000000101100100010001",
			5690 => "0000001010000000001000010100000100",
			5691 => "11111011111010000101100100010001",
			5692 => "00000001001001000101100100010001",
			5693 => "0000001000000000001111001000001000",
			5694 => "0000001110000000001000000100000100",
			5695 => "00000000000000000101100100010001",
			5696 => "00000001101000110101100100010001",
			5697 => "0000000100000000000011011000000100",
			5698 => "11111110100110010101100100010001",
			5699 => "00000000101000110101100100010001",
			5700 => "0000001100000000001011000000000100",
			5701 => "11111110011111110101100110111101",
			5702 => "0000001011000000000110100000111000",
			5703 => "0000001001000000000010101100100100",
			5704 => "0000001110000000000110111000010100",
			5705 => "0000001001000000000101010000000100",
			5706 => "11111111100011010101100110111101",
			5707 => "0000000100000000000010110000001000",
			5708 => "0000000111000000000111010000000100",
			5709 => "11111111010000100101100110111101",
			5710 => "00000000011100100101100110111101",
			5711 => "0000000110000000000101010000000100",
			5712 => "00000001010001100101100110111101",
			5713 => "00000000000000000101100110111101",
			5714 => "0000000110000000001000010000000100",
			5715 => "00000000000000000101100110111101",
			5716 => "0000000001000000001010011000001000",
			5717 => "0000000101000000001110110100000100",
			5718 => "11111110101111110101100110111101",
			5719 => "00000000000000000101100110111101",
			5720 => "00000000000000000101100110111101",
			5721 => "0000001100000000000001101000001100",
			5722 => "0000001100000000001001110100000100",
			5723 => "00000000001001010101100110111101",
			5724 => "0000000111000000000001011000000100",
			5725 => "11111111010110000101100110111101",
			5726 => "00000000000000000101100110111101",
			5727 => "0000001001000000001000010100000100",
			5728 => "00000001010101000101100110111101",
			5729 => "00000000000000000101100110111101",
			5730 => "0000000001000000001101011000010000",
			5731 => "0000001001000000000011101000001100",
			5732 => "0000000110000000000101010000001000",
			5733 => "0000000001000000001100011000000100",
			5734 => "00000000000000000101100110111101",
			5735 => "00000000100011010101100110111101",
			5736 => "11111111010001010101100110111101",
			5737 => "11111110101010010101100110111101",
			5738 => "0000001000000000000111000100001000",
			5739 => "0000001011000000000110100000000100",
			5740 => "00000000000000000101100110111101",
			5741 => "00000000110111110101100110111101",
			5742 => "11111111111111000101100110111101",
			5743 => "0000001001000000000111101100001000",
			5744 => "0000000100000000000000100000000100",
			5745 => "11111110100110110101101001101001",
			5746 => "00000000000000000101101001101001",
			5747 => "0000000110000000000100111100001100",
			5748 => "0000000111000000000111010000001000",
			5749 => "0000000100000000000110001100000100",
			5750 => "11111111110100010101101001101001",
			5751 => "00000000000000000101101001101001",
			5752 => "00000000111011010101101001101001",
			5753 => "0000000000000000000111000000011000",
			5754 => "0000001111000000001000011100001100",
			5755 => "0000001011000000000000110100001000",
			5756 => "0000000111000000000000011100000100",
			5757 => "00000000000000000101101001101001",
			5758 => "11111111010110010101101001101001",
			5759 => "00000000101000110101101001101001",
			5760 => "0000001001000000000011101000000100",
			5761 => "00000000000000000101101001101001",
			5762 => "0000001101000000000110111100000100",
			5763 => "00000000000000000101101001101001",
			5764 => "11111110101100010101101001101001",
			5765 => "0000000110000000000101010000010000",
			5766 => "0000000010000000001000000100000100",
			5767 => "00000000000000000101101001101001",
			5768 => "0000000111000000001111011100000100",
			5769 => "00000000000000000101101001101001",
			5770 => "0000000111000000000111110000000100",
			5771 => "00000001000101000101101001101001",
			5772 => "00000000000000000101101001101001",
			5773 => "0000000100000000000100001100001100",
			5774 => "0000001001000000001000100100001000",
			5775 => "0000001010000000000110011000000100",
			5776 => "00000000000000000101101001101001",
			5777 => "11111111000101000101101001101001",
			5778 => "00000000000000000101101001101001",
			5779 => "0000000000000000000011010000001000",
			5780 => "0000001001000000001010100100000100",
			5781 => "00000000000000000101101001101001",
			5782 => "00000000100110110101101001101001",
			5783 => "0000000100000000001011001000000100",
			5784 => "11111111001111010101101001101001",
			5785 => "00000000000100100101101001101001",
			5786 => "0000001100000000001011000000000100",
			5787 => "11111110011110100101101100011101",
			5788 => "0000001011000000000110100000111000",
			5789 => "0000000010000000000010110000101000",
			5790 => "0000000100000000001110100100010100",
			5791 => "0000000111000000000001011000001100",
			5792 => "0000000110000000001111000000000100",
			5793 => "00000000000000000101101100011101",
			5794 => "0000001011000000000000110100000100",
			5795 => "11111110100011100101101100011101",
			5796 => "00000000000000000101101100011101",
			5797 => "0000000001000000000100110100000100",
			5798 => "00000000000000000101101100011101",
			5799 => "00000001000010010101101100011101",
			5800 => "0000001100000000000100000100001100",
			5801 => "0000001001000000000101010000000100",
			5802 => "11111111111111000101101100011101",
			5803 => "0000000111000000001000011000000100",
			5804 => "00000000000000000101101100011101",
			5805 => "00000001000110110101101100011101",
			5806 => "0000000101000000000010000000000100",
			5807 => "11111111011101100101101100011101",
			5808 => "00000000000000000101101100011101",
			5809 => "0000001001000000000111110100001000",
			5810 => "0000001100000000000100000100000100",
			5811 => "11111110111101110101101100011101",
			5812 => "00000000000000000101101100011101",
			5813 => "0000001010000000001010110000000100",
			5814 => "00000000000000000101101100011101",
			5815 => "00000000000000000101101100011101",
			5816 => "0000000001000000001101011000010100",
			5817 => "0000000110000000001000010000000100",
			5818 => "00000000000000000101101100011101",
			5819 => "0000001100000000001111011100000100",
			5820 => "00000000000000000101101100011101",
			5821 => "0000001110000000001110100100001000",
			5822 => "0000000101000000000110010000000100",
			5823 => "00000000000000000101101100011101",
			5824 => "11111110100000010101101100011101",
			5825 => "00000000000000000101101100011101",
			5826 => "0000001010000000000110011100001000",
			5827 => "0000001011000000000110100000000100",
			5828 => "00000000000000000101101100011101",
			5829 => "00000000111010100101101100011101",
			5830 => "11111111111011000101101100011101",
			5831 => "0000000010000000001101101100001000",
			5832 => "0000001011000000001010010100000100",
			5833 => "11111110011010110101101111101001",
			5834 => "00000000000000000101101111101001",
			5835 => "0000001001000000000010101100111100",
			5836 => "0000001110000000000110111000011100",
			5837 => "0000001001000000001010100100010100",
			5838 => "0000000100000000000100001100001000",
			5839 => "0000000110000000000100111100000100",
			5840 => "00000000000000000101101111101001",
			5841 => "11111110100111010101101111101001",
			5842 => "0000001010000000000101000100001000",
			5843 => "0000001100000000000001101000000100",
			5844 => "00000001010110100101101111101001",
			5845 => "00000000000000000101101111101001",
			5846 => "11111111100000110101101111101001",
			5847 => "0000001101000000001100010100000100",
			5848 => "00000000000000000101101111101001",
			5849 => "00000001010010100101101111101001",
			5850 => "0000001100000000001000011000010000",
			5851 => "0000000100000000000000010100001100",
			5852 => "0000001011000000001110101100001000",
			5853 => "0000001111000000001000110100000100",
			5854 => "00000000000000000101101111101001",
			5855 => "11111110000010110101101111101001",
			5856 => "00000000000000000101101111101001",
			5857 => "00000000000000000101101111101001",
			5858 => "0000001100000000000100000100001100",
			5859 => "0000001010000000001010110000001000",
			5860 => "0000001001000000001010100100000100",
			5861 => "00000000000000000101101111101001",
			5862 => "00000001001111000101101111101001",
			5863 => "00000000000000000101101111101001",
			5864 => "11111110110111010101101111101001",
			5865 => "0000001100000000000110100100001100",
			5866 => "0000001100000000001001110100001000",
			5867 => "0000001000000000001001101000000100",
			5868 => "00000000000000000101101111101001",
			5869 => "00000000011000010101101111101001",
			5870 => "11111110110100000101101111101001",
			5871 => "0000001101000000000110111100000100",
			5872 => "00000001100000100101101111101001",
			5873 => "0000001100000000000111010000001100",
			5874 => "0000000011000000000101000000000100",
			5875 => "00000000100010100101101111101001",
			5876 => "0000001000000000000001010100000100",
			5877 => "11111110100000100101101111101001",
			5878 => "00000000000000000101101111101001",
			5879 => "0000001100000000001011011100000100",
			5880 => "00000001011001100101101111101001",
			5881 => "00000000000000000101101111101001",
			5882 => "0000000001000000000100110100011100",
			5883 => "0000000010000000001110000000000100",
			5884 => "11111110011001100101110011000101",
			5885 => "0000001111000000001110100100010100",
			5886 => "0000001100000000001011000000000100",
			5887 => "11111110111101110101110011000101",
			5888 => "0000001100000000001000011000001000",
			5889 => "0000000100000000001110111000000100",
			5890 => "00000000000000000101110011000101",
			5891 => "00000001100111010101110011000101",
			5892 => "0000001011000000000001001000000100",
			5893 => "00000000000000000101110011000101",
			5894 => "11111110111110100101110011000101",
			5895 => "11111110100001110101110011000101",
			5896 => "0000001100000000001000011000101000",
			5897 => "0000001110000000000110001100100100",
			5898 => "0000000100000000000011110000010000",
			5899 => "0000001011000000000001001000001100",
			5900 => "0000000110000000000100111100001000",
			5901 => "0000001110000000001111100100000100",
			5902 => "11111111010001000101110011000101",
			5903 => "00000000001110010101110011000101",
			5904 => "11111110001110100101110011000101",
			5905 => "00000001001111010101110011000101",
			5906 => "0000000110000000000101010000001000",
			5907 => "0000001011000000000100010000000100",
			5908 => "00000000000000000101110011000101",
			5909 => "00000010000000000101110011000101",
			5910 => "0000000100000000001001001100001000",
			5911 => "0000001111000000001000110100000100",
			5912 => "00000000000000000101110011000101",
			5913 => "11111111000111110101110011000101",
			5914 => "00000000100001110101110011000101",
			5915 => "11111110000100000101110011000101",
			5916 => "0000001011000000000110100000010100",
			5917 => "0000000110000000001001111100010000",
			5918 => "0000001011000000000000110100001100",
			5919 => "0000001110000000001000011100001000",
			5920 => "0000001100000000001000011000000100",
			5921 => "00000000000000000101110011000101",
			5922 => "00000001100010010101110011000101",
			5923 => "11111101001001100101110011000101",
			5924 => "00000001100101110101110011000101",
			5925 => "11111111101010000101110011000101",
			5926 => "0000000111000000000110110100000100",
			5927 => "11111010101111010101110011000101",
			5928 => "0000000000000000001010101100001000",
			5929 => "0000001111000000001000011100000100",
			5930 => "00000000111100100101110011000101",
			5931 => "11111110001100010101110011000101",
			5932 => "0000001010000000001010110000000100",
			5933 => "00000001011111010101110011000101",
			5934 => "0000000100000000000111011100000100",
			5935 => "11111110111001100101110011000101",
			5936 => "00000000010001010101110011000101",
			5937 => "0000000010000000001101101100001000",
			5938 => "0000001011000000001010010100000100",
			5939 => "11111110011010000101110110011001",
			5940 => "00000000000000000101110110011001",
			5941 => "0000000001000000001100011000111000",
			5942 => "0000000110000000000101010000101100",
			5943 => "0000000100000000001000001000010100",
			5944 => "0000001100000000001000011000001100",
			5945 => "0000000110000000000100111100000100",
			5946 => "00000000000000000101110110011001",
			5947 => "0000001000000000000101000100000100",
			5948 => "00000000000000000101110110011001",
			5949 => "11111110011111100101110110011001",
			5950 => "0000000001000000000100110100000100",
			5951 => "00000000000000000101110110011001",
			5952 => "00000000111100110101110110011001",
			5953 => "0000000001000000000111101000001100",
			5954 => "0000001111000000000010010100001000",
			5955 => "0000001001000000001011001100000100",
			5956 => "11111111101101000101110110011001",
			5957 => "00000001101011100101110110011001",
			5958 => "11111110101100110101110110011001",
			5959 => "0000001011000000000100010000000100",
			5960 => "00000000000000000101110110011001",
			5961 => "0000001101000000000010000100000100",
			5962 => "00000001101111000101110110011001",
			5963 => "00000000000000000101110110011001",
			5964 => "0000001011000000000000110100001000",
			5965 => "0000001011000000001011110100000100",
			5966 => "11111110111100110101110110011001",
			5967 => "00000000000000000101110110011001",
			5968 => "11111110011110110101110110011001",
			5969 => "0000001100000000000110100100010000",
			5970 => "0000001001000000000010101100001000",
			5971 => "0000001001000000000010101100000100",
			5972 => "00000000000000000101110110011001",
			5973 => "00000000001000110101110110011001",
			5974 => "0000000101000000000011001000000100",
			5975 => "11111110011011010101110110011001",
			5976 => "00000000000000000101110110011001",
			5977 => "0000001101000000000110111100001000",
			5978 => "0000001011000000000001001000000100",
			5979 => "00000000000000000101110110011001",
			5980 => "00000001100101000101110110011001",
			5981 => "0000001011000000001110101100000100",
			5982 => "11111110000111100101110110011001",
			5983 => "0000000001000000001101011000001000",
			5984 => "0000000001000000001101011000000100",
			5985 => "00000000110001110101110110011001",
			5986 => "11111110100111100101110110011001",
			5987 => "0000001000000000000111000100000100",
			5988 => "00000001011110110101110110011001",
			5989 => "11111111010000100101110110011001",
			5990 => "0000001001000000000100111100000100",
			5991 => "11111110111010110101111001001101",
			5992 => "0000001110000000000110111000100100",
			5993 => "0000000100000000001001000000100000",
			5994 => "0000001001000000001010100000001000",
			5995 => "0000001111000000001000011100000100",
			5996 => "11111111100001100101111001001101",
			5997 => "00000000000000000101111001001101",
			5998 => "0000001111000000000010010100001100",
			5999 => "0000000110000000001111000000000100",
			6000 => "00000000000000000101111001001101",
			6001 => "0000001100000000000001101000000100",
			6002 => "11111111011111100101111001001101",
			6003 => "00000000000000000101111001001101",
			6004 => "0000000110000000000101010000001000",
			6005 => "0000001101000000001010001000000100",
			6006 => "00000000000000000101111001001101",
			6007 => "00000000101101010101111001001101",
			6008 => "00000000000000000101111001001101",
			6009 => "00000000110010010101111001001101",
			6010 => "0000000001000000001101011000101000",
			6011 => "0000001011000000001110101100010000",
			6012 => "0000001111000000001000110100000100",
			6013 => "00000000000000000101111001001101",
			6014 => "0000001001000000001010100100000100",
			6015 => "00000000000000000101111001001101",
			6016 => "0000000110000000000100111100000100",
			6017 => "00000000000000000101111001001101",
			6018 => "11111110110101110101111001001101",
			6019 => "0000001001000000000011101000001100",
			6020 => "0000000100000000001101001000001000",
			6021 => "0000000001000000000100110100000100",
			6022 => "00000000000000000101111001001101",
			6023 => "00000000101000000101111001001101",
			6024 => "00000000000000000101111001001101",
			6025 => "0000001011000000001101000100001000",
			6026 => "0000001111000000001000011100000100",
			6027 => "00000000000000000101111001001101",
			6028 => "11111111011010100101111001001101",
			6029 => "00000000000000000101111001001101",
			6030 => "0000000110000000000100101100001000",
			6031 => "0000000011000000001000000100000100",
			6032 => "00000000000000000101111001001101",
			6033 => "00000000110001110101111001001101",
			6034 => "11111111110100010101111001001101",
			6035 => "0000001100000000001011000000000100",
			6036 => "11111110011001110101111011100011",
			6037 => "0000000001000000001011111100000100",
			6038 => "11111110100100110101111011100011",
			6039 => "0000001011000000000110100000101000",
			6040 => "0000001011000000000000110100011000",
			6041 => "0000001110000000001000011100010000",
			6042 => "0000000010000000001110000000001000",
			6043 => "0000001011000000000000110100000100",
			6044 => "11111111001000010101111011100011",
			6045 => "00000001011000110101111011100011",
			6046 => "0000000110000000001001111100000100",
			6047 => "00000001011010110101111011100011",
			6048 => "11111110111111110101111011100011",
			6049 => "0000000001000000001101011000000100",
			6050 => "11111101100001000101111011100011",
			6051 => "00000001001111010101111011100011",
			6052 => "0000000110000000001001111100001100",
			6053 => "0000000001000000000100110100001000",
			6054 => "0000001111000000000101000000000100",
			6055 => "00000000000000000101111011100011",
			6056 => "11111111011010000101111011100011",
			6057 => "00000001100101110101111011100011",
			6058 => "11111110111100010101111011100011",
			6059 => "0000000111000000000110110100000100",
			6060 => "11111100010101000101111011100011",
			6061 => "0000000000000000001010101100001000",
			6062 => "0000001111000000001000011100000100",
			6063 => "00000000110110000101111011100011",
			6064 => "11111110011110110101111011100011",
			6065 => "0000001010000000001010110000001000",
			6066 => "0000000001000000001100011000000100",
			6067 => "00000000000000000101111011100011",
			6068 => "00000001011100110101111011100011",
			6069 => "0000000001000000001001100100000100",
			6070 => "11111110101100000101111011100011",
			6071 => "00000000010100100101111011100011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1980, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(4056, initial_addr_3'length));
	end generate gen_rom_8;

	gen_rom_9: if SELECT_ROM = 9 generate
		bank <= (
			0 => "0000001101000000001110110000010100",
			1 => "0000000100000000000000101100000100",
			2 => "11111110011111000000000010110101",
			3 => "0000001000000000001101010000001000",
			4 => "0000001010000000000001110000000100",
			5 => "00000000000000000000000010110101",
			6 => "00000000010011010000000010110101",
			7 => "0000000010000000001111010100000100",
			8 => "11111111010000110000000010110101",
			9 => "00000000000000000000000010110101",
			10 => "0000001100000000000100000000010000",
			11 => "0000001111000000000011001000001000",
			12 => "0000000110000000001011001100000100",
			13 => "11111111100100000000000010110101",
			14 => "00000001100100010000000010110101",
			15 => "0000000001000000000111100100000100",
			16 => "11111110101101100000000010110101",
			17 => "00000000101010110000000010110101",
			18 => "0000001101000000001011000000011000",
			19 => "0000000100000000000011011000010000",
			20 => "0000000111000000001000111100000100",
			21 => "00000000000000000000000010110101",
			22 => "0000001000000000000110001000000100",
			23 => "00000000000000000000000010110101",
			24 => "0000001111000000001101000100000100",
			25 => "00000000000000000000000010110101",
			26 => "11111110011110000000000010110101",
			27 => "0000000110000000001001100100000100",
			28 => "00000000000000000000000010110101",
			29 => "00000000110111010000000010110101",
			30 => "0000000111000000001000111000000100",
			31 => "00000001100011010000000010110101",
			32 => "0000001011000000000110000100001100",
			33 => "0000000110000000001001100100001000",
			34 => "0000000010000000001100010000000100",
			35 => "00000001000101100000000010110101",
			36 => "11111110110100010000000010110101",
			37 => "00000001100011010000000010110101",
			38 => "0000000001000000001011101000001000",
			39 => "0000001100000000000011011100000100",
			40 => "11111111111001010000000010110101",
			41 => "11111110101001110000000010110101",
			42 => "0000001011000000001001110100000100",
			43 => "00000001011011110000000010110101",
			44 => "00000000000111000000000010110101",
			45 => "0000000101000000001010111100010100",
			46 => "0000000010000000001100000000001000",
			47 => "0000001101000000001010111000000100",
			48 => "11111110011101110000000101101001",
			49 => "00000000000000000000000101101001",
			50 => "0000001101000000000001111100000100",
			51 => "11111111011111100000000101101001",
			52 => "0000000000000000001100001000000100",
			53 => "11111111101111000000000101101001",
			54 => "00000000001111010000000101101001",
			55 => "0000001101000000001101101101000100",
			56 => "0000001100000000000000101000010100",
			57 => "0000000111000000001000111000001100",
			58 => "0000001011000000001101100000001000",
			59 => "0000000000000000000010011000000100",
			60 => "00000000000000000000000101101001",
			61 => "00000000000110000000000101101001",
			62 => "11111111010111100000000101101001",
			63 => "0000000110000000001011001100000100",
			64 => "00000000000000000000000101101001",
			65 => "00000001101101000000000101101001",
			66 => "0000000011000000000010000000100000",
			67 => "0000000000000000000010011000010000",
			68 => "0000000010000000001001100000001000",
			69 => "0000000011000000000111110000000100",
			70 => "11111111001011110000000101101001",
			71 => "00000000101100010000000101101001",
			72 => "0000001100000000000100000000000100",
			73 => "00000000000010110000000101101001",
			74 => "11111110010110100000000101101001",
			75 => "0000000010000000001100000000001000",
			76 => "0000000011000000001111011100000100",
			77 => "11111111110010100000000101101001",
			78 => "00000000111000100000000101101001",
			79 => "0000000110000000001111000000000100",
			80 => "11111110110011000000000101101001",
			81 => "00000000001111110000000101101001",
			82 => "0000000111000000000001111100000100",
			83 => "00000001101110100000000101101001",
			84 => "0000000011000000000010000100000100",
			85 => "11111110101100100000000101101001",
			86 => "0000000101000000000111100000000100",
			87 => "00000000100100010000000101101001",
			88 => "00000000000100010000000101101001",
			89 => "11111110011011100000000101101001",
			90 => "0000000001000000000110101001000000",
			91 => "0000000100000000000011011000101000",
			92 => "0000001100000000001000111000011100",
			93 => "0000000011000000000000011100001100",
			94 => "0000001100000000000100010100000100",
			95 => "00000000000000000000001010001101",
			96 => "0000000100000000000111011100000100",
			97 => "11111111010011000000001010001101",
			98 => "00000000000000000000001010001101",
			99 => "0000001111000000000111111100000100",
			100 => "00000000110001010000001010001101",
			101 => "0000000100000000000010111000000100",
			102 => "11111110111011010000001010001101",
			103 => "0000001111000000001110010000000100",
			104 => "00000000010011110000001010001101",
			105 => "00000000000000000000001010001101",
			106 => "0000001100000000000011011100001000",
			107 => "0000000111000000001000111000000100",
			108 => "00000000000000000000001010001101",
			109 => "11111110101000010000001010001101",
			110 => "00000000000000000000001010001101",
			111 => "0000001000000000001111000100001000",
			112 => "0000000110000000001011001100000100",
			113 => "00000000000000000000001010001101",
			114 => "00000001000001010000001010001101",
			115 => "0000000100000000000110110000000100",
			116 => "11111111011001010000001010001101",
			117 => "0000001111000000000100010000000100",
			118 => "00000000000000000000001010001101",
			119 => "0000000010000000001111100100000100",
			120 => "00000000001001010000001010001101",
			121 => "00000000000000000000001010001101",
			122 => "0000001110000000000101110100010100",
			123 => "0000000100000000000101010100001100",
			124 => "0000000011000000001011011100000100",
			125 => "00000000000000000000001010001101",
			126 => "0000000110000000001010011000000100",
			127 => "00000000000000000000001010001101",
			128 => "00000001010001110000001010001101",
			129 => "0000000110000000000100111100000100",
			130 => "11111111110110000000001010001101",
			131 => "00000000000000000000001010001101",
			132 => "0000001001000000001110010100001100",
			133 => "0000000110000000001000010000001000",
			134 => "0000000100000000000010010100000100",
			135 => "00000000000000000000001010001101",
			136 => "11111111001010100000001010001101",
			137 => "00000000000000000000001010001101",
			138 => "0000001001000000001101111100010100",
			139 => "0000001111000000000010000000001000",
			140 => "0000001011000000000000001100000100",
			141 => "00000000000000000000001010001101",
			142 => "11111111101010000000001010001101",
			143 => "0000001110000000000111111100001000",
			144 => "0000000100000000000110111000000100",
			145 => "00000000000000000000001010001101",
			146 => "00000001001100100000001010001101",
			147 => "00000000000000000000001010001101",
			148 => "0000001111000000001011110000010000",
			149 => "0000001000000000000001010100001000",
			150 => "0000000101000000000010011100000100",
			151 => "00000000000000000000001010001101",
			152 => "00000000100100010000001010001101",
			153 => "0000000110000000000101010000000100",
			154 => "11111111001011000000001010001101",
			155 => "00000000100101110000001010001101",
			156 => "0000000011000000001110000000001000",
			157 => "0000000000000000000111000000000100",
			158 => "00000000000000000000001010001101",
			159 => "00000000111000100000001010001101",
			160 => "0000000110000000000100101100000100",
			161 => "00000000000110010000001010001101",
			162 => "11111111011001110000001010001101",
			163 => "0000000001000000000110101001000100",
			164 => "0000001010000000000101000100100100",
			165 => "0000001100000000000000101000001000",
			166 => "0000001101000000001110110000000100",
			167 => "00000000000000000000001110110001",
			168 => "00000000000000000000001110110001",
			169 => "0000001101000000001000000000001000",
			170 => "0000000111000000000100000000000100",
			171 => "00000000000000000000001110110001",
			172 => "11111110111101000000001110110001",
			173 => "0000001110000000000101100100010000",
			174 => "0000001100000000001000111000001000",
			175 => "0000000111000000001001110000000100",
			176 => "00000000101001010000001110110001",
			177 => "00000000000000000000001110110001",
			178 => "0000000010000000001100000000000100",
			179 => "00000000000000000000001110110001",
			180 => "11111111010111000000001110110001",
			181 => "11111110111000000000001110110001",
			182 => "0000001000000000001111000100010000",
			183 => "0000000100000000001001000000000100",
			184 => "00000000000000000000001110110001",
			185 => "0000000011000000001101010100000100",
			186 => "00000000000000000000001110110001",
			187 => "0000001101000000000111001000000100",
			188 => "00000000000000000000001110110001",
			189 => "00000000111011010000001110110001",
			190 => "0000000100000000000110110000000100",
			191 => "11111111011101010000001110110001",
			192 => "0000001111000000000100010000000100",
			193 => "00000000000000000000001110110001",
			194 => "0000000010000000001111100100000100",
			195 => "00000000001000110000001110110001",
			196 => "00000000000000000000001110110001",
			197 => "0000001110000000000101110100010100",
			198 => "0000000100000000000101010100001100",
			199 => "0000000011000000001011011100000100",
			200 => "00000000000000000000001110110001",
			201 => "0000000000000000000001110000000100",
			202 => "00000000000000000000001110110001",
			203 => "00000001001110100000001110110001",
			204 => "0000001010000000000110011100000100",
			205 => "11111111111111000000001110110001",
			206 => "00000000000000000000001110110001",
			207 => "0000001001000000001011111100001000",
			208 => "0000001111000000000110010000000100",
			209 => "00000000000000000000001110110001",
			210 => "11111111000100100000001110110001",
			211 => "0000001011000000001101000100100000",
			212 => "0000000010000000001000110100010000",
			213 => "0000000010000000000011000000001000",
			214 => "0000001000000000000110001000000100",
			215 => "00000000000001010000001110110001",
			216 => "00000000111000010000001110110001",
			217 => "0000001001000000000111101100000100",
			218 => "11111111010000000000001110110001",
			219 => "00000000010010100000001110110001",
			220 => "0000001000000000000010101000001000",
			221 => "0000001100000000001001001000000100",
			222 => "00000001001001000000001110110001",
			223 => "00000000001011100000001110110001",
			224 => "0000000001000000000000111100000100",
			225 => "00000000000000000000001110110001",
			226 => "11111111110011000000001110110001",
			227 => "0000001001000000000111101100001000",
			228 => "0000000000000000000011010000000100",
			229 => "00000000000111100000001110110001",
			230 => "00000000000000000000001110110001",
			231 => "0000000000000000001010101100000100",
			232 => "00000000000000000000001110110001",
			233 => "0000001001000000001001000100000100",
			234 => "11111110111111110000001110110001",
			235 => "00000000000000000000001110110001",
			236 => "0000001101000000001110110000010100",
			237 => "0000000100000000000000101100000100",
			238 => "11111110011111110000010010011101",
			239 => "0000000000000000000011011100001000",
			240 => "0000001010000000000001010100000100",
			241 => "00000000000000000000010010011101",
			242 => "00000000010010000000010010011101",
			243 => "0000001010000000001111001000000100",
			244 => "11111111010111010000010010011101",
			245 => "00000000000000000000010010011101",
			246 => "0000000110000000000100101101010100",
			247 => "0000001111000000001000110100101000",
			248 => "0000001100000000000100000000010000",
			249 => "0000001111000000000011001000001000",
			250 => "0000000110000000001011001100000100",
			251 => "11111111100101110000010010011101",
			252 => "00000001100001010000010010011101",
			253 => "0000001011000000001100101100000100",
			254 => "11111110110000100000010010011101",
			255 => "00000000100111010000010010011101",
			256 => "0000001100000000000100000000001000",
			257 => "0000000001000000000111100100000100",
			258 => "11111110001100110000010010011101",
			259 => "00000000010000110000010010011101",
			260 => "0000000101000000000111100000001000",
			261 => "0000000100000000000110111000000100",
			262 => "00000000011111110000010010011101",
			263 => "11111111111111100000010010011101",
			264 => "0000001101000000001100010100000100",
			265 => "11111111001000010000010010011101",
			266 => "00000000001010100000010010011101",
			267 => "0000000100000000000100001100011000",
			268 => "0000000001000000001101011000001100",
			269 => "0000001000000000000001010100000100",
			270 => "00000000000000000000010010011101",
			271 => "0000000000000000001010101100000100",
			272 => "00000000000000000000010010011101",
			273 => "00000001001001000000010010011101",
			274 => "0000000000000000001010101100000100",
			275 => "00000000000000000000010010011101",
			276 => "0000000101000000000011001000000100",
			277 => "00000000000000000000010010011101",
			278 => "11111111010101100000010010011101",
			279 => "0000000101000000001110010000000100",
			280 => "11111110110001010000010010011101",
			281 => "0000001100000000001111011100001000",
			282 => "0000000011000000001110100100000100",
			283 => "00000000000000000000010010011101",
			284 => "00000001010100110000010010011101",
			285 => "0000001010000000001010110000000100",
			286 => "00000000000101000000010010011101",
			287 => "11111111011011010000010010011101",
			288 => "0000001110000000000011110000000100",
			289 => "00000000000000000000010010011101",
			290 => "0000001110000000001011100000000100",
			291 => "11111110001110000000010010011101",
			292 => "0000000110000000001010100000000100",
			293 => "00000000110000000000010010011101",
			294 => "11111111101000110000010010011101",
			295 => "0000001111000000001001010001000000",
			296 => "0000000011000000001001110100011100",
			297 => "0000000100000000000010010000001000",
			298 => "0000001101000000001000011000000100",
			299 => "11111111001010110000010110110001",
			300 => "00000000000000000000010110110001",
			301 => "0000001011000000001000111100000100",
			302 => "00000000000000000000010110110001",
			303 => "0000000010000000000010000100000100",
			304 => "00000000000000000000010110110001",
			305 => "0000000010000000001000100000001000",
			306 => "0000001011000000001100101100000100",
			307 => "00000000011100110000010110110001",
			308 => "00000000000000000000010110110001",
			309 => "00000000000000000000010110110001",
			310 => "0000000110000000001011001100011000",
			311 => "0000001100000000000100000000001000",
			312 => "0000001001000000001011101000000100",
			313 => "00000000000000000000010110110001",
			314 => "11111111011001110000010110110001",
			315 => "0000001100000000000100000000001000",
			316 => "0000001101000000000011100000000100",
			317 => "00000000000000000000010110110001",
			318 => "00000000101010000000010110110001",
			319 => "0000001001000000000001111000000100",
			320 => "11111111101011100000010110110001",
			321 => "00000000000000000000010110110001",
			322 => "0000000010000000000010000000000100",
			323 => "00000000000000000000010110110001",
			324 => "0000001101000000001001001000000100",
			325 => "00000001000110100000010110110001",
			326 => "00000000000000000000010110110001",
			327 => "0000000011000000000001011000000100",
			328 => "11111110111011010000010110110001",
			329 => "0000001000000000000001110100110000",
			330 => "0000000000000000000000111000100000",
			331 => "0000000001000000001001011000010000",
			332 => "0000001100000000001001110000001000",
			333 => "0000000110000000001001100100000100",
			334 => "11111111010010100000010110110001",
			335 => "00000000010101110000010110110001",
			336 => "0000000100000000001110111000000100",
			337 => "11111110101010010000010110110001",
			338 => "00000000000000000000010110110001",
			339 => "0000000001000000000101011100001000",
			340 => "0000000110000000001010011000000100",
			341 => "00000000000000000000010110110001",
			342 => "00000001000011100000010110110001",
			343 => "0000001111000000001110000000000100",
			344 => "11111111111010000000010110110001",
			345 => "00000000010000100000010110110001",
			346 => "0000000000000000000000110000001000",
			347 => "0000001100000000001100110000000100",
			348 => "00000001010011000000010110110001",
			349 => "00000000000000000000010110110001",
			350 => "0000001010000000001100011100000100",
			351 => "11111111101101110000010110110001",
			352 => "00000000000000000000010110110001",
			353 => "0000001010000000000101000100001000",
			354 => "0000001110000000000101100100000100",
			355 => "00000000000000000000010110110001",
			356 => "11111110110011100000010110110001",
			357 => "0000001000000000001111000100001100",
			358 => "0000001100000000000011011100000100",
			359 => "00000000111001010000010110110001",
			360 => "0000001001000000001010100100000100",
			361 => "11111111100110010000010110110001",
			362 => "00000000100000000000010110110001",
			363 => "11111111010110010000010110110001",
			364 => "0000000110000000001010011000100100",
			365 => "0000000001000000000101011100010000",
			366 => "0000001010000000001010100000001100",
			367 => "0000000000000000001100000100000100",
			368 => "11111110011100010000011011001101",
			369 => "0000001110000000001100110000000100",
			370 => "00000000000000000000011011001101",
			371 => "00000010001010010000011011001101",
			372 => "11111110011001000000011011001101",
			373 => "0000000110000000001010011000001100",
			374 => "0000001101000000000010011100001000",
			375 => "0000000111000000000110100100000100",
			376 => "11111110111111110000011011001101",
			377 => "00000001011111000000011011001101",
			378 => "00000011100110010000011011001101",
			379 => "0000001001000000000100101100000100",
			380 => "11111110100110000000011011001101",
			381 => "00000000010110010000011011001101",
			382 => "0000001010000000001001101001011100",
			383 => "0000000110000000001000010000111000",
			384 => "0000000100000000000011000000011000",
			385 => "0000000000000000001111001000001100",
			386 => "0000001010000000000011101000001000",
			387 => "0000000001000000001101111100000100",
			388 => "00000000101011110000011011001101",
			389 => "00000101111101110000011011001101",
			390 => "11111110011111100000011011001101",
			391 => "0000000010000000000000010000001000",
			392 => "0000001100000000000100011000000100",
			393 => "00000001011000110000011011001101",
			394 => "00000011100011000000011011001101",
			395 => "11111110110000010000011011001101",
			396 => "0000001100000000001000111100010000",
			397 => "0000001101000000001110110000001000",
			398 => "0000000100000000001100111100000100",
			399 => "11111110100110000000011011001101",
			400 => "00000001011011100000011011001101",
			401 => "0000000000000000000011010000000100",
			402 => "00000000100011000000011011001101",
			403 => "00000001011101110000011011001101",
			404 => "0000000011000000001011011100001000",
			405 => "0000000100000000000011010100000100",
			406 => "11111101111111010000011011001101",
			407 => "11111111110011100000011011001101",
			408 => "0000000111000000000101101100000100",
			409 => "00000001001001110000011011001101",
			410 => "11111111110011010000011011001101",
			411 => "0000000111000000001111011100010100",
			412 => "0000000100000000000111011100001100",
			413 => "0000000100000000000011110100001000",
			414 => "0000000001000000000101011100000100",
			415 => "00000000101011100000011011001101",
			416 => "00000001101011110000011011001101",
			417 => "00000010110111110000011011001101",
			418 => "0000000001000000001101011100000100",
			419 => "00000001000110100000011011001101",
			420 => "11111110011101010000011011001101",
			421 => "0000001010000000000110011000000100",
			422 => "11111110100000100000011011001101",
			423 => "0000000011000000001011110000000100",
			424 => "11111110001110110000011011001101",
			425 => "0000000110000000000101010000000100",
			426 => "00000001011011100000011011001101",
			427 => "00000000000000000000011011001101",
			428 => "0000001100000000000100000000000100",
			429 => "00000000101001100000011011001101",
			430 => "0000000000000000000110000100000100",
			431 => "11111100111101000000011011001101",
			432 => "0000000000000000001100101100000100",
			433 => "00000000011000110000011011001101",
			434 => "11111110011011100000011011001101",
			435 => "0000000011000000000111110001001000",
			436 => "0000001011000000001100101100111000",
			437 => "0000001110000000000010001000110000",
			438 => "0000001101000000001000000000100000",
			439 => "0000000111000000001000111000010000",
			440 => "0000000101000000001101010100001000",
			441 => "0000000010000000001100000000000100",
			442 => "11111111000001110000011111110001",
			443 => "00000000000000000000011111110001",
			444 => "0000000010000000000010000100000100",
			445 => "00000000101111010000011111110001",
			446 => "00000000000000000000011111110001",
			447 => "0000000100000000001110111000001000",
			448 => "0000001011000000001100101100000100",
			449 => "11111110101101100000011111110001",
			450 => "00000000000000000000011111110001",
			451 => "0000000000000000001010000000000100",
			452 => "00000000000111000000011111110001",
			453 => "11111111110011100000011111110001",
			454 => "0000000110000000001001100100001100",
			455 => "0000001001000000001001011000001000",
			456 => "0000000010000000000010000100000100",
			457 => "00000000111111100000011111110001",
			458 => "00000000000000000000011111110001",
			459 => "11111111001010110000011111110001",
			460 => "00000001011100010000011111110001",
			461 => "0000000011000000000101110100000100",
			462 => "11111110101010010000011111110001",
			463 => "00000000000000000000011111110001",
			464 => "0000000110000000001111000000001000",
			465 => "0000000010000000000001000000000100",
			466 => "00000000000000000000011111110001",
			467 => "11111110010110110000011111110001",
			468 => "0000001101000000000001101000000100",
			469 => "00000000010000000000011111110001",
			470 => "11111111101101010000011111110001",
			471 => "0000000101000000000100000100010100",
			472 => "0000000000000000001000101100000100",
			473 => "00000000000000000000011111110001",
			474 => "0000001001000000001011111100001100",
			475 => "0000001011000000001110001100000100",
			476 => "00000000100011010000011111110001",
			477 => "0000000100000000001010110100000100",
			478 => "11111111100001110000011111110001",
			479 => "00000000000000000000011111110001",
			480 => "00000001000010000000011111110001",
			481 => "0000001001000000001100011000001100",
			482 => "0000000011000000000010000000000100",
			483 => "11111110011010110000011111110001",
			484 => "0000001001000000000001111000000100",
			485 => "00000000101101010000011111110001",
			486 => "00000000000000000000011111110001",
			487 => "0000000101000000000000110100010100",
			488 => "0000000100000000001100111100010000",
			489 => "0000001001000000001000010000001000",
			490 => "0000001110000000001110101100000100",
			491 => "00000000000000000000011111110001",
			492 => "00000001010010110000011111110001",
			493 => "0000000110000000000100111100000100",
			494 => "00000000000000000000011111110001",
			495 => "00000000001010000000011111110001",
			496 => "00000000000000000000011111110001",
			497 => "0000001101000000001110101000001000",
			498 => "0000001001000000000000001000000100",
			499 => "11111110100111110000011111110001",
			500 => "00000000000000000000011111110001",
			501 => "0000001101000000001111010000001000",
			502 => "0000001110000000001100000000000100",
			503 => "00000000000000000000011111110001",
			504 => "00000000101100110000011111110001",
			505 => "0000000011000000000110111000000100",
			506 => "11111111011111100000011111110001",
			507 => "00000000010011010000011111110001",
			508 => "0000000110000000001101011000101100",
			509 => "0000000001000000000001000100010100",
			510 => "0000001000000000001001000100010000",
			511 => "0000000101000000000110110100001100",
			512 => "0000001000000000000011101000000100",
			513 => "11111110101110000000100100110101",
			514 => "0000000101000000001100101100000100",
			515 => "00000000000000000000100100110101",
			516 => "00000001111000110000100100110101",
			517 => "11111110011110100000100100110101",
			518 => "11111110011001010000100100110101",
			519 => "0000000011000000001111010100010000",
			520 => "0000000010000000000111011000001100",
			521 => "0000000100000000000111011000000100",
			522 => "00000001110010010000100100110101",
			523 => "0000001111000000001100000000000100",
			524 => "11111110101101100000100100110101",
			525 => "00000000001111010000100100110101",
			526 => "00000010111001110000100100110101",
			527 => "0000000010000000000110111100000100",
			528 => "00000000000000000000100100110101",
			529 => "11111110111011110000100100110101",
			530 => "0000001100000000001000011001010100",
			531 => "0000000110000000001000010000110000",
			532 => "0000000100000000001000000100011100",
			533 => "0000001100000000001001110000001100",
			534 => "0000000110000000001011001100000100",
			535 => "11111110101110010000100100110101",
			536 => "0000001100000000001000111000000100",
			537 => "00000001011110000000100100110101",
			538 => "00000010100100010000100100110101",
			539 => "0000001101000000000001000000001000",
			540 => "0000000100000000001100111000000100",
			541 => "00000000101110110000100100110101",
			542 => "11111110100010010000100100110101",
			543 => "0000001101000000000101110000000100",
			544 => "00000001011000100000100100110101",
			545 => "00000000000110110000100100110101",
			546 => "0000000110000000001011001100000100",
			547 => "11111110011011100000100100110101",
			548 => "0000001100000000000100000000001000",
			549 => "0000001011000000001000111100000100",
			550 => "11111110100010010000100100110101",
			551 => "00000001010100100000100100110101",
			552 => "0000000011000000001000011000000100",
			553 => "11111110101110100000100100110101",
			554 => "00000000000110100000100100110101",
			555 => "0000001010000000000001010100011100",
			556 => "0000000101000000000101110000010000",
			557 => "0000001001000000001001111100001000",
			558 => "0000001000000000000111000100000100",
			559 => "11111111101010000000100100110101",
			560 => "00000001100000110000100100110101",
			561 => "0000001000000000001100000100000100",
			562 => "00000000010100100000100100110101",
			563 => "00000001101010100000100100110101",
			564 => "0000001111000000001101001000001000",
			565 => "0000001100000000001000011000000100",
			566 => "11111110111010100000100100110101",
			567 => "00000001000000100000100100110101",
			568 => "00000001010110110000100100110101",
			569 => "0000000110000000000101010000000100",
			570 => "00000001010000110000100100110101",
			571 => "11111110110001000000100100110101",
			572 => "0000001101000000000110111100001100",
			573 => "0000000001000000000101011100001000",
			574 => "0000000101000000000010000000000100",
			575 => "11111111111100000000100100110101",
			576 => "00000001000100100000100100110101",
			577 => "11111110011011110000100100110101",
			578 => "0000001000000000001000101100010100",
			579 => "0000000010000000001000110100001000",
			580 => "0000001111000000001000011100000100",
			581 => "11111111000110010000100100110101",
			582 => "00000101000010000000100100110101",
			583 => "0000001101000000001111010100000100",
			584 => "11111110100011100000100100110101",
			585 => "0000001001000000000111101100000100",
			586 => "00000010001101110000100100110101",
			587 => "00000000010101100000100100110101",
			588 => "11111110010101100000100100110101",
			589 => "0000000101000000001010111000011000",
			590 => "0000000100000000001111100000000100",
			591 => "11111110011001000000101001001001",
			592 => "0000001101000000000001111100000100",
			593 => "11111110100101100000101001001001",
			594 => "0000001111000000001110000100001100",
			595 => "0000000110000000001011001100001000",
			596 => "0000001100000000000000101000000100",
			597 => "00000000010110110000101001001001",
			598 => "11111111101101100000101001001001",
			599 => "00000001011110010000101001001001",
			600 => "11111110110111000000101001001001",
			601 => "0000000101000000000100011000011100",
			602 => "0000001101000000001011000000010100",
			603 => "0000001011000000000101101100001000",
			604 => "0000000001000000001001111000000100",
			605 => "00000000000000000000101001001001",
			606 => "11111110101001000000101001001001",
			607 => "0000000110000000001101011000000100",
			608 => "00000000000000000000101001001001",
			609 => "0000000010000000000010000100000100",
			610 => "00000001100101010000101001001001",
			611 => "00000000000000000000101001001001",
			612 => "0000000110000000001101011000000100",
			613 => "00000000000000000000101001001001",
			614 => "00000001100110100000101001001001",
			615 => "0000001101000000001000000000011100",
			616 => "0000000100000000000010100100010000",
			617 => "0000001111000000000101110000001100",
			618 => "0000000001000000000110101000001000",
			619 => "0000000000000000001010000000000100",
			620 => "11111101111111110000101001001001",
			621 => "00000000000000000000101001001001",
			622 => "00000000100000000000101001001001",
			623 => "11111101100001110000101001001001",
			624 => "0000000010000000000111010100001000",
			625 => "0000001100000000001100110000000100",
			626 => "00000001000111110000101001001001",
			627 => "00000000000000000000101001001001",
			628 => "00000000000000000000101001001001",
			629 => "0000001011000000001100101100011100",
			630 => "0000001111000000001001011100010000",
			631 => "0000000000000000001111000100001000",
			632 => "0000000101000000000011100000000100",
			633 => "11111111110100000000101001001001",
			634 => "00000000000110110000101001001001",
			635 => "0000000101000000000011100000000100",
			636 => "00000010000101100000101001001001",
			637 => "00000000111010010000101001001001",
			638 => "0000000110000000001001100100000100",
			639 => "11111110110011100000101001001001",
			640 => "0000000010000000001111010100000100",
			641 => "00000001101000000000101001001001",
			642 => "00000000010101000000101001001001",
			643 => "0000001110000000000101100100010000",
			644 => "0000000000000000000001110100001000",
			645 => "0000001100000000000110000100000100",
			646 => "00000000000000000000101001001001",
			647 => "00000000001000010000101001001001",
			648 => "0000000110000000001111000000000100",
			649 => "11111101110011010000101001001001",
			650 => "00000000000000000000101001001001",
			651 => "0000000101000000001001001000001000",
			652 => "0000001010000000000001010000000100",
			653 => "11111111111011010000101001001001",
			654 => "00000001011010110000101001001001",
			655 => "0000001001000000000100110100000100",
			656 => "11111111010100000000101001001001",
			657 => "00000000001111100000101001001001",
			658 => "0000000110000000001010011000100100",
			659 => "0000000001000000000101011100010000",
			660 => "0000001010000000001010100000001100",
			661 => "0000000000000000001100000100000100",
			662 => "11111110011011100000101110000101",
			663 => "0000001110000000001100110000000100",
			664 => "00000000000000000000101110000101",
			665 => "00000010010111110000101110000101",
			666 => "11111110011001000000101110000101",
			667 => "0000000110000000001010011000001100",
			668 => "0000001101000000000010011100001000",
			669 => "0000000111000000000110100100000100",
			670 => "11111110111010100000101110000101",
			671 => "00000001101101010000101110000101",
			672 => "00000100110011110000101110000101",
			673 => "0000001001000000000100101100000100",
			674 => "11111110100011010000101110000101",
			675 => "00000000100000000000101110000101",
			676 => "0000001100000000001000011001010100",
			677 => "0000000110000000001000010000110000",
			678 => "0000000011000000001001110100010000",
			679 => "0000000110000000001001100100000100",
			680 => "11111110011010100000101110000101",
			681 => "0000000111000000001101100000001000",
			682 => "0000001101000000000111001000000100",
			683 => "00000000010101000000101110000101",
			684 => "00000001111010000000101110000101",
			685 => "11111101111111100000101110000101",
			686 => "0000001100000000001000111100010000",
			687 => "0000000110000000001001100100001000",
			688 => "0000001001000000001101011100000100",
			689 => "00000001011111100000101110000101",
			690 => "11111111100111000000101110000101",
			691 => "0000000011000000000000011100000100",
			692 => "00000000110110110000101110000101",
			693 => "00000001100100010000101110000101",
			694 => "0000000011000000001011011100001000",
			695 => "0000000100000000000011010100000100",
			696 => "11111101111011010000101110000101",
			697 => "11111111110111110000101110000101",
			698 => "0000001011000000000000001100000100",
			699 => "00000001011010010000101110000101",
			700 => "00000000000111010000101110000101",
			701 => "0000000100000000000111011100011000",
			702 => "0000001011000000001011110100001100",
			703 => "0000001010000000001001000100000100",
			704 => "00000000000000000000101110000101",
			705 => "0000001001000000001010011000000100",
			706 => "00000000011010000000101110000101",
			707 => "00000001110000100000101110000101",
			708 => "0000001001000000000010101100000100",
			709 => "11111110000110010000101110000101",
			710 => "0000000001000000001101011000000100",
			711 => "00000010010011100000101110000101",
			712 => "00000000010011010000101110000101",
			713 => "0000001001000000001110010100000100",
			714 => "00000001011011100000101110000101",
			715 => "0000000100000000001101110100000100",
			716 => "11111111110000010000101110000101",
			717 => "11111110001101010000101110000101",
			718 => "0000001101000000000110111100001000",
			719 => "0000000110000000001111000000000100",
			720 => "00000000001001110000101110000101",
			721 => "11111110011010100000101110000101",
			722 => "0000000111000000001011011100000100",
			723 => "00010010000000100000101110000101",
			724 => "0000001110000000001110100100010000",
			725 => "0000001011000000000110100000001000",
			726 => "0000001110000000000110111000000100",
			727 => "00000000110101110000101110000101",
			728 => "11111110100101000000101110000101",
			729 => "0000001001000000000011101000000100",
			730 => "00000001000111110000101110000101",
			731 => "00000100110011010000101110000101",
			732 => "0000000000000000001011000100001000",
			733 => "0000001011000000001111010000000100",
			734 => "11111110101111000000101110000101",
			735 => "00000000111010110000101110000101",
			736 => "11111110010100100000101110000101",
			737 => "0000000101000000000111001000011000",
			738 => "0000000100000000000001101100000100",
			739 => "11111110011101110000110010111001",
			740 => "0000001011000000000011011100010000",
			741 => "0000000010000000000111011000000100",
			742 => "11111111001000000000110010111001",
			743 => "0000000010000000000000010000001000",
			744 => "0000000101000000000011011100000100",
			745 => "00000000000000000000110010111001",
			746 => "00000000011000010000110010111001",
			747 => "11111111101011110000110010111001",
			748 => "00000000111101000000110010111001",
			749 => "0000001111000000001111010000111100",
			750 => "0000000111000000001001110000011100",
			751 => "0000001010000000001010110000001100",
			752 => "0000001100000000000100000000000100",
			753 => "11111110100111000000110010111001",
			754 => "0000001100000000000100000000000100",
			755 => "00000001010000000000110010111001",
			756 => "00000000000000000000110010111001",
			757 => "0000001110000000000100001000000100",
			758 => "00000000000000000000110010111001",
			759 => "0000000110000000001101011000000100",
			760 => "00000000000000000000110010111001",
			761 => "0000001100000000000100000000000100",
			762 => "00000001101100000000110010111001",
			763 => "00000000101010100000110010111001",
			764 => "0000001110000000001011011100011000",
			765 => "0000001111000000001110000100001100",
			766 => "0000001011000000000110000100000100",
			767 => "00000000000000000000110010111001",
			768 => "0000000010000000000001000000000100",
			769 => "00000000000000000000110010111001",
			770 => "11111110010101110000110010111001",
			771 => "0000000000000000000100010100000100",
			772 => "11111111101101100000110010111001",
			773 => "0000001011000000000000001100000100",
			774 => "00000000101001010000110010111001",
			775 => "00000000000000000000110010111001",
			776 => "0000000110000000000111101000000100",
			777 => "00000000000000000000110010111001",
			778 => "00000001010001010000110010111001",
			779 => "0000000001000000000110101000100100",
			780 => "0000001111000000000111111100010100",
			781 => "0000000111000000001001110000001000",
			782 => "0000000110000000001011001100000100",
			783 => "11111111100110010000110010111001",
			784 => "00000001011011010000110010111001",
			785 => "0000000000000000000011010000000100",
			786 => "11111101011101010000110010111001",
			787 => "0000001010000000000110011100000100",
			788 => "11111111101000100000110010111001",
			789 => "00000000000000000000110010111001",
			790 => "0000001100000000001000111000001100",
			791 => "0000000100000000000010111000000100",
			792 => "11111101111011110000110010111001",
			793 => "0000000000000000001010000000000100",
			794 => "00000000000000000000110010111001",
			795 => "11111110110001110000110010111001",
			796 => "00000000000000000000110010111001",
			797 => "0000000101000000001000000000001100",
			798 => "0000001101000000001001110100001000",
			799 => "0000001100000000000100000000000100",
			800 => "00000000111100110000110010111001",
			801 => "11111111011000100000110010111001",
			802 => "00000001100000100000110010111001",
			803 => "0000001001000000000111101000001100",
			804 => "0000001101000000000110100100000100",
			805 => "00000000100000110000110010111001",
			806 => "0000000010000000001010000100000100",
			807 => "11111110011101100000110010111001",
			808 => "00000000000000000000110010111001",
			809 => "0000000101000000001000011000000100",
			810 => "00000001100100000000110010111001",
			811 => "0000001101000000001011101100000100",
			812 => "11111111111110100000110010111001",
			813 => "11111110100100100000110010111001",
			814 => "0000001011000000000011011100001100",
			815 => "0000000010000000001111010100000100",
			816 => "11111110011010000000110110001101",
			817 => "0000000000000000001100110000000100",
			818 => "11111111011010100000110110001101",
			819 => "00000001001100000000110110001101",
			820 => "0000001010000000001001101001011000",
			821 => "0000000001000000000111100100110100",
			822 => "0000000000000000000010011000011000",
			823 => "0000000111000000001001110000001000",
			824 => "0000000000000000001111000100000100",
			825 => "11111110111010100000110110001101",
			826 => "11111001111010010000110110001101",
			827 => "0000001100000000001000111100001000",
			828 => "0000001010000000001001000100000100",
			829 => "11111111011001100000110110001101",
			830 => "00000001001011100000110110001101",
			831 => "0000001100000000000110000100000100",
			832 => "11111110001011100000110110001101",
			833 => "00000001000000010000110110001101",
			834 => "0000000100000000000010100100010000",
			835 => "0000001011000000001110001100001000",
			836 => "0000000011000000000000011100000100",
			837 => "11111111010101100000110110001101",
			838 => "00000000100011000000110110001101",
			839 => "0000001011000000001101111000000100",
			840 => "11111011101100110000110110001101",
			841 => "11111110100111100000110110001101",
			842 => "0000001100000000000011011100001000",
			843 => "0000000011000000001010001100000100",
			844 => "00000000110100100000110110001101",
			845 => "00000010000010000000110110001101",
			846 => "11111110101010000000110110001101",
			847 => "0000000101000000000001101000000100",
			848 => "00000001101000010000110110001101",
			849 => "0000001001000000001100011000010000",
			850 => "0000000111000000000001111100001000",
			851 => "0000001010000000000110011100000100",
			852 => "11111101111100000000110110001101",
			853 => "00000000000000000000110110001101",
			854 => "0000000100000000001110000000000100",
			855 => "00000001010000110000110110001101",
			856 => "11111110010110100000110110001101",
			857 => "0000001010000000000010101100001000",
			858 => "0000001001000000000101010000000100",
			859 => "11111111101001100000110110001101",
			860 => "00000001110000110000110110001101",
			861 => "0000001111000000001000110100000100",
			862 => "00000000000100010000110110001101",
			863 => "00000000101101010000110110001101",
			864 => "0000001100000000001000111100000100",
			865 => "00000001001100100000110110001101",
			866 => "11111110000111110000110110001101",
			867 => "0000000100000000000011000000111000",
			868 => "0000001011000000000000011100011000",
			869 => "0000001010000000001001000100010100",
			870 => "0000001000000000001010110000001100",
			871 => "0000000100000000001011101100001000",
			872 => "0000000000000000000110001000000100",
			873 => "11111111000111010000111011011001",
			874 => "00000000000000000000111011011001",
			875 => "00000000101110110000111011011001",
			876 => "0000000100000000000000010000000100",
			877 => "00000000000000000000111011011001",
			878 => "11111110111000110000111011011001",
			879 => "00000000101001110000111011011001",
			880 => "0000000111000000000001101000010100",
			881 => "0000001001000000001010100000010000",
			882 => "0000000001000000000101011100000100",
			883 => "00000000000000000000111011011001",
			884 => "0000000111000000001001001000000100",
			885 => "00000000000000000000111011011001",
			886 => "0000000101000000000111100000000100",
			887 => "00000001001101100000111011011001",
			888 => "00000000000000000000111011011001",
			889 => "00000000000000000000111011011001",
			890 => "0000000110000000001101011000001000",
			891 => "0000000110000000001101011000000100",
			892 => "11111111011110010000111011011001",
			893 => "00000000101011010000111011011001",
			894 => "11111111011001010000111011011001",
			895 => "0000000100000000000110001100111100",
			896 => "0000000001000000000111100100011000",
			897 => "0000000000000000000010011000000100",
			898 => "11111110001100010000111011011001",
			899 => "0000000101000000000100011000001100",
			900 => "0000001000000000001011010100000100",
			901 => "00000000000000000000111011011001",
			902 => "0000000000000000000011111100000100",
			903 => "11111110001110110000111011011001",
			904 => "00000000000000000000111011011001",
			905 => "0000000111000000001101100000000100",
			906 => "00000000111111100000111011011001",
			907 => "00000000000000000000111011011001",
			908 => "0000001011000000000000001100000100",
			909 => "00000001001011100000111011011001",
			910 => "0000000000000000000111000000010000",
			911 => "0000000000000000001010101100001000",
			912 => "0000000100000000001000000100000100",
			913 => "00000000000011000000111011011001",
			914 => "11111111001111100000111011011001",
			915 => "0000000110000000000100111100000100",
			916 => "00000000000000000000111011011001",
			917 => "00000000111000000000111011011001",
			918 => "0000001001000000000111101100001000",
			919 => "0000000100000000001000110100000100",
			920 => "11111111111100000000111011011001",
			921 => "11111101111111010000111011011001",
			922 => "0000001011000000000100010000000100",
			923 => "00000000110111110000111011011001",
			924 => "11111111001110110000111011011001",
			925 => "0000000110000000001101011000000100",
			926 => "11111110110101000000111011011001",
			927 => "0000000111000000001000111000010100",
			928 => "0000000101000000001101010100001100",
			929 => "0000001011000000001000111100000100",
			930 => "11111111110101000000111011011001",
			931 => "0000000100000000000011011000000100",
			932 => "00000000000000000000111011011001",
			933 => "00000000000100100000111011011001",
			934 => "0000001101000000000011100000000100",
			935 => "00000000010101000000111011011001",
			936 => "00000001011100000000111011011001",
			937 => "0000001000000000000111000000010000",
			938 => "0000000100000000001101001000001000",
			939 => "0000001000000000000111000100000100",
			940 => "00000000010000110000111011011001",
			941 => "11111110101000000000111011011001",
			942 => "0000000011000000001010011100000100",
			943 => "11111111011110100000111011011001",
			944 => "00000000011100110000111011011001",
			945 => "0000001110000000000100001000001000",
			946 => "0000001101000000001110110000000100",
			947 => "00000000000000000000111011011001",
			948 => "00000000011001100000111011011001",
			949 => "11111110111101100000111011011001",
			950 => "0000000110000000001010011000101000",
			951 => "0000000001000000000101011100010100",
			952 => "0000001010000000001010100000010000",
			953 => "0000001000000000001000010100001100",
			954 => "0000000100000000001010000100000100",
			955 => "11111110011100110001000000011101",
			956 => "0000000011000000000111010100000100",
			957 => "00000000001011110001000000011101",
			958 => "00000000000000000001000000011101",
			959 => "00000001111010010001000000011101",
			960 => "11111110011001010001000000011101",
			961 => "0000000110000000001010011000001100",
			962 => "0000001101000000000010011100001000",
			963 => "0000000111000000000110100100000100",
			964 => "11111111000011110001000000011101",
			965 => "00000001011000010001000000011101",
			966 => "00000011000011100001000000011101",
			967 => "0000001001000000000100101100000100",
			968 => "11111110101000110001000000011101",
			969 => "00000000010110010001000000011101",
			970 => "0000001010000000001001101001101100",
			971 => "0000000110000000001000010000111100",
			972 => "0000000100000000000011000000011100",
			973 => "0000001001000000000100101100001100",
			974 => "0000000010000000001000001100001000",
			975 => "0000001111000000001111010100000100",
			976 => "00000001011110010001000000011101",
			977 => "11111110101110110001000000011101",
			978 => "00000011010011100001000000011101",
			979 => "0000000101000000001100100100001000",
			980 => "0000001110000000000010000100000100",
			981 => "11111110100010110001000000011101",
			982 => "00000001110011000001000000011101",
			983 => "0000001101000000001001011100000100",
			984 => "11111110011101010001000000011101",
			985 => "00000001110110010001000000011101",
			986 => "0000001100000000001000111100010000",
			987 => "0000001101000000001110110000001000",
			988 => "0000000100000000001100111100000100",
			989 => "11111110100111110001000000011101",
			990 => "00000001010101100001000000011101",
			991 => "0000000110000000001001100100000100",
			992 => "00000000010001110001000000011101",
			993 => "00000001010011110001000000011101",
			994 => "0000000011000000001011011100001000",
			995 => "0000000100000000000011010100000100",
			996 => "11111110000001100001000000011101",
			997 => "11111111110101010001000000011101",
			998 => "0000000101000000001001110100000100",
			999 => "00000001001100110001000000011101",
			1000 => "11111111110100110001000000011101",
			1001 => "0000000111000000001111011100010100",
			1002 => "0000000100000000000111011100001100",
			1003 => "0000001001000000001010011000000100",
			1004 => "00000000001011110001000000011101",
			1005 => "0000001000000000000001110000000100",
			1006 => "00000000000000000001000000011101",
			1007 => "00000001101101010001000000011101",
			1008 => "0000000001000000001101011100000100",
			1009 => "00000001000000110001000000011101",
			1010 => "11111110100000110001000000011101",
			1011 => "0000001110000000000010110000010000",
			1012 => "0000001101000000000111010100001000",
			1013 => "0000000101000000000111111100000100",
			1014 => "00000000000010010001000000011101",
			1015 => "11111110100110100001000000011101",
			1016 => "0000001100000000000001011000000100",
			1017 => "00000010011111010001000000011101",
			1018 => "00000000000000000001000000011101",
			1019 => "0000000111000000000110110100000100",
			1020 => "00000010010010000001000000011101",
			1021 => "0000000100000000000001101100000100",
			1022 => "11111111100010110001000000011101",
			1023 => "00000001011101110001000000011101",
			1024 => "0000001100000000000100000000000100",
			1025 => "00000000100010110001000000011101",
			1026 => "0000001001000000001011101000001000",
			1027 => "0000000001000000001100100000000100",
			1028 => "11111110100101110001000000011101",
			1029 => "00000000011110100001000000011101",
			1030 => "11111110001011100001000000011101",
			1031 => "0000001011000000000011011100010000",
			1032 => "0000000010000000000111011000000100",
			1033 => "11111110100101000001000100101001",
			1034 => "0000000010000000000000010000001000",
			1035 => "0000001101000000000001111100000100",
			1036 => "00000000000000000001000100101001",
			1037 => "00000000001001000001000100101001",
			1038 => "11111111101101000001000100101001",
			1039 => "0000001011000000001100101100111000",
			1040 => "0000001101000000000110100100110000",
			1041 => "0000000100000000000010111000010100",
			1042 => "0000001000000000000111000100010000",
			1043 => "0000000011000000000000011100001000",
			1044 => "0000000111000000000100000000000100",
			1045 => "00000000000000000001000100101001",
			1046 => "11111110100100100001000100101001",
			1047 => "0000000010000000001110110100000100",
			1048 => "00000001011101000001000100101001",
			1049 => "11111111101010010001000100101001",
			1050 => "11111110011100010001000100101001",
			1051 => "0000001100000000000100000000001100",
			1052 => "0000000010000000001010000100001000",
			1053 => "0000000101000000000111001000000100",
			1054 => "00000000011011110001000100101001",
			1055 => "00000001100110000001000100101001",
			1056 => "00000000000000000001000100101001",
			1057 => "0000000011000000001010011100001000",
			1058 => "0000000100000000000010010000000100",
			1059 => "11111110100001010001000100101001",
			1060 => "00000000100000110001000100101001",
			1061 => "0000000010000000001111010100000100",
			1062 => "00000001000000110001000100101001",
			1063 => "11111111101101010001000100101001",
			1064 => "0000001010000000000001010000000100",
			1065 => "00000000000000000001000100101001",
			1066 => "00000001100111100001000100101001",
			1067 => "0000001100000000000100000000001100",
			1068 => "0000000100000000000110001100001000",
			1069 => "0000000110000000001001100100000100",
			1070 => "00000000000000000001000100101001",
			1071 => "00000000111100000001000100101001",
			1072 => "11111101101110000001000100101001",
			1073 => "0000000100000000001110100100010100",
			1074 => "0000001000000000001011010100010000",
			1075 => "0000001100000000001110001100001000",
			1076 => "0000000100000000000010010100000100",
			1077 => "00000000000000000001000100101001",
			1078 => "11111110010011110001000100101001",
			1079 => "0000001010000000001000100100000100",
			1080 => "00000000000000000001000100101001",
			1081 => "00000000111100000001000100101001",
			1082 => "00000001100101100001000100101001",
			1083 => "0000000011000000000110111000010000",
			1084 => "0000001010000000001010110000001000",
			1085 => "0000000000000000001111000100000100",
			1086 => "11111111100010010001000100101001",
			1087 => "11111110000110110001000100101001",
			1088 => "0000000100000000000000010100000100",
			1089 => "00000001000100010001000100101001",
			1090 => "11111111001010000001000100101001",
			1091 => "0000001000000000000001110100001000",
			1092 => "0000001000000000000001010100000100",
			1093 => "11111111010101110001000100101001",
			1094 => "00000000101010000001000100101001",
			1095 => "0000000100000000000001101100000100",
			1096 => "11111110111111100001000100101001",
			1097 => "00000000111010100001000100101001",
			1098 => "0000001001000000000001111001000000",
			1099 => "0000000111000000001101100000101000",
			1100 => "0000001100000000001001110000100000",
			1101 => "0000001111000000001001100000011100",
			1102 => "0000000001000000000110101000010000",
			1103 => "0000000100000000000010111000001000",
			1104 => "0000001111000000000101110000000100",
			1105 => "00000000000000000001001001010101",
			1106 => "11111110001000100001001001010101",
			1107 => "0000001101000000001011000000000100",
			1108 => "11111111110110000001001001010101",
			1109 => "00000001000110010001001001010101",
			1110 => "0000000110000000001011001100000100",
			1111 => "11111111011000100001001001010101",
			1112 => "0000000111000000001001110000000100",
			1113 => "00000000000000000001001001010101",
			1114 => "00000001100001110001001001010101",
			1115 => "11111110101010010001001001010101",
			1116 => "0000001010000000000101000100000100",
			1117 => "11111110000111000001001001010101",
			1118 => "00000000000000000001001001010101",
			1119 => "0000000111000000001110001100001000",
			1120 => "0000000010000000001100111000000100",
			1121 => "11111110100111110001001001010101",
			1122 => "00000000000000000001001001010101",
			1123 => "0000001010000000000001110000001100",
			1124 => "0000000101000000000111010000000100",
			1125 => "00000000000000000001001001010101",
			1126 => "0000000010000000001110010000000100",
			1127 => "00000000000000000001001001010101",
			1128 => "00000000111100000001001001010101",
			1129 => "11111111010111010001001001010101",
			1130 => "0000000101000000001010011100000100",
			1131 => "00000001100001000001001001010101",
			1132 => "0000000011000000000010000000011000",
			1133 => "0000000100000000001010110100001000",
			1134 => "0000000010000000001100010000000100",
			1135 => "00000000000000000001001001010101",
			1136 => "11111110011010000001001001010101",
			1137 => "0000000100000000001100111100001100",
			1138 => "0000000111000000001101111000001000",
			1139 => "0000000010000000001111100100000100",
			1140 => "00000000000000000001001001010101",
			1141 => "00000001010100110001001001010101",
			1142 => "00000000000000000001001001010101",
			1143 => "11111111100100000001001001010101",
			1144 => "0000000011000000001010000100011100",
			1145 => "0000001111000000001111010100010000",
			1146 => "0000001000000000001000100100001000",
			1147 => "0000000001000000000101011100000100",
			1148 => "00000000000000000001001001010101",
			1149 => "00000001000001110001001001010101",
			1150 => "0000000001000000001011111100000100",
			1151 => "11111111001000110001001001010101",
			1152 => "00000000000000000001001001010101",
			1153 => "0000000010000000000010010100001000",
			1154 => "0000001001000000000000001000000100",
			1155 => "00000001100101110001001001010101",
			1156 => "00000000000000000001001001010101",
			1157 => "11111111110111110001001001010101",
			1158 => "0000000101000000001101000100010000",
			1159 => "0000001100000000000100011000001000",
			1160 => "0000000001000000001011111100000100",
			1161 => "00000000000000000001001001010101",
			1162 => "00000001000110010001001001010101",
			1163 => "0000000110000000000100111100000100",
			1164 => "11111111000100100001001001010101",
			1165 => "00000000011110100001001001010101",
			1166 => "0000001100000000000100011000001000",
			1167 => "0000000001000000000100110100000100",
			1168 => "11111110111100110001001001010101",
			1169 => "00000000000000000001001001010101",
			1170 => "0000001100000000001011000000000100",
			1171 => "00000000110010110001001001010101",
			1172 => "00000000000000000001001001010101",
			1173 => "0000001111000000001011110001111000",
			1174 => "0000001111000000000010010101100100",
			1175 => "0000001111000000000101110000111000",
			1176 => "0000000011000000001010011100011100",
			1177 => "0000000100000000000000101100010000",
			1178 => "0000000111000000001000111000001000",
			1179 => "0000000101000000001101010100000100",
			1180 => "11111111000101000001001111000001",
			1181 => "00000000110100110001001111000001",
			1182 => "0000001011000000000001111100000100",
			1183 => "11111110101101010001001111000001",
			1184 => "00000000000000000001001111000001",
			1185 => "0000000101000000000100011000001000",
			1186 => "0000001101000000000111001000000100",
			1187 => "00000000000000000001001111000001",
			1188 => "00000001000101110001001111000001",
			1189 => "11111111011111110001001111000001",
			1190 => "0000000111000000001001110000001100",
			1191 => "0000001101000000000011100000000100",
			1192 => "00000000000000000001001111000001",
			1193 => "0000000110000000001101011000000100",
			1194 => "00000000000000000001001111000001",
			1195 => "00000001010000110001001111000001",
			1196 => "0000001000000000000001110100001000",
			1197 => "0000000001000000000111100100000100",
			1198 => "11111110110111010001001111000001",
			1199 => "00000000000000000001001111000001",
			1200 => "0000001100000000001001110000000100",
			1201 => "00000000101001100001001111000001",
			1202 => "00000000000000000001001111000001",
			1203 => "0000000011000000000101110100010100",
			1204 => "0000000110000000001111000000001100",
			1205 => "0000001011000000001100101100001000",
			1206 => "0000000100000000000011110000000100",
			1207 => "00000000010011010001001111000001",
			1208 => "11111111001001010001001111000001",
			1209 => "11111110010101010001001111000001",
			1210 => "0000000100000000001110111000000100",
			1211 => "00000000000000000001001111000001",
			1212 => "00000000100101000001001111000001",
			1213 => "0000001011000000001100101100001000",
			1214 => "0000001000000000001001101000000100",
			1215 => "00000000000000000001001111000001",
			1216 => "00000001010011110001001111000001",
			1217 => "0000000001000000000111100100001000",
			1218 => "0000000011000000001001010100000100",
			1219 => "11111111111101110001001111000001",
			1220 => "00000001010010110001001111000001",
			1221 => "0000000011000000000010000000000100",
			1222 => "11111111011100100001001111000001",
			1223 => "00000000000000000001001111000001",
			1224 => "0000000001000000000001111000000100",
			1225 => "11111110001000010001001111000001",
			1226 => "0000001011000000000010001000000100",
			1227 => "00000000010001110001001111000001",
			1228 => "0000001011000000000001001000000100",
			1229 => "11111111010101000001001111000001",
			1230 => "0000000100000000001000011100000100",
			1231 => "00000000000000000001001111000001",
			1232 => "00000000000001000001001111000001",
			1233 => "0000001010000000000110011100101100",
			1234 => "0000001011000000000100010000001000",
			1235 => "0000001111000000001110000000000100",
			1236 => "00000000000000000001001111000001",
			1237 => "00000001011000010001001111000001",
			1238 => "0000000100000000000010100100011100",
			1239 => "0000001011000000000110100000010000",
			1240 => "0000000100000000001110100100001000",
			1241 => "0000000001000000001100011000000100",
			1242 => "00000000111001010001001111000001",
			1243 => "00000000000000000001001111000001",
			1244 => "0000000001000000001110010100000100",
			1245 => "00000000000000000001001111000001",
			1246 => "11111111000101010001001111000001",
			1247 => "0000001000000000001001101000001000",
			1248 => "0000001101000000001111010100000100",
			1249 => "00000000000000000001001111000001",
			1250 => "00000000111100110001001111000001",
			1251 => "00000000000000000001001111000001",
			1252 => "0000000000000000000000111000000100",
			1253 => "00000001010000010001001111000001",
			1254 => "00000000000000000001001111000001",
			1255 => "0000001111000000001011001000001100",
			1256 => "0000000010000000001101001000000100",
			1257 => "00000000000000000001001111000001",
			1258 => "0000000110000000000100101100000100",
			1259 => "00000000000000000001001111000001",
			1260 => "11111110011100000001001111000001",
			1261 => "0000001010000000001001101000000100",
			1262 => "00000001000110000001001111000001",
			1263 => "00000000000000000001001111000001",
			1264 => "0000000110000000001011001101100000",
			1265 => "0000001111000000000110111100111100",
			1266 => "0000000110000000001101011000100100",
			1267 => "0000000001000000000101011100010000",
			1268 => "0000000001000000000110101000000100",
			1269 => "11111110010100010001010101100101",
			1270 => "0000001001000000001001011000000100",
			1271 => "00000010110011010001010101100101",
			1272 => "0000001000000000001000010100000100",
			1273 => "11111110010111010001010101100101",
			1274 => "11111111111010010001010101100101",
			1275 => "0000001000000000001000100100000100",
			1276 => "00000101010100010001010101100101",
			1277 => "0000001110000000000110010000001000",
			1278 => "0000001001000000000101010000000100",
			1279 => "00000001101010000001010101100101",
			1280 => "11111110011000100001010101100101",
			1281 => "0000001101000000001111010000000100",
			1282 => "00000101100111010001010101100101",
			1283 => "11111110011101010001010101100101",
			1284 => "0000000010000000001110110100010100",
			1285 => "0000000011000000001001110100000100",
			1286 => "11111110010111000001010101100101",
			1287 => "0000000100000000000010110000001000",
			1288 => "0000000011000000000001011000000100",
			1289 => "11111110011111010001010101100101",
			1290 => "00000100001011010001010101100101",
			1291 => "0000001100000000001000111000000100",
			1292 => "00001011101100110001010101100101",
			1293 => "00000000111111100001010101100101",
			1294 => "11111110010110000001010101100101",
			1295 => "0000001100000000000100011000010000",
			1296 => "0000000010000000001111010100000100",
			1297 => "00001010100000100001010101100101",
			1298 => "0000001111000000000000010000001000",
			1299 => "0000000111000000000001101000000100",
			1300 => "11111110011100010001010101100101",
			1301 => "00000000110110000001010101100101",
			1302 => "00000101000101100001010101100101",
			1303 => "0000000100000000001101101100001100",
			1304 => "0000001011000000001011011100001000",
			1305 => "0000001000000000000001010000000100",
			1306 => "00000100110011010001010101100101",
			1307 => "11111110011111100001010101100101",
			1308 => "11111110010111010001010101100101",
			1309 => "0000000100000000000011000000000100",
			1310 => "00001010001001110001010101100101",
			1311 => "00000000001011010001010101100101",
			1312 => "0000001100000000000110100101001000",
			1313 => "0000001010000000001000010100100000",
			1314 => "0000000110000000001111000000010000",
			1315 => "0000001001000000001001111100000100",
			1316 => "00000110010100110001010101100101",
			1317 => "0000001010000000000011101000000100",
			1318 => "00000011010010100001010101100101",
			1319 => "0000000111000000000110100100000100",
			1320 => "11111110100000000001010101100101",
			1321 => "11111111101100110001010101100101",
			1322 => "0000000111000000001001001000000100",
			1323 => "00001000111001000001010101100101",
			1324 => "0000000110000000000100111100000100",
			1325 => "00000101111110110001010101100101",
			1326 => "0000000001000000000100110100000100",
			1327 => "11111111101011100001010101100101",
			1328 => "00000100001000010001010101100101",
			1329 => "0000000100000000000011111000100000",
			1330 => "0000000110000000001001100100010000",
			1331 => "0000000111000000000101101100001000",
			1332 => "0000001011000000000011011100000100",
			1333 => "11111110100011000001010101100101",
			1334 => "00000101110101010001010101100101",
			1335 => "0000001000000000001100000100000100",
			1336 => "00000010100001100001010101100101",
			1337 => "11111110011000000001010101100101",
			1338 => "0000000111000000000111010000001000",
			1339 => "0000000111000000001101100000000100",
			1340 => "00000110100111010001010101100101",
			1341 => "00000101101100110001010101100101",
			1342 => "0000000010000000001100001100000100",
			1343 => "11111110011110010001010101100101",
			1344 => "00000100100101100001010101100101",
			1345 => "0000001100000000001000111100000100",
			1346 => "00000011000001010001010101100101",
			1347 => "11111110011010100001010101100101",
			1348 => "0000001100000000001000011000011000",
			1349 => "0000000110000000000101010000010000",
			1350 => "0000000001000000001100011000001100",
			1351 => "0000000111000000000101100100001000",
			1352 => "0000001001000000001010100000000100",
			1353 => "11111110100000110001010101100101",
			1354 => "00000000111110000001010101100101",
			1355 => "00000110000010100001010101100101",
			1356 => "11111110010110000001010101100101",
			1357 => "0000000001000000001100011000000100",
			1358 => "00000000001101010001010101100101",
			1359 => "00001011010001000001010101100101",
			1360 => "0000000001000000001000010000010000",
			1361 => "0000001001000000001000010100001100",
			1362 => "0000000110000000001111000000000100",
			1363 => "00000000000000000001010101100101",
			1364 => "0000000111000000000000011100000100",
			1365 => "11111111010000000001010101100101",
			1366 => "11111110011010000001010101100101",
			1367 => "00000000000010010001010101100101",
			1368 => "00000011101010100001010101100101",
			1369 => "0000000110000000001001100101010100",
			1370 => "0000000101000000000111001000000100",
			1371 => "11111110100110010001011010100001",
			1372 => "0000001111000000001110000100100100",
			1373 => "0000001010000000001010110000010100",
			1374 => "0000000010000000000001000000001100",
			1375 => "0000001100000000000110000100000100",
			1376 => "00000000000000000001011010100001",
			1377 => "0000000101000000001011011100000100",
			1378 => "00000000101111000001011010100001",
			1379 => "00000000000000000001011010100001",
			1380 => "0000001111000000000001000000000100",
			1381 => "11111110110100010001011010100001",
			1382 => "00000000000000000001011010100001",
			1383 => "0000000110000000001101011000000100",
			1384 => "00000000000000000001011010100001",
			1385 => "0000001100000000001000111000001000",
			1386 => "0000001110000000000100001000000100",
			1387 => "00000000000000000001011010100001",
			1388 => "00000001010011000001011010100001",
			1389 => "00000000000000000001011010100001",
			1390 => "0000000100000000001000000100011000",
			1391 => "0000001001000000001110010100001000",
			1392 => "0000000100000000001011110000000100",
			1393 => "00000000000000000001011010100001",
			1394 => "00000001000111110001011010100001",
			1395 => "0000001001000000000111101100001000",
			1396 => "0000000111000000000111010000000100",
			1397 => "11111111010001100001011010100001",
			1398 => "00000000001001100001011010100001",
			1399 => "0000001000000000001010110000000100",
			1400 => "00000000110100010001011010100001",
			1401 => "11111111101110010001011010100001",
			1402 => "0000000010000000001100010000001100",
			1403 => "0000000010000000000110010000000100",
			1404 => "11111111011010010001011010100001",
			1405 => "0000001100000000001000111000000100",
			1406 => "00000000001010110001011010100001",
			1407 => "00000000000000000001011010100001",
			1408 => "0000001100000000000111001000000100",
			1409 => "11111110011001100001011010100001",
			1410 => "00000000000000000001011010100001",
			1411 => "0000000111000000001101100000011000",
			1412 => "0000001011000000001100101100010100",
			1413 => "0000001111000000001110010000010000",
			1414 => "0000001001000000001001011000001100",
			1415 => "0000000100000000000100001100000100",
			1416 => "11111110110000100001011010100001",
			1417 => "0000000010000000001010000100000100",
			1418 => "00000001010100110001011010100001",
			1419 => "00000000000000000001011010100001",
			1420 => "00000001011011110001011010100001",
			1421 => "11111111000101110001011010100001",
			1422 => "00000001100011010001011010100001",
			1423 => "0000001100000000000100000000001000",
			1424 => "0000001000000000001011010100000100",
			1425 => "00000000000000000001011010100001",
			1426 => "11111110010100000001011010100001",
			1427 => "0000000000000000000111111000011100",
			1428 => "0000001010000000001100011100010000",
			1429 => "0000001000000000000111000100001000",
			1430 => "0000001100000000001001110000000100",
			1431 => "00000001000110000001011010100001",
			1432 => "11111111111110010001011010100001",
			1433 => "0000001111000000000110010000000100",
			1434 => "00000000000000000001011010100001",
			1435 => "11111101011110100001011010100001",
			1436 => "0000001100000000001000000000000100",
			1437 => "00000001100100000001011010100001",
			1438 => "0000001111000000000000010100000100",
			1439 => "11111110100111100001011010100001",
			1440 => "00000000110101110001011010100001",
			1441 => "0000000111000000001101100000000100",
			1442 => "00000000001010010001011010100001",
			1443 => "0000001110000000001011001000000100",
			1444 => "11111110100000100001011010100001",
			1445 => "0000001100000000000101110100000100",
			1446 => "00000000001011100001011010100001",
			1447 => "00000000000000000001011010100001",
			1448 => "0000001110000000001110101101010100",
			1449 => "0000001011000000001100101100101100",
			1450 => "0000000100000000001000000100001100",
			1451 => "0000001100000000000100000000000100",
			1452 => "00000000000000000001100000010101",
			1453 => "0000001101000000001001110100000100",
			1454 => "11111110100000100001100000010101",
			1455 => "00000000000000000001100000010101",
			1456 => "0000000011000000000000011100010000",
			1457 => "0000001010000000001010110000000100",
			1458 => "11111110111001110001100000010101",
			1459 => "0000001111000000001001010000001000",
			1460 => "0000000011000000001001110100000100",
			1461 => "11111111101100010001100000010101",
			1462 => "00000000101010000001100000010101",
			1463 => "11111111000111110001100000010101",
			1464 => "0000001111000000001110010000001000",
			1465 => "0000001101000000001011000000000100",
			1466 => "00000000000000000001100000010101",
			1467 => "00000001011001010001100000010101",
			1468 => "0000001101000000000110100100000100",
			1469 => "11111110110100010001100000010101",
			1470 => "00000000100010010001100000010101",
			1471 => "0000000001000000000111100100010100",
			1472 => "0000001101000000001001001000000100",
			1473 => "00000000000000000001100000010101",
			1474 => "0000000110000000001000010000001100",
			1475 => "0000000110000000001001011000000100",
			1476 => "00000000000000000001100000010101",
			1477 => "0000001010000000000110011100000100",
			1478 => "11111110011110110001100000010101",
			1479 => "00000000000000000001100000010101",
			1480 => "00000000000000000001100000010101",
			1481 => "0000001011000000000000001100000100",
			1482 => "00000000100001100001100000010101",
			1483 => "0000000110000000001101011000001100",
			1484 => "0000001100000000001110001100000100",
			1485 => "00000000000000000001100000010101",
			1486 => "0000001101000000000001011000000100",
			1487 => "00000000011001010001100000010101",
			1488 => "00000000000000000001100000010101",
			1489 => "11111111001111000001100000010101",
			1490 => "0000001111000000001111100100110100",
			1491 => "0000000110000000000100111100110000",
			1492 => "0000001111000000000110111100011000",
			1493 => "0000000010000000001100010000010000",
			1494 => "0000001110000000000101001000001000",
			1495 => "0000000111000000000011100000000100",
			1496 => "00000000110101110001100000010101",
			1497 => "00000000000000000001100000010101",
			1498 => "0000001011000000000101100100000100",
			1499 => "11111111101010010001100000010101",
			1500 => "00000000000000000001100000010101",
			1501 => "0000001011000000000000001100000100",
			1502 => "00000000000000000001100000010101",
			1503 => "11111110110111000001100000010101",
			1504 => "0000000011000000001010000100001100",
			1505 => "0000000001000000001101111100001000",
			1506 => "0000000011000000001100010000000100",
			1507 => "00000000000000000001100000010101",
			1508 => "00000000111011010001100000010101",
			1509 => "00000000000000000001100000010101",
			1510 => "0000000111000000000110100100000100",
			1511 => "11111111011101100001100000010101",
			1512 => "0000000100000000001111100100000100",
			1513 => "00000000000000000001100000010101",
			1514 => "00000000011101010001100000010101",
			1515 => "00000001000101100001100000010101",
			1516 => "0000000011000000001110110100000100",
			1517 => "11111110111011110001100000010101",
			1518 => "0000000001000000000111101000010100",
			1519 => "0000001000000000000010101000001100",
			1520 => "0000001000000000001011010100001000",
			1521 => "0000001010000000000110011000000100",
			1522 => "00000000011111000001100000010101",
			1523 => "11111111010001000001100000010101",
			1524 => "00000001000000010001100000010101",
			1525 => "0000000001000000000000111100000100",
			1526 => "00000000000000000001100000010101",
			1527 => "11111111110011010001100000010101",
			1528 => "0000000001000000000001111000001100",
			1529 => "0000001010000000001100011100001000",
			1530 => "0000001011000000001011011100000100",
			1531 => "00000000000000000001100000010101",
			1532 => "11111110010011100001100000010101",
			1533 => "00000000000000000001100000010101",
			1534 => "0000000100000000000100001100001000",
			1535 => "0000000000000000000001110100000100",
			1536 => "11111111100110110001100000010101",
			1537 => "00000000011010000001100000010101",
			1538 => "0000001010000000000001010100000100",
			1539 => "11111111000011100001100000010101",
			1540 => "00000000000111000001100000010101",
			1541 => "0000000110000000001011001101011000",
			1542 => "0000001001000000001000010000110100",
			1543 => "0000000110000000001011001100100000",
			1544 => "0000000110000000001001011000001000",
			1545 => "0000000000000000001100000100000100",
			1546 => "11111110011111110001100110110001",
			1547 => "00000011010001110001100110110001",
			1548 => "0000000110000000001101011000001100",
			1549 => "0000001110000000001011011100000100",
			1550 => "11111110010111010001100110110001",
			1551 => "0000001101000000000100010000000100",
			1552 => "00000001001000000001100110110001",
			1553 => "11111110011000000001100110110001",
			1554 => "0000001110000000001011000000000100",
			1555 => "11111110011011000001100110110001",
			1556 => "0000001110000000000110100100000100",
			1557 => "00000010001000100001100110110001",
			1558 => "11111110100100000001100110110001",
			1559 => "0000000010000000000010000100010000",
			1560 => "0000001110000000001010111000000100",
			1561 => "11111110011110000001100110110001",
			1562 => "0000001010000000001010110000001000",
			1563 => "0000000000000000000010011000000100",
			1564 => "00000000101001010001100110110001",
			1565 => "11111110011111010001100110110001",
			1566 => "00000010111000110001100110110001",
			1567 => "11111110011010100001100110110001",
			1568 => "0000001110000000001110110100001100",
			1569 => "0000000111000000001110110000001000",
			1570 => "0000000100000000001100111000000100",
			1571 => "00000100111111000001100110110001",
			1572 => "11111110110000010001100110110001",
			1573 => "11111110011010000001100110110001",
			1574 => "0000001100000000000100011000001000",
			1575 => "0000000101000000000110100000000100",
			1576 => "00000000010010110001100110110001",
			1577 => "11111110010011000001100110110001",
			1578 => "0000000100000000001101101100001100",
			1579 => "0000000101000000000111100000001000",
			1580 => "0000001010000000000010101100000100",
			1581 => "00000011011010010001100110110001",
			1582 => "11111111101001110001100110110001",
			1583 => "11111110011110000001100110110001",
			1584 => "00000101001010010001100110110001",
			1585 => "0000001011000000000001001001001100",
			1586 => "0000001000000000000001010100100000",
			1587 => "0000000100000000001000110100011100",
			1588 => "0000001001000000000111101100001100",
			1589 => "0000001100000000000100011000001000",
			1590 => "0000000110000000001011001100000100",
			1591 => "11111110001111000001100110110001",
			1592 => "00000001100100000001100110110001",
			1593 => "00000100011101000001100110110001",
			1594 => "0000001010000000000111110100001000",
			1595 => "0000001010000000000011101000000100",
			1596 => "00000000010100100001100110110001",
			1597 => "11111110011001010001100110110001",
			1598 => "0000001011000000000110110100000100",
			1599 => "00000010000100110001100110110001",
			1600 => "11111111000000000001100110110001",
			1601 => "11111110010000110001100110110001",
			1602 => "0000000100000000000100001100010100",
			1603 => "0000001101000000001110110000000100",
			1604 => "11111110001010100001100110110001",
			1605 => "0000000001000000001011101000001000",
			1606 => "0000000111000000000101101100000100",
			1607 => "00000010000010100001100110110001",
			1608 => "11111110110011110001100110110001",
			1609 => "0000000000000000001010101100000100",
			1610 => "00000000001111110001100110110001",
			1611 => "00000010001100100001100110110001",
			1612 => "0000001100000000001000111000001100",
			1613 => "0000000101000000000100001000000100",
			1614 => "11111110100000010001100110110001",
			1615 => "0000001001000000001101101000000100",
			1616 => "00000011111000100001100110110001",
			1617 => "00000001111100100001100110110001",
			1618 => "0000000110000000001111000000000100",
			1619 => "11111110011001000001100110110001",
			1620 => "0000001100000000000110000100000100",
			1621 => "00000001100000110001100110110001",
			1622 => "11111111000010110001100110110001",
			1623 => "0000001001000000001000100100100100",
			1624 => "0000000111000000000001011000001100",
			1625 => "0000001101000000001100010000000100",
			1626 => "11111110011011100001100110110001",
			1627 => "0000001110000000001000000100000100",
			1628 => "00000110100110000001100110110001",
			1629 => "00000000100001000001100110110001",
			1630 => "0000000001000000000001111000001100",
			1631 => "0000001010000000001010110000001000",
			1632 => "0000001101000000000110111100000100",
			1633 => "00000000011011010001100110110001",
			1634 => "00000110011111110001100110110001",
			1635 => "11111110011000010001100110110001",
			1636 => "0000001101000000001010000100000100",
			1637 => "11111110010111110001100110110001",
			1638 => "0000001110000000001110100100000100",
			1639 => "00000110011100100001100110110001",
			1640 => "11111110011110100001100110110001",
			1641 => "0000001110000000000000010100000100",
			1642 => "11111110100010010001100110110001",
			1643 => "00000010001000100001100110110001",
			1644 => "0000000110000000001011001100111100",
			1645 => "0000000001000000000101011100011100",
			1646 => "0000000110000000001001011000001000",
			1647 => "0000000001000000000111100100000100",
			1648 => "11111110100001010001101100100101",
			1649 => "00000010110101100001101100100101",
			1650 => "0000001110000000001011000000000100",
			1651 => "11111110010111110001101100100101",
			1652 => "0000001101000000000100010000001100",
			1653 => "0000000111000000001101010100001000",
			1654 => "0000000000000000001110111100000100",
			1655 => "11111110110001010001101100100101",
			1656 => "00000001110001010001101100100101",
			1657 => "00000101000011010001101100100101",
			1658 => "11111110011000010001101100100101",
			1659 => "0000001111000000001111010100010000",
			1660 => "0000001110000000000111111100000100",
			1661 => "00000001100101000001101100100101",
			1662 => "0000001110000000001110110100000100",
			1663 => "11111110011100000001101100100101",
			1664 => "0000000101000000001101000100000100",
			1665 => "00000001011011000001101100100101",
			1666 => "11111110100101100001101100100101",
			1667 => "0000000101000000000101110000001100",
			1668 => "0000000101000000000111100000001000",
			1669 => "0000000101000000001100100100000100",
			1670 => "00000000011100010001101100100101",
			1671 => "00000101100011100001101100100101",
			1672 => "11111110011100000001101100100101",
			1673 => "00000101000001010001101100100101",
			1674 => "0000001100000000001000011001011100",
			1675 => "0000000110000000001000010000111000",
			1676 => "0000000111000000001101100000011100",
			1677 => "0000001101000000001110110000001100",
			1678 => "0000000100000000000000101100001000",
			1679 => "0000001111000000000000110100000100",
			1680 => "11111111111101110001101100100101",
			1681 => "11111110001111010001101100100101",
			1682 => "00000010010101010001101100100101",
			1683 => "0000001111000000001001011100001000",
			1684 => "0000001101000000001011000000000100",
			1685 => "00000001100101000001101100100101",
			1686 => "00000010011111110001101100100101",
			1687 => "0000001001000000001001011000000100",
			1688 => "11111101100011110001101100100101",
			1689 => "00000001101011010001101100100101",
			1690 => "0000000101000000000010110100010000",
			1691 => "0000000100000000001111101000001000",
			1692 => "0000000001000000001110010100000100",
			1693 => "00000011000001010001101100100101",
			1694 => "11111110100010000001101100100101",
			1695 => "0000000111000000000101101100000100",
			1696 => "00000000100011110001101100100101",
			1697 => "11111110011001010001101100100101",
			1698 => "0000000001000000001100011000001000",
			1699 => "0000000000000000000110001000000100",
			1700 => "11111111110111000001101100100101",
			1701 => "00000001100010110001101100100101",
			1702 => "11111110001011100001101100100101",
			1703 => "0000000000000000001010101100001000",
			1704 => "0000001111000000001111101000000100",
			1705 => "00000000100000000001101100100101",
			1706 => "11111101111111010001101100100101",
			1707 => "0000001011000000001011110100010000",
			1708 => "0000000100000000000100001100001000",
			1709 => "0000000001000000001011101000000100",
			1710 => "00000001011100010001101100100101",
			1711 => "00000010001000010001101100100101",
			1712 => "0000001100000000001110001100000100",
			1713 => "00000001111010110001101100100101",
			1714 => "11111110110001000001101100100101",
			1715 => "0000000110000000001000010000000100",
			1716 => "00000101100111010001101100100101",
			1717 => "0000001111000000001000001000000100",
			1718 => "11111110100010010001101100100101",
			1719 => "00000001111000100001101100100101",
			1720 => "0000000001000000001000010000100000",
			1721 => "0000001010000000000110011100011100",
			1722 => "0000000001000000000111101000010000",
			1723 => "0000001101000000000110111100001000",
			1724 => "0000000100000000000100001100000100",
			1725 => "11111110100010100001101100100101",
			1726 => "00000010111111100001101100100101",
			1727 => "0000001010000000000001010000000100",
			1728 => "00001100101001110001101100100101",
			1729 => "00000010101010100001101100100101",
			1730 => "0000000100000000000011101100001000",
			1731 => "0000001101000000001010000100000100",
			1732 => "11111110011110000001101100100101",
			1733 => "11111111110000110001101100100101",
			1734 => "00000010111100100001101100100101",
			1735 => "11111110010111100001101100100101",
			1736 => "00000001101000010001101100100101",
			1737 => "0000001011000000000011011100001100",
			1738 => "0000000010000000001111010100000100",
			1739 => "11111110011010010001110000011001",
			1740 => "0000000000000000001100110000000100",
			1741 => "11111111011101010001110000011001",
			1742 => "00000001000101000001110000011001",
			1743 => "0000001000000000001111000101101000",
			1744 => "0000000110000000000100111100110100",
			1745 => "0000001000000000001010110000011000",
			1746 => "0000000100000000001111100100001100",
			1747 => "0000001011000000000101100100001000",
			1748 => "0000001110000000000111011000000100",
			1749 => "00000000111101010001110000011001",
			1750 => "11111110101111100001110000011001",
			1751 => "11111110100111110001110000011001",
			1752 => "0000001100000000001001110100001000",
			1753 => "0000001100000000000100011000000100",
			1754 => "00000000000001010001110000011001",
			1755 => "00000010001100010001110000011001",
			1756 => "11111111001111110001110000011001",
			1757 => "0000001100000000001000111100001100",
			1758 => "0000000110000000001101011000000100",
			1759 => "11111110100100100001110000011001",
			1760 => "0000001111000000000010000000000100",
			1761 => "00000000100101010001110000011001",
			1762 => "11111110011011000001110000011001",
			1763 => "0000000100000000001000000100001000",
			1764 => "0000001000000000001001101000000100",
			1765 => "00000000010101010001110000011001",
			1766 => "11111110011101100001110000011001",
			1767 => "0000001001000000001001111100000100",
			1768 => "11111111011011000001110000011001",
			1769 => "11111101111001010001110000011001",
			1770 => "0000001100000000001100110000011000",
			1771 => "0000001100000000000100000000001000",
			1772 => "0000000101000000001001110100000100",
			1773 => "11111101111000010001110000011001",
			1774 => "00000000111001000001110000011001",
			1775 => "0000001001000000001010011000001000",
			1776 => "0000000010000000001111010100000100",
			1777 => "00000000110110110001110000011001",
			1778 => "00000001111011010001110000011001",
			1779 => "0000001100000000000011011100000100",
			1780 => "00000000000000000001110000011001",
			1781 => "00000001001101110001110000011001",
			1782 => "0000001001000000001100011000001100",
			1783 => "0000000001000000001011101000000100",
			1784 => "11111101110101110001110000011001",
			1785 => "0000000001000000001111001100000100",
			1786 => "00000001100101000001110000011001",
			1787 => "00000000000000000001110000011001",
			1788 => "0000001101000000000111111100001000",
			1789 => "0000000001000000001110010100000100",
			1790 => "00000000001110000001110000011001",
			1791 => "00000001100000010001110000011001",
			1792 => "0000001111000000001000110100000100",
			1793 => "11111111001110100001110000011001",
			1794 => "00000000100011010001110000011001",
			1795 => "0000001100000000001000111100000100",
			1796 => "00000001010010010001110000011001",
			1797 => "11111110001001010001110000011001",
			1798 => "0000000110000000001101011001001100",
			1799 => "0000001001000000001000010000100100",
			1800 => "0000000001000000000110101000001100",
			1801 => "0000000011000000001010001100000100",
			1802 => "11111110011000010001110110101101",
			1803 => "0000000011000000000100000100000100",
			1804 => "00000001000010000001110110101101",
			1805 => "11111110100001100001110110101101",
			1806 => "0000001001000000001001011000000100",
			1807 => "00000010011100110001110110101101",
			1808 => "0000001101000000000010110100010000",
			1809 => "0000000001000000001101011100001000",
			1810 => "0000001110000000000010001000000100",
			1811 => "11111110010011100001110110101101",
			1812 => "00000000000000110001110110101101",
			1813 => "0000001011000000000011100000000100",
			1814 => "11111111100001110001110110101101",
			1815 => "00000101100010010001110110101101",
			1816 => "11111110011001100001110110101101",
			1817 => "0000000111000000001001001000001000",
			1818 => "0000001101000000001110101100000100",
			1819 => "00000001110011000001110110101101",
			1820 => "11111110011001100001110110101101",
			1821 => "0000000111000000000110100100010000",
			1822 => "0000001110000000000010000000000100",
			1823 => "11111110111101110001110110101101",
			1824 => "0000000001000000000001000100000100",
			1825 => "11111111010000010001110110101101",
			1826 => "0000001000000000001001000100000100",
			1827 => "00000101001001100001110110101101",
			1828 => "00000010010010110001110110101101",
			1829 => "0000000000000000001001101000001000",
			1830 => "0000001011000000000101100100000100",
			1831 => "00000001010111010001110110101101",
			1832 => "11111110011110110001110110101101",
			1833 => "0000001100000000001001110100000100",
			1834 => "00000011000011100001110110101101",
			1835 => "11111110101011000001110110101101",
			1836 => "0000001100000000001000011001011000",
			1837 => "0000000110000000001000010000110100",
			1838 => "0000001100000000001000111100010100",
			1839 => "0000001011000000000011011100001000",
			1840 => "0000000100000000000110110000000100",
			1841 => "11111110010101000001110110101101",
			1842 => "00000000110000100001110110101101",
			1843 => "0000000001000000000111100100001000",
			1844 => "0000001111000000001110010000000100",
			1845 => "00000001100101110001110110101101",
			1846 => "00000000000111100001110110101101",
			1847 => "00000010000011110001110110101101",
			1848 => "0000001000000000001001101000010000",
			1849 => "0000001000000000000001110000001000",
			1850 => "0000001011000000000110110100000100",
			1851 => "00000000101110100001110110101101",
			1852 => "11111111001011010001110110101101",
			1853 => "0000000110000000001001100100000100",
			1854 => "11111111010111100001110110101101",
			1855 => "00000001111010000001110110101101",
			1856 => "0000000111000000000101101100001000",
			1857 => "0000000011000000001011011100000100",
			1858 => "11111110111000010001110110101101",
			1859 => "00000001100010010001110110101101",
			1860 => "0000001010000000000110011100000100",
			1861 => "11111110000100100001110110101101",
			1862 => "11111111100101010001110110101101",
			1863 => "0000001011000000001011110100010100",
			1864 => "0000000100000000000011010100001100",
			1865 => "0000000011000000001100010100000100",
			1866 => "00000001000101110001110110101101",
			1867 => "0000001010000000001001000100000100",
			1868 => "00000001000010110001110110101101",
			1869 => "00000001111100000001110110101101",
			1870 => "0000001100000000000110000100000100",
			1871 => "00000001111110010001110110101101",
			1872 => "11111110111001110001110110101101",
			1873 => "0000001110000000001011110000000100",
			1874 => "11111110000010000001110110101101",
			1875 => "0000001100000000001001110100000100",
			1876 => "11111110110011100001110110101101",
			1877 => "0000000110000000000101010000000100",
			1878 => "11111110111011100001110110101101",
			1879 => "00000010011100110001110110101101",
			1880 => "0000001001000000001000010100100000",
			1881 => "0000001010000000001010110000011100",
			1882 => "0000001101000000001010000100010000",
			1883 => "0000001001000000001001111100001000",
			1884 => "0000001101000000001100000000000100",
			1885 => "11111110111101100001110110101101",
			1886 => "00000011010001010001110110101101",
			1887 => "0000001011000000000110100000000100",
			1888 => "11111110100110010001110110101101",
			1889 => "11111111101010010001110110101101",
			1890 => "0000001000000000000001010100000100",
			1891 => "00000111100000100001110110101101",
			1892 => "0000001001000000001010100000000100",
			1893 => "00000011001011010001110110101101",
			1894 => "11111110100100010001110110101101",
			1895 => "11111110011001010001110110101101",
			1896 => "0000001111000000000000010100000100",
			1897 => "11111111000101000001110110101101",
			1898 => "00000001110011110001110110101101",
			1899 => "0000000100000000001011110001001100",
			1900 => "0000000110000000001001100100111100",
			1901 => "0000001100000000000100001000001100",
			1902 => "0000000010000000000010110100000100",
			1903 => "00000000000000000001111101011001",
			1904 => "0000001100000000000100000000000100",
			1905 => "00000000000000000001111101011001",
			1906 => "11111111000101100001111101011001",
			1907 => "0000001100000000000100011000011000",
			1908 => "0000001110000000001100000000001100",
			1909 => "0000000101000000001001010100001000",
			1910 => "0000000001000000001011111100000100",
			1911 => "00000000100000000001111101011001",
			1912 => "00000000000000000001111101011001",
			1913 => "11111111101100010001111101011001",
			1914 => "0000000101000000000111100000001000",
			1915 => "0000001011000000000000011100000100",
			1916 => "00000000000000000001111101011001",
			1917 => "00000000100111100001111101011001",
			1918 => "00000000000000000001111101011001",
			1919 => "0000001110000000001100000000001100",
			1920 => "0000001111000000001111010100000100",
			1921 => "11111111111011010001111101011001",
			1922 => "0000001111000000000111010100000100",
			1923 => "00000000100110110001111101011001",
			1924 => "00000000000000000001111101011001",
			1925 => "0000001010000000000010101100000100",
			1926 => "00000000000000000001111101011001",
			1927 => "0000000001000000001011111100000100",
			1928 => "00000000000000000001111101011001",
			1929 => "11111111010011110001111101011001",
			1930 => "0000001010000000000111110100000100",
			1931 => "00000000000000000001111101011001",
			1932 => "0000001110000000001100111000001000",
			1933 => "0000000111000000001111011100000100",
			1934 => "00000000111110100001111101011001",
			1935 => "00000000000000000001111101011001",
			1936 => "00000000000000000001111101011001",
			1937 => "0000000100000000001110111001000100",
			1938 => "0000000110000000000100111100011000",
			1939 => "0000000111000000001000111000001100",
			1940 => "0000001101000000001011000000001000",
			1941 => "0000001011000000000101101100000100",
			1942 => "11111111100011000001111101011001",
			1943 => "00000000000000000001111101011001",
			1944 => "00000000110011110001111101011001",
			1945 => "0000001011000000000001001000001000",
			1946 => "0000000010000000000110010000000100",
			1947 => "00000000000000000001111101011001",
			1948 => "11111111001111000001111101011001",
			1949 => "00000000000000000001111101011001",
			1950 => "0000000110000000001000010000010000",
			1951 => "0000000011000000001101000100000100",
			1952 => "00000000000000000001111101011001",
			1953 => "0000000100000000001100001100000100",
			1954 => "00000000000000000001111101011001",
			1955 => "0000000001000000001010011000000100",
			1956 => "00000000110101010001111101011001",
			1957 => "00000000000000000001111101011001",
			1958 => "0000001011000000000101110100010000",
			1959 => "0000000001000000000001000100001000",
			1960 => "0000001010000000001100011100000100",
			1961 => "11111111001110100001111101011001",
			1962 => "00000000000000000001111101011001",
			1963 => "0000001000000000000001110000000100",
			1964 => "00000000000000000001111101011001",
			1965 => "00000001000001000001111101011001",
			1966 => "0000000001000000001010011000001000",
			1967 => "0000001000000000001001101000000100",
			1968 => "11111110111000100001111101011001",
			1969 => "00000000000000000001111101011001",
			1970 => "00000000000000000001111101011001",
			1971 => "0000001110000000000110010000101000",
			1972 => "0000000001000000001001111000011000",
			1973 => "0000001100000000000100000000001100",
			1974 => "0000000101000000001010111100000100",
			1975 => "00000000000000000001111101011001",
			1976 => "0000001011000000000101101100000100",
			1977 => "00000001000000010001111101011001",
			1978 => "00000000000000000001111101011001",
			1979 => "0000000100000000000010010000001000",
			1980 => "0000000111000000000100000000000100",
			1981 => "00000000000000000001111101011001",
			1982 => "11111110111011100001111101011001",
			1983 => "00000000000000000001111101011001",
			1984 => "0000001000000000001111000100001100",
			1985 => "0000000110000000001001100100000100",
			1986 => "00000000000000000001111101011001",
			1987 => "0000000100000000000011111000000100",
			1988 => "00000001000011010001111101011001",
			1989 => "00000000000000000001111101011001",
			1990 => "00000000000000000001111101011001",
			1991 => "0000001110000000000010110000001100",
			1992 => "0000001101000000000111010100001000",
			1993 => "0000001100000000001000000000000100",
			1994 => "11111111111011100001111101011001",
			1995 => "11111110111000100001111101011001",
			1996 => "00000000000000000001111101011001",
			1997 => "0000001101000000001101101100001100",
			1998 => "0000000001000000001101111100000100",
			1999 => "00000000000000000001111101011001",
			2000 => "0000000001000000000100111100000100",
			2001 => "00000000101101110001111101011001",
			2002 => "00000000000000000001111101011001",
			2003 => "0000001100000000000101110100000100",
			2004 => "11111111101010110001111101011001",
			2005 => "00000000000000000001111101011001",
			2006 => "0000000110000000001101011000101000",
			2007 => "0000000001000000000001000100010100",
			2008 => "0000001000000000001001000100010000",
			2009 => "0000000000000000000001110000000100",
			2010 => "11111110011101010010000011000101",
			2011 => "0000000001000000001101011100001000",
			2012 => "0000001001000000000010001100000100",
			2013 => "00000000000000000010000011000101",
			2014 => "00000010000111110010000011000101",
			2015 => "11111110111101000010000011000101",
			2016 => "11111110011001010010000011000101",
			2017 => "0000000011000000001010000100010000",
			2018 => "0000001101000000000010011100001100",
			2019 => "0000001001000000000100101100001000",
			2020 => "0000001011000000000101100100000100",
			2021 => "11111110100100110010000011000101",
			2022 => "00000000101000110010000011000101",
			2023 => "00000010011011100010000011000101",
			2024 => "00000100000000110010000011000101",
			2025 => "11111110110100010010000011000101",
			2026 => "0000000101000000000111111101100000",
			2027 => "0000000110000000001000010000110100",
			2028 => "0000000100000000001110000000011000",
			2029 => "0000000001000000000111100100001000",
			2030 => "0000001011000000001100101100000100",
			2031 => "00000000000100100010000011000101",
			2032 => "11111110000100000010000011000101",
			2033 => "0000000000000000000001110100001000",
			2034 => "0000001010000000000011101000000100",
			2035 => "00000001001110100010000011000101",
			2036 => "11111111011110010010000011000101",
			2037 => "0000000110000000001001100100000100",
			2038 => "11111111111010110010000011000101",
			2039 => "00000001101001100010000011000101",
			2040 => "0000001011000000001100101100001100",
			2041 => "0000001011000000000011011100000100",
			2042 => "11111110011000100010000011000101",
			2043 => "0000000111000000001000111000000100",
			2044 => "00000001010101100010000011000101",
			2045 => "00000000001101100010000011000101",
			2046 => "0000001000000000001111001000001000",
			2047 => "0000001010000000001010110000000100",
			2048 => "11111111010111110010000011000101",
			2049 => "00000001100111000010000011000101",
			2050 => "0000001001000000001100011000000100",
			2051 => "11111101111011110010000011000101",
			2052 => "00000000110101100010000011000101",
			2053 => "0000000100000000000100001100011000",
			2054 => "0000000000000000001010101100001000",
			2055 => "0000001011000000000010001000000100",
			2056 => "11111101111110010010000011000101",
			2057 => "00000001101001000010000011000101",
			2058 => "0000000111000000001111011100001000",
			2059 => "0000000001000000001011101000000100",
			2060 => "00000000111011010010000011000101",
			2061 => "00000001101000100010000011000101",
			2062 => "0000001111000000001000110100000100",
			2063 => "11111110010000000010000011000101",
			2064 => "00000001101001000010000011000101",
			2065 => "0000000001000000000111100100001000",
			2066 => "0000000110000000001000010000000100",
			2067 => "00000010001100100010000011000101",
			2068 => "00000001001001100010000011000101",
			2069 => "0000000100000000001100111100001000",
			2070 => "0000001100000000001000000000000100",
			2071 => "00000000001110010010000011000101",
			2072 => "11111110010011100010000011000101",
			2073 => "11111101110110100010000011000101",
			2074 => "0000000000000000001011000100101100",
			2075 => "0000001101000000001111010100011100",
			2076 => "0000001001000000000100101100001100",
			2077 => "0000001100000000001111011100001000",
			2078 => "0000001101000000001100000000000100",
			2079 => "00000000011000010010000011000101",
			2080 => "00000001111001000010000011000101",
			2081 => "11111111000010000010000011000101",
			2082 => "0000001101000000000110111100001000",
			2083 => "0000001111000000001010110100000100",
			2084 => "11111110100011110010000011000101",
			2085 => "00000001011011100010000011000101",
			2086 => "0000001010000000001000010100000100",
			2087 => "00000100000110110010000011000101",
			2088 => "11111110110010000010000011000101",
			2089 => "0000000000000000000111000000000100",
			2090 => "00000011001111000010000011000101",
			2091 => "0000001001000000000111101100000100",
			2092 => "00000010100001000010000011000101",
			2093 => "0000000110000000001001111100000100",
			2094 => "11111110100010000010000011000101",
			2095 => "00000000101001000010000011000101",
			2096 => "11111110010100110010000011000101",
			2097 => "0000001001000000000111101110000100",
			2098 => "0000001000000000001011010101000100",
			2099 => "0000001010000000001000010100100100",
			2100 => "0000001100000000000100011000010000",
			2101 => "0000001101000000001111010000001100",
			2102 => "0000001100000000000110000100000100",
			2103 => "11111111011011000010001001011001",
			2104 => "0000000001000000001011101000000100",
			2105 => "00000000111011010010001001011001",
			2106 => "11111111111000110010001001011001",
			2107 => "11111110101111010010001001011001",
			2108 => "0000000000000000001111001000001100",
			2109 => "0000000111000000000001101000000100",
			2110 => "11111111011111010010001001011001",
			2111 => "0000001100000000001001110100000100",
			2112 => "00000000011101010010001001011001",
			2113 => "11111111100111110010001001011001",
			2114 => "0000000011000000001010000100000100",
			2115 => "00000000111011110010001001011001",
			2116 => "00000000000000000010001001011001",
			2117 => "0000000100000000000110111000001100",
			2118 => "0000001011000000001101111000001000",
			2119 => "0000000001000000000111100100000100",
			2120 => "00000000000000000010001001011001",
			2121 => "00000000110101110010001001011001",
			2122 => "11111111100011100010001001011001",
			2123 => "0000000011000000001111101000001100",
			2124 => "0000000111000000001000111000000100",
			2125 => "00000000000000000010001001011001",
			2126 => "0000001100000000000000101000000100",
			2127 => "00000000000000000010001001011001",
			2128 => "11111110010010110010001001011001",
			2129 => "0000001110000000001111101000000100",
			2130 => "00000000000101000010001001011001",
			2131 => "00000000000000000010001001011001",
			2132 => "0000000001000000001011101000100100",
			2133 => "0000001100000000001100110000100000",
			2134 => "0000000011000000001010011100010000",
			2135 => "0000000111000000001000111000001000",
			2136 => "0000000110000000001001100100000100",
			2137 => "11111111101100100010001001011001",
			2138 => "00000000110110110010001001011001",
			2139 => "0000000100000000000010010000000100",
			2140 => "11111110110011000010001001011001",
			2141 => "00000000000000000010001001011001",
			2142 => "0000001110000000000110100100001000",
			2143 => "0000000111000000001101100000000100",
			2144 => "00000001001110010010001001011001",
			2145 => "00000000000000000010001001011001",
			2146 => "0000000011000000000101110100000100",
			2147 => "11111111101111010010001001011001",
			2148 => "00000000001111000010001001011001",
			2149 => "11111110101001100010001001011001",
			2150 => "0000000101000000001010010100001100",
			2151 => "0000000100000000000000100000001000",
			2152 => "0000000110000000001000010000000100",
			2153 => "00000000000000000010001001011001",
			2154 => "00000001100101000010001001011001",
			2155 => "00000000000000000010001001011001",
			2156 => "0000000101000000000111100000000100",
			2157 => "11111110111100010010001001011001",
			2158 => "0000000100000000000011110100000100",
			2159 => "00000000000000000010001001011001",
			2160 => "0000001010000000000110011100000100",
			2161 => "00000001000111110010001001011001",
			2162 => "00000000000000000010001001011001",
			2163 => "0000001001000000001010100000100100",
			2164 => "0000001110000000001100010000000100",
			2165 => "11111111011011000010001001011001",
			2166 => "0000000100000000000100001100011000",
			2167 => "0000000000000000000111000100001100",
			2168 => "0000001010000000000011101000001000",
			2169 => "0000000111000000000001101000000100",
			2170 => "00000000100001100010001001011001",
			2171 => "00000000000000000010001001011001",
			2172 => "11111111100101010010001001011001",
			2173 => "0000001010000000000111110100000100",
			2174 => "00000000000000000010001001011001",
			2175 => "0000000111000000001000011000000100",
			2176 => "00000001010010110010001001011001",
			2177 => "00000000000100110010001001011001",
			2178 => "0000001010000000001010110000000100",
			2179 => "00000000000000000010001001011001",
			2180 => "11111111011101110010001001011001",
			2181 => "0000001110000000000011010100100000",
			2182 => "0000001011000000001101000100011100",
			2183 => "0000000001000000000100110100001100",
			2184 => "0000001110000000001000110100001000",
			2185 => "0000001101000000000101110000000100",
			2186 => "00000000000000000010001001011001",
			2187 => "11111111001001100010001001011001",
			2188 => "00000000000000000010001001011001",
			2189 => "0000000001000000001100011000001000",
			2190 => "0000001000000000000101000100000100",
			2191 => "00000000000000000010001001011001",
			2192 => "00000001000101000010001001011001",
			2193 => "0000001011000000000110100000000100",
			2194 => "11111111110010110010001001011001",
			2195 => "00000000110001110010001001011001",
			2196 => "11111110101001110010001001011001",
			2197 => "00000000101110110010001001011001",
			2198 => "0000001000000000001001000100011100",
			2199 => "0000000111000000000001101000011000",
			2200 => "0000001100000000001110001100000100",
			2201 => "00000000000000000010001111000101",
			2202 => "0000001011000000001011011100010000",
			2203 => "0000001000000000000010101100000100",
			2204 => "00000000000000000010001111000101",
			2205 => "0000001101000000000101110000001000",
			2206 => "0000000101000000000111100000000100",
			2207 => "00000000111100100010001111000101",
			2208 => "00000000000000000010001111000101",
			2209 => "00000000000000000010001111000101",
			2210 => "00000000000000000010001111000101",
			2211 => "00000000000000000010001111000101",
			2212 => "0000000000000000000011010001010000",
			2213 => "0000000001000000000111100100100100",
			2214 => "0000000111000000001101100000011000",
			2215 => "0000000101000000000100011000010000",
			2216 => "0000001011000000000101101100001000",
			2217 => "0000000100000000000010110000000100",
			2218 => "11111111001101110010001111000101",
			2219 => "00000000000000000010001111000101",
			2220 => "0000000111000000001001110000000100",
			2221 => "00000000010101010010001111000101",
			2222 => "00000000000000000010001111000101",
			2223 => "0000001100000000001100001000000100",
			2224 => "00000000000000000010001111000101",
			2225 => "11111110101000100010001111000101",
			2226 => "0000001100000000000100000000000100",
			2227 => "00000000010110100010001111000101",
			2228 => "0000001111000000000010011100000100",
			2229 => "00000000000000000010001111000101",
			2230 => "11111111110000000010001111000101",
			2231 => "0000001101000000000101100100010000",
			2232 => "0000001111000000000010000100001100",
			2233 => "0000000001000000000111100100000100",
			2234 => "00000000000000000010001111000101",
			2235 => "0000000000000000001000101100000100",
			2236 => "00000000000000000010001111000101",
			2237 => "00000001001000110010001111000101",
			2238 => "00000000000000000010001111000101",
			2239 => "0000000001000000001001011000001100",
			2240 => "0000000001000000001011101000000100",
			2241 => "00000000000000000010001111000101",
			2242 => "0000001011000000001010111000000100",
			2243 => "00000000000000000010001111000101",
			2244 => "11111110100111110010001111000101",
			2245 => "0000001001000000000101010000001000",
			2246 => "0000000000000000001101010000000100",
			2247 => "00000000111011110010001111000101",
			2248 => "00000000000000000010001111000101",
			2249 => "0000001010000000001001000100000100",
			2250 => "11111111110010100010001111000101",
			2251 => "00000000001100100010001111000101",
			2252 => "0000001100000000001100110000101000",
			2253 => "0000000011000000000101110100011100",
			2254 => "0000000010000000001110110100001100",
			2255 => "0000000011000000001010011100001000",
			2256 => "0000000100000000001110111000000100",
			2257 => "11111111010101100010001111000101",
			2258 => "00000000000000000010001111000101",
			2259 => "00000001010100110010001111000101",
			2260 => "0000000000000000000000111000001000",
			2261 => "0000000000000000000011010000000100",
			2262 => "00000000000000000010001111000101",
			2263 => "11111110110011110010001111000101",
			2264 => "0000000011000000000000011100000100",
			2265 => "11111111110100000010001111000101",
			2266 => "00000000100101100010001111000101",
			2267 => "0000001111000000001111100100001000",
			2268 => "0000001000000000001111001000000100",
			2269 => "00000000000000000010001111000101",
			2270 => "00000001010100010010001111000101",
			2271 => "00000000000000000010001111000101",
			2272 => "0000000000000000000000111000001100",
			2273 => "0000001100000000001000011000001000",
			2274 => "0000001000000000000110001000000100",
			2275 => "00000000000000000010001111000101",
			2276 => "00000000110110000010001111000101",
			2277 => "00000000000000000010001111000101",
			2278 => "0000000011000000000011011000010000",
			2279 => "0000001000000000000111000100001000",
			2280 => "0000001000000000000111000100000100",
			2281 => "11111111110000000010001111000101",
			2282 => "00000000001110000010001111000101",
			2283 => "0000000100000000001011100000000100",
			2284 => "00000000000000000010001111000101",
			2285 => "11111110101111110010001111000101",
			2286 => "0000001000000000001110111100000100",
			2287 => "00000000100010000010001111000101",
			2288 => "00000000000000000010001111000101",
			2289 => "0000000101000000001010111100001000",
			2290 => "0000001000000000000000101000000100",
			2291 => "11111110110110000010010011011001",
			2292 => "00000000000000000010010011011001",
			2293 => "0000001100000000000100000000011000",
			2294 => "0000000100000000000010111000001000",
			2295 => "0000001001000000000101011100000100",
			2296 => "11111111001000010010010011011001",
			2297 => "00000000011000010010010011011001",
			2298 => "0000000101000000001010111100000100",
			2299 => "00000000000000000010010011011001",
			2300 => "0000000110000000001011001100001000",
			2301 => "0000000110000000001101011000000100",
			2302 => "00000000000000000010010011011001",
			2303 => "00000000000101010010010011011001",
			2304 => "00000001100010100010010011011001",
			2305 => "0000000011000000000010000100111000",
			2306 => "0000001000000000000110001000100000",
			2307 => "0000000100000000000011000000010000",
			2308 => "0000000110000000001001100100001000",
			2309 => "0000001100000000000110000100000100",
			2310 => "11111111001101110010010011011001",
			2311 => "00000000001000110010010011011001",
			2312 => "0000000010000000001100010000000100",
			2313 => "00000000101111000010010011011001",
			2314 => "00000000000000000010010011011001",
			2315 => "0000001111000000000101110000001000",
			2316 => "0000000111000000001001110000000100",
			2317 => "00000000011111100010010011011001",
			2318 => "11111111010001010010010011011001",
			2319 => "0000001100000000000100000000000100",
			2320 => "00000000000000000010010011011001",
			2321 => "11111110100010100010010011011001",
			2322 => "0000001100000000000100000000001100",
			2323 => "0000001000000000001111001000000100",
			2324 => "00000000000000000010010011011001",
			2325 => "0000000011000000000110100100000100",
			2326 => "00000000000000000010010011011001",
			2327 => "11111110011110100010010011011001",
			2328 => "0000001100000000001100110000001000",
			2329 => "0000000011000000001000011000000100",
			2330 => "11111111100010110010010011011001",
			2331 => "00000000010111000010010011011001",
			2332 => "11111110110100000010010011011001",
			2333 => "0000000101000000000001000000010100",
			2334 => "0000001000000000000111000000010000",
			2335 => "0000000010000000001000101000001000",
			2336 => "0000001001000000001010100000000100",
			2337 => "00000000100100100010010011011001",
			2338 => "11111111100011100010010011011001",
			2339 => "0000001111000000001000101000000100",
			2340 => "00000000000000000010010011011001",
			2341 => "00000001010111010010010011011001",
			2342 => "11111111101111010010010011011001",
			2343 => "0000000101000000001001010000010000",
			2344 => "0000000001000000000100110100001000",
			2345 => "0000000011000000000110111000000100",
			2346 => "11111110000110110010010011011001",
			2347 => "00000000000000000010010011011001",
			2348 => "0000000101000000000101001000000100",
			2349 => "00000000100000110010010011011001",
			2350 => "00000000000000000010010011011001",
			2351 => "0000001100000000000001011000001000",
			2352 => "0000000100000000000011101100000100",
			2353 => "00000000000100000010010011011001",
			2354 => "00000000111101100010010011011001",
			2355 => "0000000101000000001111100100000100",
			2356 => "11111110101101100010010011011001",
			2357 => "00000000000000000010010011011001",
			2358 => "0000001101000000001010111100001000",
			2359 => "0000000010000000000000010000000100",
			2360 => "11111110100101110010011000000101",
			2361 => "00000000000000000010011000000101",
			2362 => "0000001111000000000010011101001000",
			2363 => "0000000011000000000000011100110000",
			2364 => "0000000100000000001001001100010100",
			2365 => "0000000111000000000100000000001000",
			2366 => "0000001011000000000101101100000100",
			2367 => "11111111101000010010011000000101",
			2368 => "00000000010110010010011000000101",
			2369 => "0000001111000000001100100100001000",
			2370 => "0000001101000000000011100000000100",
			2371 => "11111111010001000010011000000101",
			2372 => "00000000000011000010011000000101",
			2373 => "11111110011110100010011000000101",
			2374 => "0000000010000000001100010000001100",
			2375 => "0000000110000000001101011000000100",
			2376 => "00000000000000000010011000000101",
			2377 => "0000001100000000001000111000000100",
			2378 => "00000001100001100010011000000101",
			2379 => "00000000000000000010011000000101",
			2380 => "0000000110000000001111000000001000",
			2381 => "0000000111000000001000111000000100",
			2382 => "00000000000000000010011000000101",
			2383 => "11111110100100100010011000000101",
			2384 => "0000001100000000001000111000000100",
			2385 => "00000001000010000010011000000101",
			2386 => "11111111010100000010011000000101",
			2387 => "0000001010000000001000010100010000",
			2388 => "0000000010000000001110000100001100",
			2389 => "0000000111000000000001111100000100",
			2390 => "00000000000000000010011000000101",
			2391 => "0000001011000000001011000000000100",
			2392 => "00000000110100000010011000000101",
			2393 => "00000000000000000010011000000101",
			2394 => "11111111001101000010011000000101",
			2395 => "0000000100000000000000101100000100",
			2396 => "00000001100100100010011000000101",
			2397 => "00000000000000000010011000000101",
			2398 => "0000000011000000001011011100001100",
			2399 => "0000000110000000001111000000000100",
			2400 => "11111101111101000010011000000101",
			2401 => "0000001111000000001001011100000100",
			2402 => "00000001001100110010011000000101",
			2403 => "00000000000000000010011000000101",
			2404 => "0000001100000000000110100100100000",
			2405 => "0000001011000000000101110100010000",
			2406 => "0000000110000000001000010000001000",
			2407 => "0000000010000000001111010100000100",
			2408 => "00000000010001100010011000000101",
			2409 => "11111111100111000010011000000101",
			2410 => "0000000100000000001001000000000100",
			2411 => "00000001011010000010011000000101",
			2412 => "11111111010100000010011000000101",
			2413 => "0000001101000000001100010100001000",
			2414 => "0000001001000000001010100000000100",
			2415 => "11111100010110000010011000000101",
			2416 => "00000000000000000010011000000101",
			2417 => "0000001101000000001110110100000100",
			2418 => "00000000100100110010011000000101",
			2419 => "11111110101001110010011000000101",
			2420 => "0000000110000000001001111100001100",
			2421 => "0000000100000000001011110000000100",
			2422 => "11111111001001010010011000000101",
			2423 => "0000000001000000001100011000000100",
			2424 => "00000001000111100010011000000101",
			2425 => "00000000001010010010011000000101",
			2426 => "0000001110000000000011010100001000",
			2427 => "0000001011000000001001011100000100",
			2428 => "11111110101000100010011000000101",
			2429 => "00000000000000000010011000000101",
			2430 => "0000001101000000001100111000000100",
			2431 => "00000001000000100010011000000101",
			2432 => "00000000000000000010011000000101",
			2433 => "0000000110000000001001100101100000",
			2434 => "0000001111000000000000010001010100",
			2435 => "0000000110000000001011001100100100",
			2436 => "0000001001000000000101010000010100",
			2437 => "0000000110000000001101011000001100",
			2438 => "0000000001000000000110101000000100",
			2439 => "11010001011011100010011111000001",
			2440 => "0000001001000000001001011000000100",
			2441 => "11010101000111110010011111000001",
			2442 => "11010001100001000010011111000001",
			2443 => "0000000011000000000100000100000100",
			2444 => "11010001100111010010011111000001",
			2445 => "11010011001000100010011111000001",
			2446 => "0000001010000000000010101100001100",
			2447 => "0000001011000000001011011100001000",
			2448 => "0000000010000000001100000000000100",
			2449 => "11010011010010000010011111000001",
			2450 => "11100011011010000010011111000001",
			2451 => "11010001100101110010011111000001",
			2452 => "11010001011101100010011111000001",
			2453 => "0000001100000000000100000000011000",
			2454 => "0000001101000000000011100000001100",
			2455 => "0000000101000000000111001000000100",
			2456 => "11010001011110100010011111000001",
			2457 => "0000000001000000001001111000000100",
			2458 => "11011011101001110010011111000001",
			2459 => "11010001101110000010011111000001",
			2460 => "0000000010000000001100010000001000",
			2461 => "0000000011000000000000011100000100",
			2462 => "11100000110100100010011111000001",
			2463 => "11101011010111010010011111000001",
			2464 => "11010001101010010010011111000001",
			2465 => "0000001010000000000010101100001000",
			2466 => "0000001100000000000100011000000100",
			2467 => "11011001000100010010011111000001",
			2468 => "11010001110101000010011111000001",
			2469 => "0000001100000000001011000000001000",
			2470 => "0000000010000000001001010000000100",
			2471 => "11010011101100000010011111000001",
			2472 => "11010001100101010010011111000001",
			2473 => "0000000011000000001111010100000100",
			2474 => "11011000011011000010011111000001",
			2475 => "11010001100101100010011111000001",
			2476 => "0000001100000000000100011000000100",
			2477 => "11011110000110010010011111000001",
			2478 => "0000000100000000001000101000000100",
			2479 => "11010001100001000010011111000001",
			2480 => "11010111111000010010011111000001",
			2481 => "0000001100000000001001110101010100",
			2482 => "0000000110000000000100111100101100",
			2483 => "0000000010000000001111010100011000",
			2484 => "0000001100000000001001110000001100",
			2485 => "0000000101000000001010111100000100",
			2486 => "11010011101100000010011111000001",
			2487 => "0000000110000000001001100100000100",
			2488 => "11100101000100000010011111000001",
			2489 => "11101011011100000010011111000001",
			2490 => "0000000001000000000111100100001000",
			2491 => "0000000001000000000111100100000100",
			2492 => "11010011111001010010011111000001",
			2493 => "11010001110101000010011111000001",
			2494 => "11011001000100010010011111000001",
			2495 => "0000001011000000001100101100000100",
			2496 => "11011100001111110010011111000001",
			2497 => "0000001111000000001011101100001000",
			2498 => "0000000100000000000011000000000100",
			2499 => "11010010111101010010011111000001",
			2500 => "11010001011111100010011111000001",
			2501 => "0000001000000000000101000100000100",
			2502 => "11010011001000100010011111000001",
			2503 => "11100101111111100010011111000001",
			2504 => "0000000101000000000010011100011100",
			2505 => "0000001000000000000001010100001100",
			2506 => "0000001011000000001011011100000100",
			2507 => "11100010000001000010011111000001",
			2508 => "0000001101000000000100101000000100",
			2509 => "11010110011110110010011111000001",
			2510 => "11010001101011000010011111000001",
			2511 => "0000000100000000001001000000001000",
			2512 => "0000000110000000001000010000000100",
			2513 => "11100110111010010010011111000001",
			2514 => "11101100101111100010011111000001",
			2515 => "0000001100000000001100110000000100",
			2516 => "11100110000110000010011111000001",
			2517 => "11010010101111000010011111000001",
			2518 => "0000000010000000000011110000001000",
			2519 => "0000000110000000001000010000000100",
			2520 => "11010111011010100010011111000001",
			2521 => "11010001101101000010011111000001",
			2522 => "11011111100001010010011111000001",
			2523 => "0000001100000000000001101000010000",
			2524 => "0000000110000000000101010000001100",
			2525 => "0000000110000000000100111100001000",
			2526 => "0000000001000000001100011000000100",
			2527 => "11011001000100010010011111000001",
			2528 => "11010001101110000010011111000001",
			2529 => "11010001100000110010011111000001",
			2530 => "11100001010010100010011111000001",
			2531 => "0000001001000000001000010100010100",
			2532 => "0000001101000000001100010100000100",
			2533 => "11010111111000010010011111000001",
			2534 => "0000000110000000001111000000001000",
			2535 => "0000000001000000001100011000000100",
			2536 => "11010110011110110010011111000001",
			2537 => "11010001110101000010011111000001",
			2538 => "0000001011000000000001001000000100",
			2539 => "11010010111000000010011111000001",
			2540 => "11010001100000100010011111000001",
			2541 => "0000000011000000001110111000000100",
			2542 => "11010001101110000010011111000001",
			2543 => "11011110001111000010011111000001",
			2544 => "0000000010000000001110000010100000",
			2545 => "0000000010000000000110111101000000",
			2546 => "0000000011000000000001101000010100",
			2547 => "0000001010000000000001010100001000",
			2548 => "0000000001000000000111100100000100",
			2549 => "11111110110011110010100110000101",
			2550 => "00000000000000000010100110000101",
			2551 => "0000001000000000001111000100001000",
			2552 => "0000000101000000001010111100000100",
			2553 => "00000000000000000010100110000101",
			2554 => "00000000110010010010100110000101",
			2555 => "11111111100010110010100110000101",
			2556 => "0000000000000000001111000100011000",
			2557 => "0000000001000000000111100100001000",
			2558 => "0000000010000000001100010100000100",
			2559 => "00000000000000000010100110000101",
			2560 => "11111110011000010010100110000101",
			2561 => "0000000101000000000100000100001000",
			2562 => "0000000001000000001101101000000100",
			2563 => "00000000000000000010100110000101",
			2564 => "00000000111101010010100110000101",
			2565 => "0000001100000000000100011000000100",
			2566 => "11111111000111010010100110000101",
			2567 => "00000000001100000010100110000101",
			2568 => "0000001110000000000010001000010000",
			2569 => "0000000010000000000010000100001000",
			2570 => "0000001100000000001000111000000100",
			2571 => "00000000111111000010100110000101",
			2572 => "11111110110111110010100110000101",
			2573 => "0000000110000000001111000000000100",
			2574 => "11111111000110000010100110000101",
			2575 => "00000000110000010010100110000101",
			2576 => "00000001011111110010100110000101",
			2577 => "0000000001000000000001111000111000",
			2578 => "0000000000000000000000111000011100",
			2579 => "0000000100000000001100001100010000",
			2580 => "0000000010000000000000010000001000",
			2581 => "0000000101000000000001101000000100",
			2582 => "00000000000000000010100110000101",
			2583 => "11111110111110110010100110000101",
			2584 => "0000001110000000001111100100000100",
			2585 => "00000000101001110010100110000101",
			2586 => "11111111100000010010100110000101",
			2587 => "0000001011000000001101111000000100",
			2588 => "00000000000000000010100110000101",
			2589 => "0000001010000000001100011100000100",
			2590 => "11111110001100010010100110000101",
			2591 => "00000000000000000010100110000101",
			2592 => "0000000110000000000100111100001100",
			2593 => "0000000010000000001111010100001000",
			2594 => "0000001100000000000100000000000100",
			2595 => "00000000100010010010100110000101",
			2596 => "11111111110000100010100110000101",
			2597 => "11111110100101010010100110000101",
			2598 => "0000000111000000000110000100001000",
			2599 => "0000000010000000001010000100000100",
			2600 => "00000000000000000010100110000101",
			2601 => "00000001011000110010100110000101",
			2602 => "0000000011000000001001011100000100",
			2603 => "11111110100111010010100110000101",
			2604 => "00000000101001000010100110000101",
			2605 => "0000001100000000001010111000001100",
			2606 => "0000001110000000001100010000000100",
			2607 => "00000000000000000010100110000101",
			2608 => "0000000001000000000100110100000100",
			2609 => "00000001010000100010100110000101",
			2610 => "00000000000000000010100110000101",
			2611 => "0000000000000000001010101100001100",
			2612 => "0000001110000000001100111000001000",
			2613 => "0000001000000000000101000100000100",
			2614 => "11111111100001100010100110000101",
			2615 => "00000000010000000010100110000101",
			2616 => "11111111000000100010100110000101",
			2617 => "0000001011000000000100010000001000",
			2618 => "0000001000000000000001010100000100",
			2619 => "00000000000000000010100110000101",
			2620 => "00000001000111000010100110000101",
			2621 => "0000001011000000000001001000000100",
			2622 => "11111111001100000010100110000101",
			2623 => "00000000101100110010100110000101",
			2624 => "0000001010000000000110011100101100",
			2625 => "0000001011000000000100010000001000",
			2626 => "0000000101000000000010110100000100",
			2627 => "00000000000000000010100110000101",
			2628 => "00000001010011000010100110000101",
			2629 => "0000000100000000000010100100011100",
			2630 => "0000001011000000000110100000010000",
			2631 => "0000000101000000000111111100001000",
			2632 => "0000000010000000000101000000000100",
			2633 => "11111111101101100010100110000101",
			2634 => "00000000011110110010100110000101",
			2635 => "0000000111000000000101110100000100",
			2636 => "11111110110001100010100110000101",
			2637 => "00000000000000000010100110000101",
			2638 => "0000001000000000001001101000001000",
			2639 => "0000000011000000001100001100000100",
			2640 => "00000000000000000010100110000101",
			2641 => "00000000111001110010100110000101",
			2642 => "00000000000000000010100110000101",
			2643 => "0000000000000000000000111000000100",
			2644 => "00000001001100110010100110000101",
			2645 => "00000000000000000010100110000101",
			2646 => "0000001010000000000101000100000100",
			2647 => "11111110101111100010100110000101",
			2648 => "0000001100000000000101100100010000",
			2649 => "0000000101000000000010011100001000",
			2650 => "0000001011000000000001101000000100",
			2651 => "00000000011101010010100110000101",
			2652 => "11111110111101100010100110000101",
			2653 => "0000000001000000000100110100000100",
			2654 => "00000000000000000010100110000101",
			2655 => "00000001010011100010100110000101",
			2656 => "11111111001000000010100110000101",
			2657 => "0000000011000000001011000000010000",
			2658 => "0000000110000000001001100100000100",
			2659 => "11111110011001100010101011111011",
			2660 => "0000000100000000000001001100000100",
			2661 => "11111111011101110010101011111011",
			2662 => "0000000010000000001111100100000100",
			2663 => "00000010000111100010101011111011",
			2664 => "11111111000010000010101011111011",
			2665 => "0000000110000000000100111101100000",
			2666 => "0000001100000000001000111100100100",
			2667 => "0000000110000000001101011000000100",
			2668 => "11111110100001100010101011111011",
			2669 => "0000000010000000000010000100010000",
			2670 => "0000000010000000001100010100001000",
			2671 => "0000001110000000000110100100000100",
			2672 => "00000001110010010010101011111011",
			2673 => "11111110100000000010101011111011",
			2674 => "0000000101000000000111001000000100",
			2675 => "11111111110000100010101011111011",
			2676 => "00000001111011000010101011111011",
			2677 => "0000000110000000001001100100001000",
			2678 => "0000001011000000000110000100000100",
			2679 => "11111111110001100010101011111011",
			2680 => "11111100110011100010101011111011",
			2681 => "0000000001000000000110101000000100",
			2682 => "00000000010000100010101011111011",
			2683 => "00000001110000010010101011111011",
			2684 => "0000000100000000001111101000011100",
			2685 => "0000000110000000001100011000001100",
			2686 => "0000001001000000000101011100001000",
			2687 => "0000001100000000001100110000000100",
			2688 => "11111111110011000010101011111011",
			2689 => "00000001010010010010101011111011",
			2690 => "11111110011111110010101011111011",
			2691 => "0000000110000000001101011000001000",
			2692 => "0000001100000000000100011000000100",
			2693 => "00000000110001010010101011111011",
			2694 => "00000010011000100010101011111011",
			2695 => "0000000000000000001111001000000100",
			2696 => "11111111101010000010101011111011",
			2697 => "00000001001110110010101011111011",
			2698 => "0000001011000000001110001100010000",
			2699 => "0000000011000000000001011000001000",
			2700 => "0000001111000000001001010000000100",
			2701 => "11111111110000000010101011111011",
			2702 => "11111101110101010010101011111011",
			2703 => "0000001111000000001110010000000100",
			2704 => "00000001111110000010101011111011",
			2705 => "11111111101010100010101011111011",
			2706 => "0000001110000000000111010100001000",
			2707 => "0000001100000000001000111000000100",
			2708 => "11111111101001010010101011111011",
			2709 => "11111110100001100010101011111011",
			2710 => "0000000101000000001111010000000100",
			2711 => "00000000100000100010101011111011",
			2712 => "11111110110011100010101011111011",
			2713 => "0000000101000000000001000000011000",
			2714 => "0000000100000000000111011100001100",
			2715 => "0000001110000000000011001000001000",
			2716 => "0000001011000000000001111100000100",
			2717 => "00000001101101110010101011111011",
			2718 => "11111111000110110010101011111011",
			2719 => "00000001101010000010101011111011",
			2720 => "0000001001000000000001000100000100",
			2721 => "00000001110010100010101011111011",
			2722 => "0000000100000000001100111100000100",
			2723 => "00000000001001110010101011111011",
			2724 => "11111110000100000010101011111011",
			2725 => "0000001111000000001000000100011000",
			2726 => "0000001001000000000011101000010000",
			2727 => "0000001111000000001110000000001000",
			2728 => "0000000001000000001010011000000100",
			2729 => "11111110001000110010101011111011",
			2730 => "00000000000000000010101011111011",
			2731 => "0000001011000000000001001000000100",
			2732 => "00000000000000000010101011111011",
			2733 => "11111111011111110010101011111011",
			2734 => "0000000011000000001011110000000100",
			2735 => "00000010101000010010101011111011",
			2736 => "11111110110000110010101011111011",
			2737 => "0000001000000000000001010100010000",
			2738 => "0000001011000000000000110100001000",
			2739 => "0000001001000000000011101000000100",
			2740 => "00011101011110100010101011111011",
			2741 => "00000000000000000010101011111011",
			2742 => "0000000011000000001100001100000100",
			2743 => "11111110101110000010101011111011",
			2744 => "00000110011111100010101011111011",
			2745 => "0000000000000000001011000100001000",
			2746 => "0000000001000000001010011000000100",
			2747 => "00000001000101100010101011111011",
			2748 => "11111111111010100010101011111011",
			2749 => "11111110011001010010101011111011",
			2750 => "0000000011000000001001110100100000",
			2751 => "0000000100000000000010010000001000",
			2752 => "0000001101000000001000011000000100",
			2753 => "11111110011101010010101111001101",
			2754 => "00000000000000000010101111001101",
			2755 => "0000001110000000001001110000010000",
			2756 => "0000000010000000000000010000000100",
			2757 => "11111110101010000010101111001101",
			2758 => "0000000010000000000000010000001000",
			2759 => "0000001010000000001000110000000100",
			2760 => "00000000101010000010101111001101",
			2761 => "00000000000000000010101111001101",
			2762 => "00000000000000000010101111001101",
			2763 => "0000000101000000000100011000000100",
			2764 => "00000001000111000010101111001101",
			2765 => "00000000000000000010101111001101",
			2766 => "0000000010000000000110010000101000",
			2767 => "0000000001000000001001111000001000",
			2768 => "0000001110000000001011000000000100",
			2769 => "00000010010101110010101111001101",
			2770 => "00000000000000000010101111001101",
			2771 => "0000000011000000000000011100001100",
			2772 => "0000000000000000000011010000000100",
			2773 => "11111110011111110010101111001101",
			2774 => "0000000011000000001000011000000100",
			2775 => "11111110100111010010101111001101",
			2776 => "00000000111011110010101111001101",
			2777 => "0000000000000000001111000100010000",
			2778 => "0000000001000000000111100100001000",
			2779 => "0000001100000000000100000000000100",
			2780 => "00000000001110100010101111001101",
			2781 => "11111101111001000010101111001101",
			2782 => "0000000100000000001100010000000100",
			2783 => "00000000000000000010101111001101",
			2784 => "00000001011101110010101111001101",
			2785 => "00000010000110000010101111001101",
			2786 => "0000000101000000001010111000001000",
			2787 => "0000000010000000000010000100000100",
			2788 => "00000000001110100010101111001101",
			2789 => "11111110011001110010101111001101",
			2790 => "0000001000000000001111000100011000",
			2791 => "0000000101000000000100011000001100",
			2792 => "0000000000000000000011111100000100",
			2793 => "11111110110010100010101111001101",
			2794 => "0000000110000000001011001100000100",
			2795 => "00000000010010010010101111001101",
			2796 => "00000001101111110010101111001101",
			2797 => "0000001101000000001000000000000100",
			2798 => "11111101101110010010101111001101",
			2799 => "0000000100000000000010111000000100",
			2800 => "00000000010011110010101111001101",
			2801 => "11111111101101000010101111001101",
			2802 => "11111110010000010010101111001101",
			2803 => "0000000011000000001001110100100000",
			2804 => "0000000110000000001011001100001000",
			2805 => "0000000001000000000111100100000100",
			2806 => "11111110011011000010110011010001",
			2807 => "00000000000000000010110011010001",
			2808 => "0000001001000000001011101000010000",
			2809 => "0000000101000000000100001000000100",
			2810 => "11111111011000100010110011010001",
			2811 => "0000001111000000000110100000001000",
			2812 => "0000000000000000000100011000000100",
			2813 => "00000001100101000010110011010001",
			2814 => "00000000000000000010110011010001",
			2815 => "00000000000000000010110011010001",
			2816 => "0000000001000000001001111000000100",
			2817 => "11111101110100100010110011010001",
			2818 => "00000000000000000010110011010001",
			2819 => "0000001111000000000101001000100000",
			2820 => "0000001000000000001111001000010000",
			2821 => "0000000011000000000100000100000100",
			2822 => "11111110100001010010110011010001",
			2823 => "0000001111000000000001000000001000",
			2824 => "0000001111000000001110101000000100",
			2825 => "11111111100100110010110011010001",
			2826 => "00000010010001110010110011010001",
			2827 => "11111111100001000010110011010001",
			2828 => "0000000011000000000001101000001000",
			2829 => "0000000001000000001001111000000100",
			2830 => "00000001101101010010110011010001",
			2831 => "11111110011001110010110011010001",
			2832 => "0000001011000000001100101100000100",
			2833 => "00000001111110010010110011010001",
			2834 => "00000000000000000010110011010001",
			2835 => "0000000011000000000010001000100000",
			2836 => "0000001011000000001100101100010100",
			2837 => "0000001111000000001110010000010000",
			2838 => "0000000110000000001011001100001000",
			2839 => "0000001011000000000101101100000100",
			2840 => "11111111111111000010110011010001",
			2841 => "11111110011110000010110011010001",
			2842 => "0000000011000000000001011000000100",
			2843 => "00000000000000000010110011010001",
			2844 => "00000001101100000010110011010001",
			2845 => "11111101101110100010110011010001",
			2846 => "0000000010000000001100010000000100",
			2847 => "11111011111110100010110011010001",
			2848 => "0000000110000000001111000000000100",
			2849 => "11111110101000000010110011010001",
			2850 => "00000000000000000010110011010001",
			2851 => "0000000001000000000110101000001000",
			2852 => "0000000000000000001110111100000100",
			2853 => "11111101100100010010110011010001",
			2854 => "00000000111100100010110011010001",
			2855 => "0000000101000000001000000000001100",
			2856 => "0000001111000000000010000000001000",
			2857 => "0000000101000000000100011000000100",
			2858 => "00000000100110000010110011010001",
			2859 => "00000001101011100010110011010001",
			2860 => "00000000000000000010110011010001",
			2861 => "0000000001000000000000111100001000",
			2862 => "0000000110000000001111000000000100",
			2863 => "11111111000111100010110011010001",
			2864 => "00000000010011010010110011010001",
			2865 => "0000000100000000001000001000000100",
			2866 => "00000000100011010010110011010001",
			2867 => "11111111110001110010110011010001",
			2868 => "0000000111000000001001110000110100",
			2869 => "0000001111000000000010011100100000",
			2870 => "0000000011000000000000011100011100",
			2871 => "0000000100000000000100001100001000",
			2872 => "0000000011000000001010001100000100",
			2873 => "11111110110001000010110111001101",
			2874 => "00000000000000000010110111001101",
			2875 => "0000001011000000000011011100001000",
			2876 => "0000000011000000001010111100000100",
			2877 => "11111111011101110010110111001101",
			2878 => "00000000000000000010110111001101",
			2879 => "0000001111000000000101001000001000",
			2880 => "0000000110000000001101011000000100",
			2881 => "00000000000000000010110111001101",
			2882 => "00000001001111000010110111001101",
			2883 => "11111111101111110010110111001101",
			2884 => "00000001010000010010110111001101",
			2885 => "0000000011000000000101110100010000",
			2886 => "0000001110000000000100000100001100",
			2887 => "0000000001000000001001111000001000",
			2888 => "0000000100000000000010100100000100",
			2889 => "11111111100111100010110111001101",
			2890 => "00000000000000000010110111001101",
			2891 => "00000000001000010010110111001101",
			2892 => "11111110010110000010110111001101",
			2893 => "00000000111111010010110111001101",
			2894 => "0000000111000000001001110000010000",
			2895 => "0000000011000000001000011000001000",
			2896 => "0000001100000000001100001000000100",
			2897 => "00000000000000000010110111001101",
			2898 => "11111111100010010010110111001101",
			2899 => "0000001000000000001001101000000100",
			2900 => "00000000000000000010110111001101",
			2901 => "00000001010111110010110111001101",
			2902 => "0000001101000000001000000000001000",
			2903 => "0000000100000000000010010000000100",
			2904 => "11111110101110110010110111001101",
			2905 => "00000000000000000010110111001101",
			2906 => "0000000101000000001000000000010100",
			2907 => "0000000110000000001001100100001000",
			2908 => "0000001100000000000100000000000100",
			2909 => "00000000000000000010110111001101",
			2910 => "11111111001011110010110111001101",
			2911 => "0000000000000000000011111100001000",
			2912 => "0000001111000000001110010000000100",
			2913 => "00000000111000100010110111001101",
			2914 => "11111111101001110010110111001101",
			2915 => "00000001100100010010110111001101",
			2916 => "0000001100000000001101010100010000",
			2917 => "0000001010000000001010110000001000",
			2918 => "0000000100000000001000000100000100",
			2919 => "00000000000000000010110111001101",
			2920 => "11111110100010100010110111001101",
			2921 => "0000000111000000000110000100000100",
			2922 => "00000000110100000010110111001101",
			2923 => "11111111101001010010110111001101",
			2924 => "0000000100000000000101010100001000",
			2925 => "0000001000000000000001110000000100",
			2926 => "00000000000110110010110111001101",
			2927 => "00000000110110110010110111001101",
			2928 => "0000001111000000001100001100000100",
			2929 => "11111111000100000010110111001101",
			2930 => "00000000001111010010110111001101",
			2931 => "0000001011000000000011011100001100",
			2932 => "0000000100000000000110110000000100",
			2933 => "11111110101010010010111010001001",
			2934 => "0000000000000000000110000100000100",
			2935 => "00000000000000000010111010001001",
			2936 => "11111111110111100010111010001001",
			2937 => "0000000111000000001000111000010000",
			2938 => "0000000110000000001011001100000100",
			2939 => "11111111111100010010111010001001",
			2940 => "0000000111000000001000111100001000",
			2941 => "0000000111000000000100000000000100",
			2942 => "00000000011100110010111010001001",
			2943 => "00000000000000000010111010001001",
			2944 => "00000001010101000010111010001001",
			2945 => "0000000111000000001001110000001000",
			2946 => "0000000100000000001000000100000100",
			2947 => "00000000000000000010111010001001",
			2948 => "11111110000100010010111010001001",
			2949 => "0000001101000000000111111100011100",
			2950 => "0000001110000000001011101100010000",
			2951 => "0000001010000000001010110000001000",
			2952 => "0000000100000000001000000100000100",
			2953 => "00000000001000110010111010001001",
			2954 => "11111110111100110010111010001001",
			2955 => "0000001001000000001001011000000100",
			2956 => "11111111101110100010111010001001",
			2957 => "00000000101101000010111010001001",
			2958 => "0000000101000000000101001000001000",
			2959 => "0000000001000000000111101000000100",
			2960 => "00000000000000000010111010001001",
			2961 => "00000001010100110010111010001001",
			2962 => "00000000000000000010111010001001",
			2963 => "0000000101000000001001010000010000",
			2964 => "0000001101000000001110010000001000",
			2965 => "0000001110000000001111101000000100",
			2966 => "11111111000100000010111010001001",
			2967 => "00000000100001000010111010001001",
			2968 => "0000000011000000001110000000000100",
			2969 => "11111101001110010010111010001001",
			2970 => "00000000000000000010111010001001",
			2971 => "0000001000000000000001010100001000",
			2972 => "0000000111000000000100010000000100",
			2973 => "00000000100110000010111010001001",
			2974 => "00000000000000000010111010001001",
			2975 => "0000001011000000000101110100000100",
			2976 => "00000000110010100010111010001001",
			2977 => "11111111101000100010111010001001",
			2978 => "0000000101000000000111001000010100",
			2979 => "0000000100000000000001101100001000",
			2980 => "0000000011000000001000011000000100",
			2981 => "11111110011011000010111110011101",
			2982 => "00000000000000000010111110011101",
			2983 => "0000001011000000000011011100001000",
			2984 => "0000000011000000000100001000000100",
			2985 => "11111111010101110010111110011101",
			2986 => "00000000000000000010111110011101",
			2987 => "00000000111001000010111110011101",
			2988 => "0000001111000000001111010000110100",
			2989 => "0000000111000000001001110000011000",
			2990 => "0000001010000000001010110000001100",
			2991 => "0000001100000000000100000000000100",
			2992 => "11111110101010010010111110011101",
			2993 => "0000001100000000000100000000000100",
			2994 => "00000001001100100010111110011101",
			2995 => "00000000000000000010111110011101",
			2996 => "0000000011000000001001110100000100",
			2997 => "00000000000000000010111110011101",
			2998 => "0000001100000000000100000000000100",
			2999 => "00000001101011000010111110011101",
			3000 => "00000000100110110010111110011101",
			3001 => "0000001110000000001011011100010100",
			3002 => "0000001111000000001100100100001000",
			3003 => "0000000000000000000001110100000100",
			3004 => "00000000000000000010111110011101",
			3005 => "11111110011000100010111110011101",
			3006 => "0000001010000000001100011100000100",
			3007 => "11111111001001010010111110011101",
			3008 => "0000001100000000001001110000000100",
			3009 => "00000000110001010010111110011101",
			3010 => "00000000000000000010111110011101",
			3011 => "0000000110000000000111101000000100",
			3012 => "00000000000000000010111110011101",
			3013 => "00000001001100110010111110011101",
			3014 => "0000001001000000001110010100101000",
			3015 => "0000001110000000000101110100011000",
			3016 => "0000000011000000000001011000001000",
			3017 => "0000000110000000001111000000000100",
			3018 => "11111110001011110010111110011101",
			3019 => "00000000000000000010111110011101",
			3020 => "0000001101000000000001101000001000",
			3021 => "0000001111000000001110010000000100",
			3022 => "00000000110011110010111110011101",
			3023 => "11111111011100110010111110011101",
			3024 => "0000000011000000000111110000000100",
			3025 => "11111110010111000010111110011101",
			3026 => "00000000100010110010111110011101",
			3027 => "0000000011000000000001001000000100",
			3028 => "11111101111011010010111110011101",
			3029 => "0000001011000000001100101000000100",
			3030 => "00000000111000100010111110011101",
			3031 => "0000000110000000000100111100000100",
			3032 => "00000000001101000010111110011101",
			3033 => "11111110100100100010111110011101",
			3034 => "0000000101000000001000011000001000",
			3035 => "0000000000000000001000110000000100",
			3036 => "00000000000000000010111110011101",
			3037 => "00000001100100010010111110011101",
			3038 => "0000000011000000000111100000000100",
			3039 => "11111110011000100010111110011101",
			3040 => "0000001101000000001011101100001000",
			3041 => "0000001111000000001000110100000100",
			3042 => "11111111110110100010111110011101",
			3043 => "00000000100000010010111110011101",
			3044 => "0000001110000000000001101100000100",
			3045 => "11111110011010100010111110011101",
			3046 => "00000000000000000010111110011101",
			3047 => "0000000101000000001010111000100100",
			3048 => "0000000100000000001111100000001100",
			3049 => "0000000111000000001001110000000100",
			3050 => "11111110010111000011000010111001",
			3051 => "0000000111000000001101100000000100",
			3052 => "00000000000000000011000010111001",
			3053 => "11111111011110100011000010111001",
			3054 => "0000001101000000000001111100000100",
			3055 => "11111110100111100011000010111001",
			3056 => "0000001111000000001110000100010000",
			3057 => "0000000110000000001011001100001100",
			3058 => "0000001010000000000110011100001000",
			3059 => "0000001010000000001100011100000100",
			3060 => "00000000000000000011000010111001",
			3061 => "00000000011001010011000010111001",
			3062 => "11111111110111110011000010111001",
			3063 => "00000001011011110011000010111001",
			3064 => "11111110111001110011000010111001",
			3065 => "0000000101000000000100011000100000",
			3066 => "0000001101000000001011000000010100",
			3067 => "0000001011000000000101101100001000",
			3068 => "0000001001000000001111001100000100",
			3069 => "00000000000000000011000010111001",
			3070 => "11111110100000110011000010111001",
			3071 => "0000000111000000001001110000001000",
			3072 => "0000000110000000001101011000000100",
			3073 => "00000000000000000011000010111001",
			3074 => "00000001100010110011000010111001",
			3075 => "11111111110101000011000010111001",
			3076 => "0000000110000000001101011000000100",
			3077 => "00000000000000000011000010111001",
			3078 => "0000000111000000001101100000000100",
			3079 => "00000001101010000011000010111001",
			3080 => "00000000000000000011000010111001",
			3081 => "0000001101000000001000000000011000",
			3082 => "0000000100000000000010100100010000",
			3083 => "0000001111000000000101110000001100",
			3084 => "0000000111000000001001110000000100",
			3085 => "00000000001011110011000010111001",
			3086 => "0000000001000000001001111000000100",
			3087 => "00000000000000000011000010111001",
			3088 => "11111110000110110011000010111001",
			3089 => "11111101101011000011000010111001",
			3090 => "0000001011000000001100101100000100",
			3091 => "00000000110000110011000010111001",
			3092 => "00000000000000000011000010111001",
			3093 => "0000001011000000001100101100010100",
			3094 => "0000000000000000000000111000010000",
			3095 => "0000001101000000001001001000001000",
			3096 => "0000000001000000000110101000000100",
			3097 => "00000000001111000011000010111001",
			3098 => "11111110011001010011000010111001",
			3099 => "0000001011000000001100101100000100",
			3100 => "00000000001011010011000010111001",
			3101 => "00000001110000100011000010111001",
			3102 => "00000001110111100011000010111001",
			3103 => "0000001110000000000101100100010000",
			3104 => "0000000000000000000001110100001000",
			3105 => "0000000111000000001100101000000100",
			3106 => "00000000000000000011000010111001",
			3107 => "00000000001000100011000010111001",
			3108 => "0000000110000000001111000000000100",
			3109 => "11111101111000100011000010111001",
			3110 => "00000000000000000011000010111001",
			3111 => "0000000111000000001101100000001000",
			3112 => "0000000001000000000111100100000100",
			3113 => "00000000000000000011000010111001",
			3114 => "00000001100010110011000010111001",
			3115 => "0000001001000000001100011000000100",
			3116 => "11111111000001000011000010111001",
			3117 => "00000000001101010011000010111001",
			3118 => "0000000000000000000011010000110100",
			3119 => "0000000001000000000110101000001000",
			3120 => "0000000100000000000010110000000100",
			3121 => "11111110011100000011000111011101",
			3122 => "00000000000000000011000111011101",
			3123 => "0000000000000000000011010000101000",
			3124 => "0000001100000000000100000000001000",
			3125 => "0000000110000000001011001100000100",
			3126 => "00000000000000000011000111011101",
			3127 => "00000001001010010011000111011101",
			3128 => "0000000111000000000001111100010000",
			3129 => "0000000010000000001001100000001000",
			3130 => "0000000100000000001110000000000100",
			3131 => "00000000000000000011000111011101",
			3132 => "00000000100001100011000111011101",
			3133 => "0000000110000000001000010000000100",
			3134 => "11111111000000000011000111011101",
			3135 => "00000000000000000011000111011101",
			3136 => "0000001000000000001011010100001000",
			3137 => "0000001101000000001001011100000100",
			3138 => "00000000001100000011000111011101",
			3139 => "11111111101101110011000111011101",
			3140 => "0000001100000000000001101000000100",
			3141 => "00000001001010100011000111011101",
			3142 => "00000000000000000011000111011101",
			3143 => "11111110111011010011000111011101",
			3144 => "0000001100000000001100110000111100",
			3145 => "0000000110000000001001100100011100",
			3146 => "0000000010000000001110110100010000",
			3147 => "0000001110000000001110110000001000",
			3148 => "0000001110000000000111001000000100",
			3149 => "11111111011110010011000111011101",
			3150 => "00000000000000000011000111011101",
			3151 => "0000001010000000001010110000000100",
			3152 => "00000000000000000011000111011101",
			3153 => "00000001010001000011000111011101",
			3154 => "0000000100000000000011011000001000",
			3155 => "0000000111000000000100000000000100",
			3156 => "00000000000000000011000111011101",
			3157 => "11111110101101010011000111011101",
			3158 => "00000000000000000011000111011101",
			3159 => "0000001010000000001001101000011000",
			3160 => "0000000110000000000100111100010000",
			3161 => "0000000010000000001111010100001000",
			3162 => "0000000100000000001000001000000100",
			3163 => "00000000000000000011000111011101",
			3164 => "00000000101110110011000111011101",
			3165 => "0000001111000000000011001000000100",
			3166 => "00000000000000000011000111011101",
			3167 => "11111111011011000011000111011101",
			3168 => "0000000000000000000011010000000100",
			3169 => "00000000000000000011000111011101",
			3170 => "00000001011100000011000111011101",
			3171 => "0000001010000000001111001000000100",
			3172 => "11111111010110100011000111011101",
			3173 => "00000000000000000011000111011101",
			3174 => "0000000000000000000000111000001100",
			3175 => "0000001100000000001000011000001000",
			3176 => "0000000110000000001000010000000100",
			3177 => "00000000000000000011000111011101",
			3178 => "00000000110001110011000111011101",
			3179 => "00000000000000000011000111011101",
			3180 => "0000001110000000000011010100010000",
			3181 => "0000000100000000000111011100001100",
			3182 => "0000001000000000000001110100001000",
			3183 => "0000001000000000000111000100000100",
			3184 => "00000000000000000011000111011101",
			3185 => "11111111000011100011000111011101",
			3186 => "00000000001001110011000111011101",
			3187 => "11111110101000000011000111011101",
			3188 => "0000000111000000001001010100000100",
			3189 => "00000000101101000011000111011101",
			3190 => "11111111111110100011000111011101",
			3191 => "0000000011000000001001110100010100",
			3192 => "0000000110000000001011001100001000",
			3193 => "0000000001000000000111100100000100",
			3194 => "11111110011011010011001010110001",
			3195 => "00000000000000000011001010110001",
			3196 => "0000000111000000001101100000001000",
			3197 => "0000001011000000001001110000000100",
			3198 => "11111111010110000011001010110001",
			3199 => "00000001011011010011001010110001",
			3200 => "11111101101101100011001010110001",
			3201 => "0000000000000000001001110001010100",
			3202 => "0000000000000000000011010000100100",
			3203 => "0000000011000000000000011100001000",
			3204 => "0000000000000000000011111100000100",
			3205 => "11111110011001010011001010110001",
			3206 => "11111011101110100011001010110001",
			3207 => "0000001111000000001001010000001100",
			3208 => "0000000000000000000010011000001000",
			3209 => "0000000111000000000001111100000100",
			3210 => "11111111101110000011001010110001",
			3211 => "00000001011100010011001010110001",
			3212 => "00000010010101000011001010110001",
			3213 => "0000000001000000000111100100001000",
			3214 => "0000001111000000000011001000000100",
			3215 => "11111111110100110011001010110001",
			3216 => "11111101001101010011001010110001",
			3217 => "0000000101000000000001101000000100",
			3218 => "00000001011100100011001010110001",
			3219 => "00000000000100100011001010110001",
			3220 => "0000000000000000001110111100010000",
			3221 => "0000001010000000001010110000000100",
			3222 => "11111110110011110011001010110001",
			3223 => "0000001100000000001111011100001000",
			3224 => "0000000110000000001111000000000100",
			3225 => "00000000100001110011001010110001",
			3226 => "00000001010111000011001010110001",
			3227 => "11111110111100000011001010110001",
			3228 => "0000001010000000000101000100010000",
			3229 => "0000001000000000000010101000001000",
			3230 => "0000001010000000000110011100000100",
			3231 => "11111110101000110011001010110001",
			3232 => "00000000111011010011001010110001",
			3233 => "0000001111000000000111111100000100",
			3234 => "11111111111111010011001010110001",
			3235 => "11111101111101010011001010110001",
			3236 => "0000001100000000000110000100001000",
			3237 => "0000000000000000001000111100000100",
			3238 => "00000001011001010011001010110001",
			3239 => "00000000000000000011001010110001",
			3240 => "0000001011000000001110101000000100",
			3241 => "11111110011111110011001010110001",
			3242 => "00000001001100000011001010110001",
			3243 => "11111110001100000011001010110001",
			3244 => "0000000111000000001001110000111100",
			3245 => "0000001111000000000010011100100100",
			3246 => "0000000011000000000000011100100000",
			3247 => "0000000100000000000100001100001000",
			3248 => "0000000011000000001010001100000100",
			3249 => "11111110110100010011001111110101",
			3250 => "00000000000000000011001111110101",
			3251 => "0000001011000000000011011100001100",
			3252 => "0000000010000000000111011000001000",
			3253 => "0000000111000000001000111000000100",
			3254 => "11111111010110010011001111110101",
			3255 => "00000000000000000011001111110101",
			3256 => "00000000000000000011001111110101",
			3257 => "0000001111000000000101001000001000",
			3258 => "0000000110000000001101011000000100",
			3259 => "00000000000000000011001111110101",
			3260 => "00000001001011100011001111110101",
			3261 => "11111111110001000011001111110101",
			3262 => "00000001001101100011001111110101",
			3263 => "0000000011000000000101110100010100",
			3264 => "0000000001000000000110101000010000",
			3265 => "0000000111000000001000111000001100",
			3266 => "0000000100000000001010110100000100",
			3267 => "00000000011100110011001111110101",
			3268 => "0000000100000000000011010100000100",
			3269 => "11111111110000000011001111110101",
			3270 => "00000000000000000011001111110101",
			3271 => "11111111001010100011001111110101",
			3272 => "11111110011011010011001111110101",
			3273 => "00000000111101000011001111110101",
			3274 => "0000000111000000001001110000011000",
			3275 => "0000000000000000000000110000001100",
			3276 => "0000000110000000001101011000000100",
			3277 => "00000000000000000011001111110101",
			3278 => "0000001011000000001110001100000100",
			3279 => "00000001011111100011001111110101",
			3280 => "00000000000000000011001111110101",
			3281 => "0000000101000000000111001000001000",
			3282 => "0000000101000000001101010100000100",
			3283 => "00000000000000000011001111110101",
			3284 => "11111111110001010011001111110101",
			3285 => "00000000000000000011001111110101",
			3286 => "0000000011000000001011011100011100",
			3287 => "0000001010000000000110011100001100",
			3288 => "0000000111000000001100101000001000",
			3289 => "0000001011000000000110000100000100",
			3290 => "00000000000000000011001111110101",
			3291 => "11111110100010010011001111110101",
			3292 => "00000000000000000011001111110101",
			3293 => "0000000011000000001001110100001000",
			3294 => "0000001101000000000100011000000100",
			3295 => "00000000000000000011001111110101",
			3296 => "11111111110001110011001111110101",
			3297 => "0000000111000000001101100000000100",
			3298 => "00000000110101100011001111110101",
			3299 => "00000000000000000011001111110101",
			3300 => "0000000101000000001001110100010100",
			3301 => "0000000000000000000011111100001100",
			3302 => "0000000001000000000111100100000100",
			3303 => "11111111001001100011001111110101",
			3304 => "0000000110000000001001100100000100",
			3305 => "11111111101101010011001111110101",
			3306 => "00000001001011010011001111110101",
			3307 => "0000000100000000000000010100000100",
			3308 => "00000001100100010011001111110101",
			3309 => "00000000000000000011001111110101",
			3310 => "0000001011000000001010111000010000",
			3311 => "0000000110000000001000010000001000",
			3312 => "0000001011000000000000001100000100",
			3313 => "00000000000000000011001111110101",
			3314 => "11111110101010100011001111110101",
			3315 => "0000001011000000000001111100000100",
			3316 => "00000000011101000011001111110101",
			3317 => "00000000000000000011001111110101",
			3318 => "0000000000000000000010011000001000",
			3319 => "0000000101000000000001000000000100",
			3320 => "00000000011001110011001111110101",
			3321 => "11111111111110010011001111110101",
			3322 => "0000001010000000001010110000000100",
			3323 => "11111110100010100011001111110101",
			3324 => "00000000000000000011001111110101",
			3325 => "0000000110000000000100111101011100",
			3326 => "0000000111000000000001101001010100",
			3327 => "0000000001000000001101101000111000",
			3328 => "0000000101000000000011100000100000",
			3329 => "0000001101000000001011000000010000",
			3330 => "0000001100000000001100001000001000",
			3331 => "0000000101000000001010111100000100",
			3332 => "11111111010111110011010100011001",
			3333 => "00000000100001010011010100011001",
			3334 => "0000001000000000000001110100000100",
			3335 => "11111110111100100011010100011001",
			3336 => "00000000000000000011010100011001",
			3337 => "0000001100000000000100000000001000",
			3338 => "0000000111000000001001110000000100",
			3339 => "11111110111101100011010100011001",
			3340 => "00000000010011000011010100011001",
			3341 => "0000000111000000001101100000000100",
			3342 => "00000001000001110011010100011001",
			3343 => "11111111111111110011010100011001",
			3344 => "0000001100000000000100000000001100",
			3345 => "0000001010000000001010110000001000",
			3346 => "0000001001000000000101011100000100",
			3347 => "00000000100111010011010100011001",
			3348 => "00000000000000000011010100011001",
			3349 => "11111111011100010011010100011001",
			3350 => "0000000110000000001111000000001000",
			3351 => "0000000001000000000111100100000100",
			3352 => "11111110100101100011010100011001",
			3353 => "00000000000000000011010100011001",
			3354 => "00000000000000000011010100011001",
			3355 => "0000001110000000000111010100010100",
			3356 => "0000001100000000000100011000001100",
			3357 => "0000001110000000001011011100000100",
			3358 => "00000000000000000011010100011001",
			3359 => "0000001001000000001010100000000100",
			3360 => "00000000110001000011010100011001",
			3361 => "00000000000000000011010100011001",
			3362 => "0000000101000000000110100000000100",
			3363 => "00000000000000000011010100011001",
			3364 => "11111111100111010011010100011001",
			3365 => "0000001010000000001000100100000100",
			3366 => "11111111001001010011010100011001",
			3367 => "00000000100001000011010100011001",
			3368 => "0000000111000000000101100100000100",
			3369 => "11111110010111100011010100011001",
			3370 => "00000000000000000011010100011001",
			3371 => "0000000101000000001010011100001100",
			3372 => "0000001100000000000000101000000100",
			3373 => "00000000000000000011010100011001",
			3374 => "0000000010000000001100000000000100",
			3375 => "00000000000000000011010100011001",
			3376 => "00000001010001010011010100011001",
			3377 => "0000001001000000001100011000001100",
			3378 => "0000000011000000000010000000000100",
			3379 => "11111110011111100011010100011001",
			3380 => "0000000001000000001101101000000100",
			3381 => "00000000101001110011010100011001",
			3382 => "00000000000000000011010100011001",
			3383 => "0000000101000000001010010100001000",
			3384 => "0000001100000000000011011100000100",
			3385 => "00000000000000000011010100011001",
			3386 => "00000001001010000011010100011001",
			3387 => "0000001110000000001111100100001000",
			3388 => "0000001001000000000111101100000100",
			3389 => "11111110110011010011010100011001",
			3390 => "00000000000000000011010100011001",
			3391 => "0000000000000000001111000100001000",
			3392 => "0000001010000000001000100100000100",
			3393 => "00000000000000000011010100011001",
			3394 => "00000000011111000011010100011001",
			3395 => "0000001010000000000001010000000100",
			3396 => "11111110111011100011010100011001",
			3397 => "00000000000111000011010100011001",
			3398 => "0000000110000000001011001101010000",
			3399 => "0000001001000000001000010000110000",
			3400 => "0000000110000000001101011000010100",
			3401 => "0000000001000000000110101000000100",
			3402 => "11111110010110000011011001100101",
			3403 => "0000000000000000000001110000000100",
			3404 => "11111110011001110011011001100101",
			3405 => "0000001111000000000010000100001000",
			3406 => "0000001100000000001110001100000100",
			3407 => "11111111101001100011011001100101",
			3408 => "00001010011110000011011001100101",
			3409 => "11111110011000100011011001100101",
			3410 => "0000000011000000001001110100000100",
			3411 => "11111110010111110011011001100101",
			3412 => "0000001111000000000001000000001100",
			3413 => "0000001100000000001000111100001000",
			3414 => "0000000000000000000000111000000100",
			3415 => "00000001100101110011011001100101",
			3416 => "00000110001101010011011001100101",
			3417 => "00000000010001110011011001100101",
			3418 => "0000001001000000001111000000001000",
			3419 => "0000000010000000001110110100000100",
			3420 => "00000000001111110011011001100101",
			3421 => "11111110010111100011011001100101",
			3422 => "00000110010000110011011001100101",
			3423 => "0000000010000000000000010000011100",
			3424 => "0000001010000000001010100000000100",
			3425 => "00000100101000010011011001100101",
			3426 => "0000001110000000000110010000001000",
			3427 => "0000001111000000000110010000000100",
			3428 => "00000001000111100011011001100101",
			3429 => "11111110011000110011011001100101",
			3430 => "0000001101000000001111010000001000",
			3431 => "0000000001000000000001111000000100",
			3432 => "00000100101010010011011001100101",
			3433 => "11111110101110000011011001100101",
			3434 => "0000001100000000000100011000000100",
			3435 => "00000000000100000011011001100101",
			3436 => "11111110011000010011011001100101",
			3437 => "00000011111011000011011001100101",
			3438 => "0000001100000000000001101000110100",
			3439 => "0000001010000000001000010100011000",
			3440 => "0000000001000000001011111100000100",
			3441 => "00000100100111010011011001100101",
			3442 => "0000001101000000000001000000001000",
			3443 => "0000001110000000000110111100000100",
			3444 => "11111110011000000011011001100101",
			3445 => "00000000010010100011011001100101",
			3446 => "0000000000000000001111001000000100",
			3447 => "11111110010111110011011001100101",
			3448 => "0000000100000000000001011100000100",
			3449 => "00001001011011000011011001100101",
			3450 => "00000000111111110011011001100101",
			3451 => "0000000100000000000011111000010100",
			3452 => "0000000101000000001101010100001000",
			3453 => "0000000100000000001101110100000100",
			3454 => "11111110011000100011011001100101",
			3455 => "00000001110100100011011001100101",
			3456 => "0000000000000000001010101100000100",
			3457 => "11111111100001010011011001100101",
			3458 => "0000000101000000000111111100000100",
			3459 => "00000010110100100011011001100101",
			3460 => "00000000100010010011011001100101",
			3461 => "0000000110000000001111000000000100",
			3462 => "11111110011100000011011001100101",
			3463 => "00000001110010000011011001100101",
			3464 => "0000001001000000001000010100011100",
			3465 => "0000000101000000000111111100001000",
			3466 => "0000000101000000000010011100000100",
			3467 => "11111110100010000011011001100101",
			3468 => "00000010111110000011011001100101",
			3469 => "0000000110000000001111000000000100",
			3470 => "00000001010110010011011001100101",
			3471 => "0000001101000000000110111100001000",
			3472 => "0000000001000000000101011100000100",
			3473 => "11111111111101010011011001100101",
			3474 => "11111110011000000011011001100101",
			3475 => "0000001010000000001010110000000100",
			3476 => "00000000000111010011011001100101",
			3477 => "11111110010110110011011001100101",
			3478 => "0000000011000000000100001100000100",
			3479 => "11111110100010110011011001100101",
			3480 => "00000100000010110011011001100101",
			3481 => "0000000011000000001001110100011000",
			3482 => "0000001010000000000001010100001000",
			3483 => "0000000001000000000111100100000100",
			3484 => "11111110011101000011011101010001",
			3485 => "00000000000000000011011101010001",
			3486 => "0000000111000000001101100000001100",
			3487 => "0000001011000000001001110000001000",
			3488 => "0000001011000000000100000000000100",
			3489 => "11111110110010010011011101010001",
			3490 => "00000000000000000011011101010001",
			3491 => "00000001010100110011011101010001",
			3492 => "11111110100010000011011101010001",
			3493 => "0000000000000000001001110001011100",
			3494 => "0000001101000000000110111100111100",
			3495 => "0000000101000000000001000000011100",
			3496 => "0000000111000000000001101000010000",
			3497 => "0000000000000000000011010000001000",
			3498 => "0000000011000000000000011100000100",
			3499 => "11111101110001110011011101010001",
			3500 => "00000000000100010011011101010001",
			3501 => "0000000000000000001010000000000100",
			3502 => "00000000111111110011011101010001",
			3503 => "00000000000011000011011101010001",
			3504 => "0000001111000000001010000100000100",
			3505 => "11111110110111100011011101010001",
			3506 => "0000001011000000001011011100000100",
			3507 => "00000001100011000011011101010001",
			3508 => "00000000010011110011011101010001",
			3509 => "0000000011000000000010010100010000",
			3510 => "0000000101000000000101110000001000",
			3511 => "0000000111000000001000011000000100",
			3512 => "11111111110001110011011101010001",
			3513 => "11111110001100000011011101010001",
			3514 => "0000000001000000001110010100000100",
			3515 => "00000000101000100011011101010001",
			3516 => "11111110110101000011011101010001",
			3517 => "0000001110000000001000101000001000",
			3518 => "0000000100000000001110000000000100",
			3519 => "00000000000000000011011101010001",
			3520 => "00000001111000010011011101010001",
			3521 => "0000000011000000000110111000000100",
			3522 => "11111110000010010011011101010001",
			3523 => "00000000000000000011011101010001",
			3524 => "0000000111000000000110110100001000",
			3525 => "0000000111000000001011011100000100",
			3526 => "00000001101000010011011101010001",
			3527 => "00000100111111100011011101010001",
			3528 => "0000001001000000000111101100001100",
			3529 => "0000000101000000001110110100000100",
			3530 => "00000000000000000011011101010001",
			3531 => "0000000000000000000011010000000100",
			3532 => "00000001011111000011011101010001",
			3533 => "00000000000000000011011101010001",
			3534 => "0000001011000000001111010000001000",
			3535 => "0000001100000000001010001100000100",
			3536 => "00000000011010110011011101010001",
			3537 => "11111110101000010011011101010001",
			3538 => "00000001000001110011011101010001",
			3539 => "11111110001111000011011101010001",
			3540 => "0000001000000000001001000100011100",
			3541 => "0000000111000000000001101000011000",
			3542 => "0000000111000000001100101000000100",
			3543 => "00000000000000000011100000101101",
			3544 => "0000001011000000001011011100010000",
			3545 => "0000001000000000000010101100000100",
			3546 => "00000000000000000011100000101101",
			3547 => "0000001101000000000101110000001000",
			3548 => "0000000101000000000111100000000100",
			3549 => "00000000111000000011100000101101",
			3550 => "00000000000000000011100000101101",
			3551 => "00000000000000000011100000101101",
			3552 => "00000000000000000011100000101101",
			3553 => "00000000000000000011100000101101",
			3554 => "0000000110000000001010011000000100",
			3555 => "11111110111010110011100000101101",
			3556 => "0000001011000000001100110000010100",
			3557 => "0000001101000000001110110000010000",
			3558 => "0000000111000000001000111000001000",
			3559 => "0000000111000000001100001000000100",
			3560 => "00000000000000000011100000101101",
			3561 => "00000000000000000011100000101101",
			3562 => "0000000111000000001001110000000100",
			3563 => "11111111111010000011100000101101",
			3564 => "00000000000000000011100000101101",
			3565 => "00000001000011010011100000101101",
			3566 => "0000000011000000000111110000011100",
			3567 => "0000000100000000000011110000001100",
			3568 => "0000000001000000000110101000000100",
			3569 => "11111110011110000011100000101101",
			3570 => "0000000100000000001000000100000100",
			3571 => "11111110111111010011100000101101",
			3572 => "00000000001110100011100000101101",
			3573 => "0000000011000000001010011100001000",
			3574 => "0000000010000000000110111100000100",
			3575 => "11111111000011100011100000101101",
			3576 => "00000000000000000011100000101101",
			3577 => "0000000010000000000010000100000100",
			3578 => "00000001001011000011100000101101",
			3579 => "00000000000000000011100000101101",
			3580 => "0000001111000000000110010000010000",
			3581 => "0000001011000000000000001100001000",
			3582 => "0000001110000000001001010100000100",
			3583 => "00000001010101100011100000101101",
			3584 => "00000000000000000011100000101101",
			3585 => "0000000111000000000001111100000100",
			3586 => "00000000000000000011100000101101",
			3587 => "00000000011000000011100000101101",
			3588 => "0000001000000000000111000100001000",
			3589 => "0000000100000000000011101100000100",
			3590 => "11111111111110000011100000101101",
			3591 => "00000000111001110011100000101101",
			3592 => "0000001110000000000011010100000100",
			3593 => "11111111011011010011100000101101",
			3594 => "00000000010111010011100000101101",
			3595 => "0000000011000000000110111001111100",
			3596 => "0000001101000000001001011101011100",
			3597 => "0000000011000000001011111000111100",
			3598 => "0000000010000000000110010000011100",
			3599 => "0000000010000000001100010100010000",
			3600 => "0000001110000000000010001000001000",
			3601 => "0000000110000000001001011000000100",
			3602 => "00000000000000000011100101111001",
			3603 => "11111111000101010011100101111001",
			3604 => "0000001011000000001000000000000100",
			3605 => "00000000010000100011100101111001",
			3606 => "00000000000000000011100101111001",
			3607 => "0000001100000000000100010100000100",
			3608 => "00000000000000000011100101111001",
			3609 => "0000001100000000000100000000000100",
			3610 => "00000001000100010011100101111001",
			3611 => "00000000000000010011100101111001",
			3612 => "0000000000000000000011010000010000",
			3613 => "0000000111000000000111001000001000",
			3614 => "0000001100000000001000111000000100",
			3615 => "11111111110111010011100101111001",
			3616 => "11111110101011000011100101111001",
			3617 => "0000001000000000001100011100000100",
			3618 => "11111111110011010011100101111001",
			3619 => "00000000011011110011100101111001",
			3620 => "0000000000000000000011010000001000",
			3621 => "0000001010000000001010110000000100",
			3622 => "00000000000000000011100101111001",
			3623 => "00000001001111010011100101111001",
			3624 => "0000000011000000001100010100000100",
			3625 => "11111111101111100011100101111001",
			3626 => "00000000010011100011100101111001",
			3627 => "0000000000000000000001110100010000",
			3628 => "0000000011000000001100111000001100",
			3629 => "0000000100000000000001011100000100",
			3630 => "00000000000000000011100101111001",
			3631 => "0000001100000000001011000000000100",
			3632 => "00000000010100010011100101111001",
			3633 => "00000000000000000011100101111001",
			3634 => "11111111101110110011100101111001",
			3635 => "0000001001000000000010101100001100",
			3636 => "0000000110000000001001111100001000",
			3637 => "0000001011000000000010001000000100",
			3638 => "00000001001011100011100101111001",
			3639 => "00000000000000000011100101111001",
			3640 => "00000000000000000011100101111001",
			3641 => "00000000000000000011100101111001",
			3642 => "0000000010000000000010010100010100",
			3643 => "0000001011000000000101110100001000",
			3644 => "0000001100000000001001110100000100",
			3645 => "11111111001001000011100101111001",
			3646 => "00000000000000000011100101111001",
			3647 => "0000001100000000000001101000001000",
			3648 => "0000000000000000001011010100000100",
			3649 => "00000000000000000011100101111001",
			3650 => "00000000111000100011100101111001",
			3651 => "00000000000000000011100101111001",
			3652 => "0000001001000000000111101100000100",
			3653 => "00000000000000000011100101111001",
			3654 => "0000001101000000001010001000000100",
			3655 => "00000000000000000011100101111001",
			3656 => "11111110010111010011100101111001",
			3657 => "0000001101000000001100111000100100",
			3658 => "0000001111000000001000110100001100",
			3659 => "0000000000000000000001110100000100",
			3660 => "00000000000000000011100101111001",
			3661 => "0000000011000000000110111000000100",
			3662 => "00000000000000000011100101111001",
			3663 => "11111111011011110011100101111001",
			3664 => "0000000111000000000001101000000100",
			3665 => "00000000000000000011100101111001",
			3666 => "0000001010000000001000100100000100",
			3667 => "00000000000000000011100101111001",
			3668 => "0000001001000000000000001000001000",
			3669 => "0000000110000000001001111100000100",
			3670 => "00000000001110110011100101111001",
			3671 => "00000000000000000011100101111001",
			3672 => "0000000110000000000100111100000100",
			3673 => "00000000000000000011100101111001",
			3674 => "00000000110000110011100101111001",
			3675 => "0000001100000000000101110100000100",
			3676 => "11111111000110100011100101111001",
			3677 => "00000000000000000011100101111001",
			3678 => "0000000001000000000100110101110000",
			3679 => "0000000010000000000110010000110000",
			3680 => "0000000010000000001100010100010000",
			3681 => "0000001110000000000010001000001000",
			3682 => "0000000110000000001001011000000100",
			3683 => "00000000000000000011101010111101",
			3684 => "11111111001000010011101010111101",
			3685 => "0000001011000000001000000000000100",
			3686 => "00000000001111000011101010111101",
			3687 => "00000000000000000011101010111101",
			3688 => "0000001100000000000100010100000100",
			3689 => "00000000000000000011101010111101",
			3690 => "0000001100000000000100000000001100",
			3691 => "0000000110000000001101011000000100",
			3692 => "00000000000000000011101010111101",
			3693 => "0000001011000000000011011100000100",
			3694 => "00000000000000000011101010111101",
			3695 => "00000001000111100011101010111101",
			3696 => "0000001100000000001000111000001000",
			3697 => "0000001101000000001001110100000100",
			3698 => "11111111010111100011101010111101",
			3699 => "00000000000000000011101010111101",
			3700 => "0000001001000000001100011000000100",
			3701 => "00000000101010100011101010111101",
			3702 => "00000000000000000011101010111101",
			3703 => "0000001101000000001100010000101100",
			3704 => "0000001101000000001001011100011100",
			3705 => "0000001101000000001001010100010000",
			3706 => "0000000111000000001101100000001000",
			3707 => "0000000100000000000011110000000100",
			3708 => "11111111011010000011101010111101",
			3709 => "00000000001001100011101010111101",
			3710 => "0000000110000000001000010000000100",
			3711 => "11111110110111100011101010111101",
			3712 => "00000000000000000011101010111101",
			3713 => "0000000001000000001111001100000100",
			3714 => "00000000111101000011101010111101",
			3715 => "0000000100000000000100001100000100",
			3716 => "00000000000011100011101010111101",
			3717 => "11111111001100000011101010111101",
			3718 => "0000001001000000000101010000001000",
			3719 => "0000000001000000000101011100000100",
			3720 => "00000000000000000011101010111101",
			3721 => "00000000001000110011101010111101",
			3722 => "0000001110000000001000110100000100",
			3723 => "11111110110101010011101010111101",
			3724 => "00000000000000000011101010111101",
			3725 => "0000001101000000000011000000010000",
			3726 => "0000000110000000001001111100001100",
			3727 => "0000000001000000000000111100000100",
			3728 => "00000000000000000011101010111101",
			3729 => "0000000101000000001100010100000100",
			3730 => "00000000000000000011101010111101",
			3731 => "00000000111001110011101010111101",
			3732 => "00000000000000000011101010111101",
			3733 => "00000000000000000011101010111101",
			3734 => "0000001100000000000101100100110000",
			3735 => "0000000001000000001100011000001100",
			3736 => "0000000111000000000111010000001000",
			3737 => "0000001110000000001000101000000100",
			3738 => "00000001000101110011101010111101",
			3739 => "00000000000000000011101010111101",
			3740 => "00000000000000000011101010111101",
			3741 => "0000000001000000001101011000010100",
			3742 => "0000001000000000000110001000010000",
			3743 => "0000001111000000001000110100001000",
			3744 => "0000000111000000001000011000000100",
			3745 => "00000000000000000011101010111101",
			3746 => "11111111100001100011101010111101",
			3747 => "0000000111000000000110110100000100",
			3748 => "00000000110001110011101010111101",
			3749 => "11111111111010110011101010111101",
			3750 => "11111111011100000011101010111101",
			3751 => "0000001111000000001000011100000100",
			3752 => "00000000000000000011101010111101",
			3753 => "0000001110000000001000000100000100",
			3754 => "00000000000000000011101010111101",
			3755 => "0000000110000000001000010000000100",
			3756 => "00000000000000000011101010111101",
			3757 => "00000000111001100011101010111101",
			3758 => "11111111001101100011101010111101",
			3759 => "0000000101000000001010111100001000",
			3760 => "0000001000000000000000101000000100",
			3761 => "11111110110011110011101110110001",
			3762 => "00000000000000000011101110110001",
			3763 => "0000001100000000000100000000010100",
			3764 => "0000000100000000000010111000001000",
			3765 => "0000001001000000000101011100000100",
			3766 => "11111111000101000011101110110001",
			3767 => "00000000011011010011101110110001",
			3768 => "0000000101000000001010111100000100",
			3769 => "00000000000000000011101110110001",
			3770 => "0000000110000000001101011000000100",
			3771 => "00000000000000000011101110110001",
			3772 => "00000001011010010011101110110001",
			3773 => "0000000100000000000011000000101100",
			3774 => "0000001011000000000000011100010100",
			3775 => "0000001010000000001001000100010000",
			3776 => "0000001100000000000100011000001000",
			3777 => "0000001110000000000001111100000100",
			3778 => "00000000000000000011101110110001",
			3779 => "11111111001110110011101110110001",
			3780 => "0000000000000000000110001000000100",
			3781 => "00000000000000000011101110110001",
			3782 => "00000000010000010011101110110001",
			3783 => "00000000101011110011101110110001",
			3784 => "0000000101000000000110100000001000",
			3785 => "0000000001000000001011111100000100",
			3786 => "00000000000000000011101110110001",
			3787 => "00000001100010110011101110110001",
			3788 => "0000001010000000000010101100001000",
			3789 => "0000001001000000000101010000000100",
			3790 => "11111111100010100011101110110001",
			3791 => "00000000110101110011101110110001",
			3792 => "0000000100000000001011101100000100",
			3793 => "11111111001010010011101110110001",
			3794 => "00000000000000000011101110110001",
			3795 => "0000000110000000000100111100011100",
			3796 => "0000001100000000001011000000010000",
			3797 => "0000000000000000000010011000001000",
			3798 => "0000000100000000001010110100000100",
			3799 => "11111110100000110011101110110001",
			3800 => "00000000000110000011101110110001",
			3801 => "0000000111000000001000111000000100",
			3802 => "00000000110011010011101110110001",
			3803 => "11111111100100110011101110110001",
			3804 => "0000000001000000001110010100000100",
			3805 => "00000000110110010011101110110001",
			3806 => "0000001000000000000101000100000100",
			3807 => "11111111011111110011101110110001",
			3808 => "00000000001011010011101110110001",
			3809 => "0000001011000000001101111000001000",
			3810 => "0000000001000000001001111000000100",
			3811 => "00000000000000000011101110110001",
			3812 => "00000001010111010011101110110001",
			3813 => "0000001100000000000001011000001000",
			3814 => "0000001001000000001110010100000100",
			3815 => "11111111000000000011101110110001",
			3816 => "00000000001011000011101110110001",
			3817 => "0000000101000000001111100100000100",
			3818 => "11111110101010110011101110110001",
			3819 => "00000000000000000011101110110001",
			3820 => "0000001011000000000011011100001000",
			3821 => "0000000010000000000111011000000100",
			3822 => "11111110101011110011110010111101",
			3823 => "00000000000000000011110010111101",
			3824 => "0000000000000000000000111001000000",
			3825 => "0000001000000000001111001000110100",
			3826 => "0000001010000000001010110000100000",
			3827 => "0000000100000000001000001000010000",
			3828 => "0000000001000000000111101000001000",
			3829 => "0000000001000000000111101000000100",
			3830 => "11111111111101100011110010111101",
			3831 => "11111101011000100011110010111101",
			3832 => "0000000000000000001010101100000100",
			3833 => "00000000000100100011110010111101",
			3834 => "00000000101110010011110010111101",
			3835 => "0000000010000000001110100100001000",
			3836 => "0000000000000000001111000100000100",
			3837 => "11111111110001100011110010111101",
			3838 => "11111101110110000011110010111101",
			3839 => "0000000100000000001110111000000100",
			3840 => "00000000100000010011110010111101",
			3841 => "11111111100001100011110010111101",
			3842 => "0000000000000000000011111100001100",
			3843 => "0000000001000000001011101000000100",
			3844 => "11111111011111010011110010111101",
			3845 => "0000000101000000000101110000000100",
			3846 => "00000001000000110011110010111101",
			3847 => "11111111111110010011110010111101",
			3848 => "0000000110000000001001111100000100",
			3849 => "00000001011101000011110010111101",
			3850 => "00000000000000000011110010111101",
			3851 => "0000000001000000001111001100000100",
			3852 => "11111110100100110011110010111101",
			3853 => "0000000001000000000100110100000100",
			3854 => "00000000000000000011110010111101",
			3855 => "11111111010100000011110010111101",
			3856 => "0000000010000000001010110100110000",
			3857 => "0000000000000000000000110000010100",
			3858 => "0000000100000000001101001000001000",
			3859 => "0000000110000000001111000000000100",
			3860 => "11111110011000110011110010111101",
			3861 => "00000000000101100011110010111101",
			3862 => "0000001001000000001111001100000100",
			3863 => "00000000000000000011110010111101",
			3864 => "0000001010000000001010110000000100",
			3865 => "00000000000000000011110010111101",
			3866 => "00000001101010000011110010111101",
			3867 => "0000001010000000001100011100001100",
			3868 => "0000000010000000000010000000001000",
			3869 => "0000000100000000000100001100000100",
			3870 => "00000000000000000011110010111101",
			3871 => "00000000001111110011110010111101",
			3872 => "11111110110010010011110010111101",
			3873 => "0000001000000000000010101000001000",
			3874 => "0000000110000000001011001100000100",
			3875 => "00000000000000000011110010111101",
			3876 => "00000001010001100011110010111101",
			3877 => "0000001010000000000101000100000100",
			3878 => "11111111001111000011110010111101",
			3879 => "00000000010000100011110010111101",
			3880 => "0000001110000000000010100100001000",
			3881 => "0000000110000000000100101100000100",
			3882 => "00000000000000000011110010111101",
			3883 => "11111110011010000011110010111101",
			3884 => "0000000110000000000000001000000100",
			3885 => "00000001000001010011110010111101",
			3886 => "11111111111110100011110010111101",
			3887 => "0000000100000000001000000101000100",
			3888 => "0000000100000000001111100100011000",
			3889 => "0000000011000000001010000100010100",
			3890 => "0000001010000000000010101100010000",
			3891 => "0000001011000000000101100100001100",
			3892 => "0000000001000000001011111100000100",
			3893 => "00000000000000000011111000101001",
			3894 => "0000001011000000000000011100000100",
			3895 => "00000000000000000011111000101001",
			3896 => "00000000111010010011111000101001",
			3897 => "00000000000000000011111000101001",
			3898 => "00000000000000000011111000101001",
			3899 => "11111111100110100011111000101001",
			3900 => "0000000011000000001100111000011100",
			3901 => "0000001100000000001110001100010000",
			3902 => "0000001100000000001000111000001000",
			3903 => "0000000011000000000010001000000100",
			3904 => "00000000000000000011111000101001",
			3905 => "00000000101110110011111000101001",
			3906 => "0000001100000000001001110000000100",
			3907 => "00000000000000000011111000101001",
			3908 => "11111111100001000011111000101001",
			3909 => "0000001100000000001000000000001000",
			3910 => "0000001001000000000010101100000100",
			3911 => "00000000111001100011111000101001",
			3912 => "00000000000000000011111000101001",
			3913 => "00000000000000000011111000101001",
			3914 => "0000001100000000001001001000001000",
			3915 => "0000000010000000000011000000000100",
			3916 => "11111111001101010011111000101001",
			3917 => "00000000000000000011111000101001",
			3918 => "0000001100000000000001101000000100",
			3919 => "00000000101001100011111000101001",
			3920 => "00000000000000000011111000101001",
			3921 => "0000000100000000001000110100001100",
			3922 => "0000000110000000001000010000001000",
			3923 => "0000000000000000000010011000000100",
			3924 => "11111110101111100011111000101001",
			3925 => "00000000000000000011111000101001",
			3926 => "00000000000000000011111000101001",
			3927 => "0000000010000000001011110000111000",
			3928 => "0000001011000000001110001100011100",
			3929 => "0000000011000000000001011000010000",
			3930 => "0000000001000000001001111000001000",
			3931 => "0000001011000000000011011100000100",
			3932 => "11111111111010000011111000101001",
			3933 => "00000000100100000011111000101001",
			3934 => "0000001011000000001100110000000100",
			3935 => "00000000000000000011111000101001",
			3936 => "11111111010101110011111000101001",
			3937 => "0000001111000000001001011100000100",
			3938 => "00000001010000110011111000101001",
			3939 => "0000000110000000001001100100000100",
			3940 => "11111111011101010011111000101001",
			3941 => "00000000001001110011111000101001",
			3942 => "0000000100000000001100001100001100",
			3943 => "0000000110000000000100111100000100",
			3944 => "00000000000000000011111000101001",
			3945 => "0000001010000000001000010100000100",
			3946 => "00000000000000000011111000101001",
			3947 => "00000000011110010011111000101001",
			3948 => "0000001010000000001100011100001000",
			3949 => "0000001001000000000111101100000100",
			3950 => "11111110110100000011111000101001",
			3951 => "00000000000000000011111000101001",
			3952 => "0000001011000000001101010100000100",
			3953 => "00000000100000000011111000101001",
			3954 => "11111111011000010011111000101001",
			3955 => "0000000110000000000100101100011000",
			3956 => "0000000100000000000110001100001100",
			3957 => "0000000011000000001100001100001000",
			3958 => "0000001011000000001011110100000100",
			3959 => "00000000000000000011111000101001",
			3960 => "11111111101010000011111000101001",
			3961 => "00000000000000000011111000101001",
			3962 => "0000001010000000000001110000001000",
			3963 => "0000001110000000000101010100000100",
			3964 => "00000000100110000011111000101001",
			3965 => "00000000000000000011111000101001",
			3966 => "00000000000000000011111000101001",
			3967 => "0000001110000000000011010100010000",
			3968 => "0000000010000000001101001000001000",
			3969 => "0000000001000000000100110100000100",
			3970 => "00000000000000000011111000101001",
			3971 => "00000000000001000011111000101001",
			3972 => "0000001000000000000111000100000100",
			3973 => "00000000000000000011111000101001",
			3974 => "11111110101100000011111000101001",
			3975 => "0000001101000000001011101100000100",
			3976 => "00000000010101000011111000101001",
			3977 => "00000000000000000011111000101001",
			3978 => "0000000000000000001111000101011100",
			3979 => "0000000111000000001100101000010000",
			3980 => "0000001100000000001000111000001000",
			3981 => "0000000110000000001011001100000100",
			3982 => "00000000000000000011111110111101",
			3983 => "00000000000110100011111110111101",
			3984 => "0000000111000000001001110000000100",
			3985 => "00000000000000000011111110111101",
			3986 => "11111111001010010011111110111101",
			3987 => "0000001101000000001001011100100100",
			3988 => "0000000000000000000111000100010100",
			3989 => "0000001010000000000011101000001100",
			3990 => "0000000101000000000111100000001000",
			3991 => "0000001100000000001000000000000100",
			3992 => "00000000011011110011111110111101",
			3993 => "00000000000000000011111110111101",
			3994 => "00000000000000000011111110111101",
			3995 => "0000001000000000000110011100000100",
			3996 => "11111111011011100011111110111101",
			3997 => "00000000000000000011111110111101",
			3998 => "0000001001000000001010100100001100",
			3999 => "0000001100000000001110001100000100",
			4000 => "00000000000000000011111110111101",
			4001 => "0000001010000000000111110100000100",
			4002 => "00000000000000000011111110111101",
			4003 => "00000000111010010011111110111101",
			4004 => "00000000000000000011111110111101",
			4005 => "0000001100000000001001001000001100",
			4006 => "0000000000000000001000101100001000",
			4007 => "0000000011000000001100111000000100",
			4008 => "00000000000000000011111110111101",
			4009 => "11111110111001110011111110111101",
			4010 => "00000000000000000011111110111101",
			4011 => "0000000110000000001000010000001100",
			4012 => "0000001101000000001100010100000100",
			4013 => "00000000000000000011111110111101",
			4014 => "0000000101000000000010000100000100",
			4015 => "00000000100101000011111110111101",
			4016 => "00000000000000000011111110111101",
			4017 => "0000001000000000001001101000001000",
			4018 => "0000001101000000001100010100000100",
			4019 => "00000000000000000011111110111101",
			4020 => "11111111100100010011111110111101",
			4021 => "0000001110000000001011110000000100",
			4022 => "00000000000000000011111110111101",
			4023 => "00000000010011110011111110111101",
			4024 => "0000000101000000001000000000101000",
			4025 => "0000001101000000001001001000100000",
			4026 => "0000000111000000001001110000010100",
			4027 => "0000001111000000001110010000010000",
			4028 => "0000001101000000001011000000001000",
			4029 => "0000001100000000001100001000000100",
			4030 => "00000000010011110011111110111101",
			4031 => "11111111101111010011111110111101",
			4032 => "0000000011000000001111011100000100",
			4033 => "00000000000000000011111110111101",
			4034 => "00000000111010110011111110111101",
			4035 => "11111111001101000011111110111101",
			4036 => "0000000011000000000001011000001000",
			4037 => "0000000010000000000111010100000100",
			4038 => "11111111000100110011111110111101",
			4039 => "00000000000000000011111110111101",
			4040 => "00000000000000000011111110111101",
			4041 => "0000000011000000000100000100000100",
			4042 => "00000000000000000011111110111101",
			4043 => "00000001000010010011111110111101",
			4044 => "0000000010000000001011110000100100",
			4045 => "0000001010000000000001010000001000",
			4046 => "0000001110000000000101100100000100",
			4047 => "00000000000000000011111110111101",
			4048 => "11111110101101010011111110111101",
			4049 => "0000000111000000000110000100010000",
			4050 => "0000001100000000000100000000001000",
			4051 => "0000001101000000000110100100000100",
			4052 => "00000000001001010011111110111101",
			4053 => "11111111010000100011111110111101",
			4054 => "0000000110000000001001100100000100",
			4055 => "00000000000000000011111110111101",
			4056 => "00000000111101110011111110111101",
			4057 => "0000001110000000001110110100001000",
			4058 => "0000001011000000001101111000000100",
			4059 => "00000000000000000011111110111101",
			4060 => "11111110111010010011111110111101",
			4061 => "00000000000111000011111110111101",
			4062 => "0000000110000000000100101100011000",
			4063 => "0000000010000000001000001000001100",
			4064 => "0000001100000000001011000000000100",
			4065 => "00000000001110110011111110111101",
			4066 => "0000001110000000001011110000000100",
			4067 => "11111111010010100011111110111101",
			4068 => "00000000000000000011111110111101",
			4069 => "0000000111000000000010001000001000",
			4070 => "0000001000000000000010101000000100",
			4071 => "00000000111101110011111110111101",
			4072 => "00000000000000000011111110111101",
			4073 => "00000000000000000011111110111101",
			4074 => "0000000010000000001010110100000100",
			4075 => "00000000001001100011111110111101",
			4076 => "0000001110000000001011100000000100",
			4077 => "11111110110010010011111110111101",
			4078 => "00000000000000000011111110111101",
			4079 => "0000000011000000000001101000111000",
			4080 => "0000000011000000001001110100101000",
			4081 => "0000000011000000001010111000011000",
			4082 => "0000000011000000000100001000000100",
			4083 => "11111110010101010100000100111001",
			4084 => "0000000010000000000111011000001100",
			4085 => "0000000010000000000110010000000100",
			4086 => "11111110010101010100000100111001",
			4087 => "0000000010000000000110010000000100",
			4088 => "00000000010011000100000100111001",
			4089 => "11111110100001100100000100111001",
			4090 => "0000000010000000000000010000000100",
			4091 => "00000001011111000100000100111001",
			4092 => "11111110110010010100000100111001",
			4093 => "0000001010000000000001110000001000",
			4094 => "0000001011000000001100101000000100",
			4095 => "11111110010101010100000100111001",
			4096 => "00000010011011110100000100111001",
			4097 => "0000000111000000001001110000000100",
			4098 => "00000100110001000100000100111001",
			4099 => "11111110011110010100000100111001",
			4100 => "0000000000000000000111111000000100",
			4101 => "11111110010101100100000100111001",
			4102 => "0000000111000000001101100000001000",
			4103 => "0000001111000000001001010000000100",
			4104 => "00000110010101010100000100111001",
			4105 => "11111110100000100100000100111001",
			4106 => "11111110011010110100000100111001",
			4107 => "0000001100000000000001101001101000",
			4108 => "0000001010000000001000100100110100",
			4109 => "0000001111000000000110111100011000",
			4110 => "0000000011000000001110101100001100",
			4111 => "0000000111000000000001111100000100",
			4112 => "11111110011001010100000100111001",
			4113 => "0000001111000000000101110100000100",
			4114 => "11111110110000000100000100111001",
			4115 => "00001010111100110100000100111001",
			4116 => "0000000001000000000101011100000100",
			4117 => "11111110010101110100000100111001",
			4118 => "0000001000000000001000100100000100",
			4119 => "00000011110111010100000100111001",
			4120 => "11111110110001110100000100111001",
			4121 => "0000000101000000000111100000010000",
			4122 => "0000001001000000001001111100001000",
			4123 => "0000001100000000000100011000000100",
			4124 => "00000011000100100100000100111001",
			4125 => "00001000010000100100000100111001",
			4126 => "0000001101000000000001000000000100",
			4127 => "11111110110110000100000100111001",
			4128 => "00000001101111100100000100111001",
			4129 => "0000001101000000001100010100000100",
			4130 => "11111110010110100100000100111001",
			4131 => "0000000001000000000100110100000100",
			4132 => "00000110110101110100000100111001",
			4133 => "11111110110000100100000100111001",
			4134 => "0000000011000000000001011000011100",
			4135 => "0000001100000000001000111100010000",
			4136 => "0000001010000000001010110000001000",
			4137 => "0000001101000000001000000000000100",
			4138 => "11111110011011100100000100111001",
			4139 => "00000000110111100100000100111001",
			4140 => "0000001101000000001110110000000100",
			4141 => "11111110011001100100000100111001",
			4142 => "00000100011100100100000100111001",
			4143 => "0000000111000000001101100000001000",
			4144 => "0000001111000000001111010000000100",
			4145 => "00000011100000110100000100111001",
			4146 => "11111110001110110100000100111001",
			4147 => "11111110010111000100000100111001",
			4148 => "0000000101000000000111111100010000",
			4149 => "0000001110000000000111010100001000",
			4150 => "0000001100000000001100110000000100",
			4151 => "00000100001101110100000100111001",
			4152 => "11111111110001010100000100111001",
			4153 => "0000000000000000001010101100000100",
			4154 => "00000010001111100100000100111001",
			4155 => "00000100011000100100000100111001",
			4156 => "0000000000000000000010111100000100",
			4157 => "11111110011000000100000100111001",
			4158 => "00000100111001000100000100111001",
			4159 => "0000001001000000001000010100011000",
			4160 => "0000001101000000001100010100000100",
			4161 => "00000010010001000100000100111001",
			4162 => "0000001011000000000001001000001000",
			4163 => "0000001100000000001000011000000100",
			4164 => "00000011101000010100000100111001",
			4165 => "11111110011101110100000100111001",
			4166 => "0000000101000000001110010000000100",
			4167 => "00000000001100100100000100111001",
			4168 => "0000000111000000000000011100000100",
			4169 => "11111111111101110100000100111001",
			4170 => "11111110011100000100000100111001",
			4171 => "0000000000000000000011010000000100",
			4172 => "11111110100110100100000100111001",
			4173 => "00000100011100100100000100111001",
			4174 => "0000000001000000000100110110001000",
			4175 => "0000000010000000000110111101000000",
			4176 => "0000000011000000000111110000100100",
			4177 => "0000001010000000000001010000001100",
			4178 => "0000000101000000000011100000000100",
			4179 => "00000000000000000100001010011101",
			4180 => "0000000100000000001000101000000100",
			4181 => "00000000000000000100001010011101",
			4182 => "11111110100111010100001010011101",
			4183 => "0000000111000000001101100000001100",
			4184 => "0000001001000000000001000100001000",
			4185 => "0000000111000000001001110000000100",
			4186 => "00000000000000000100001010011101",
			4187 => "00000000110100010100001010011101",
			4188 => "11111111100000100100001010011101",
			4189 => "0000000011000000000010001000001000",
			4190 => "0000000001000000000010001100000100",
			4191 => "00000000000000000100001010011101",
			4192 => "11111111001010110100001010011101",
			4193 => "00000000000000000100001010011101",
			4194 => "0000000011000000001101000100001000",
			4195 => "0000000110000000000111101000000100",
			4196 => "00000000000000000100001010011101",
			4197 => "00000001000010100100001010011101",
			4198 => "0000000010000000000110111100010000",
			4199 => "0000001100000000001001001000001000",
			4200 => "0000001100000000001010111000000100",
			4201 => "00000000000000000100001010011101",
			4202 => "11111111011011000100001010011101",
			4203 => "0000001100000000001001110100000100",
			4204 => "00000000001000000100001010011101",
			4205 => "00000000000000000100001010011101",
			4206 => "00000000001101010100001010011101",
			4207 => "0000000110000000001000010000110000",
			4208 => "0000001100000000001101010100011000",
			4209 => "0000001010000000001010110000001100",
			4210 => "0000001001000000000111101100001000",
			4211 => "0000000100000000000110111000000100",
			4212 => "00000000000000000100001010011101",
			4213 => "11111110100110100100001010011101",
			4214 => "00000000000000000100001010011101",
			4215 => "0000001000000000000111000100000100",
			4216 => "00000001001000100100001010011101",
			4217 => "0000001111000000001001011100000100",
			4218 => "00000000000000000100001010011101",
			4219 => "11111111000111110100001010011101",
			4220 => "0000000001000000001110010100001100",
			4221 => "0000000110000000001000010000001000",
			4222 => "0000000110000000001101011000000100",
			4223 => "11111111111001110100001010011101",
			4224 => "00000000110101100100001010011101",
			4225 => "11111111110001110100001010011101",
			4226 => "0000000111000000001000011000001000",
			4227 => "0000000111000000000001101000000100",
			4228 => "11111111110011110100001010011101",
			4229 => "00000000010100110100001010011101",
			4230 => "11111110100011010100001010011101",
			4231 => "0000001100000000000110000100001000",
			4232 => "0000001010000000001001101000000100",
			4233 => "00000000111101000100001010011101",
			4234 => "00000000000000000100001010011101",
			4235 => "0000001000000000000111000100001100",
			4236 => "0000000111000000001111011100000100",
			4237 => "00000000111101010100001010011101",
			4238 => "0000000010000000000010110000000100",
			4239 => "11111110111011010100001010011101",
			4240 => "00000000101101100100001010011101",
			4241 => "11111110111001100100001010011101",
			4242 => "0000001100000000000101100100101000",
			4243 => "0000000001000000001100011000001000",
			4244 => "0000000111000000000111010000000100",
			4245 => "00000000111101110100001010011101",
			4246 => "00000000000000000100001010011101",
			4247 => "0000000001000000001101011000011000",
			4248 => "0000000011000000001100001100010000",
			4249 => "0000001111000000001000110100001000",
			4250 => "0000000111000000001000011000000100",
			4251 => "00000000000000000100001010011101",
			4252 => "11111111100100000100001010011101",
			4253 => "0000000111000000000110110100000100",
			4254 => "00000000110001010100001010011101",
			4255 => "00000000000000000100001010011101",
			4256 => "0000000001000000001010011000000100",
			4257 => "11111111010111000100001010011101",
			4258 => "00000000000000000100001010011101",
			4259 => "0000000011000000001100001100000100",
			4260 => "00000000000000000100001010011101",
			4261 => "00000000110110010100001010011101",
			4262 => "11111111010000010100001010011101",
			4263 => "0000000100000000001100001101001100",
			4264 => "0000000000000000000010111101000100",
			4265 => "0000001100000000000100011000011100",
			4266 => "0000001010000000001010110000011000",
			4267 => "0000000000000000001111000100010000",
			4268 => "0000000100000000000010010100001000",
			4269 => "0000000000000000000110001000000100",
			4270 => "11111111110110000100001111101001",
			4271 => "00000000001001000100001111101001",
			4272 => "0000001001000000000111101100000100",
			4273 => "11111111000011010100001111101001",
			4274 => "00000000000000000100001111101001",
			4275 => "0000000011000000000001011000000100",
			4276 => "00000000000000000100001111101001",
			4277 => "00000000110001010100001111101001",
			4278 => "11111110111110000100001111101001",
			4279 => "0000001100000000000001101000010100",
			4280 => "0000000001000000001001011000000100",
			4281 => "00000000000000000100001111101001",
			4282 => "0000001001000000001010100100001000",
			4283 => "0000000010000000000110111000000100",
			4284 => "00000000101001000100001111101001",
			4285 => "00000000000000000100001111101001",
			4286 => "0000000100000000001110000000000100",
			4287 => "00000000001011000100001111101001",
			4288 => "00000000000000000100001111101001",
			4289 => "0000001111000000001000110100001000",
			4290 => "0000000101000000000110010000000100",
			4291 => "11111111100110010100001111101001",
			4292 => "00000000000000000100001111101001",
			4293 => "0000001000000000000001010100000100",
			4294 => "00000000000000000100001111101001",
			4295 => "0000000000000000001010101100000100",
			4296 => "00000000010010000100001111101001",
			4297 => "00000000000000000100001111101001",
			4298 => "0000000011000000000000011100000100",
			4299 => "00000000000000000100001111101001",
			4300 => "00000001000111010100001111101001",
			4301 => "0000000100000000000110001100010000",
			4302 => "0000001010000000001000010100000100",
			4303 => "00000000000000000100001111101001",
			4304 => "0000001100000000001000111100000100",
			4305 => "00000000000000000100001111101001",
			4306 => "0000000100000000001100001100000100",
			4307 => "00000000000000000100001111101001",
			4308 => "11111110011101100100001111101001",
			4309 => "0000000000000000001111000100010100",
			4310 => "0000000011000000000000010000000100",
			4311 => "00000000000000000100001111101001",
			4312 => "0000001001000000000011101000001100",
			4313 => "0000001010000000001010110000001000",
			4314 => "0000001000000000000001010100000100",
			4315 => "00000000000000000100001111101001",
			4316 => "00000000110000000100001111101001",
			4317 => "00000000000000000100001111101001",
			4318 => "00000000000000000100001111101001",
			4319 => "0000001010000000001010110000011000",
			4320 => "0000000010000000001110100100001100",
			4321 => "0000001110000000000110111000001000",
			4322 => "0000000000000000001111000100000100",
			4323 => "00000000000000000100001111101001",
			4324 => "11111110100011100100001111101001",
			4325 => "00000000000000000100001111101001",
			4326 => "0000000001000000001100011000001000",
			4327 => "0000001110000000001000001000000100",
			4328 => "00000000100001110100001111101001",
			4329 => "00000000000000000100001111101001",
			4330 => "00000000000000000100001111101001",
			4331 => "0000000010000000001111010100010000",
			4332 => "0000000011000000001011011100001000",
			4333 => "0000000010000000001100010000000100",
			4334 => "00000000011011100100001111101001",
			4335 => "11111111100000110100001111101001",
			4336 => "0000001010000000001100011100000100",
			4337 => "00000001010100000100001111101001",
			4338 => "00000000000000000100001111101001",
			4339 => "0000000000000000000000111000001000",
			4340 => "0000001110000000000010000100000100",
			4341 => "11111111000011110100001111101001",
			4342 => "00000000000000000100001111101001",
			4343 => "0000000000000000000111111000000100",
			4344 => "00000000010101100100001111101001",
			4345 => "11111111100101100100001111101001",
			4346 => "0000000011000000001001110100010100",
			4347 => "0000000001000000000111100100010000",
			4348 => "0000000011000000000100001000000100",
			4349 => "11111110010101100100010100011101",
			4350 => "0000001000000000001000110000000100",
			4351 => "11111110010101100100010100011101",
			4352 => "0000000111000000001001110000000100",
			4353 => "00000100010000000100010100011101",
			4354 => "11111110011100110100010100011101",
			4355 => "00000001110110000100010100011101",
			4356 => "0000001100000000000001101001100100",
			4357 => "0000001000000000000101000100101000",
			4358 => "0000000000000000001100000100001100",
			4359 => "0000000001000000000001000100001000",
			4360 => "0000001000000000001000010100000100",
			4361 => "11111110011000110100010100011101",
			4362 => "00000000110111110100010100011101",
			4363 => "00000011000110100100010100011101",
			4364 => "0000000100000000001000001100001100",
			4365 => "0000001101000000001111010000001000",
			4366 => "0000001100000000000100001000000100",
			4367 => "11111110101011100100010100011101",
			4368 => "00000101010011010100010100011101",
			4369 => "11111110011010110100010100011101",
			4370 => "0000000011000000001100010000001000",
			4371 => "0000001100000000000100011000000100",
			4372 => "11111110010111010100010100011101",
			4373 => "00000000001000010100010100011101",
			4374 => "0000000000000000000001110100000100",
			4375 => "11111111110010100100010100011101",
			4376 => "00000101111100110100010100011101",
			4377 => "0000000011000000000001011000100000",
			4378 => "0000000100000000001001001100010000",
			4379 => "0000000011000000000100000100001000",
			4380 => "0000000011000000001010001100000100",
			4381 => "11111110010101010100010100011101",
			4382 => "11111111100110100100010100011101",
			4383 => "0000000010000000001110110100000100",
			4384 => "00000011001010000100010100011101",
			4385 => "11111110001101110100010100011101",
			4386 => "0000001111000000001001010000001000",
			4387 => "0000000111000000001101100000000100",
			4388 => "00000100101101010100010100011101",
			4389 => "11111110011010100100010100011101",
			4390 => "0000000011000000000000011100000100",
			4391 => "11111110010110100100010100011101",
			4392 => "00000001000101100100010100011101",
			4393 => "0000000100000000000100001100010000",
			4394 => "0000001000000000000001110000001000",
			4395 => "0000000100000000001110000000000100",
			4396 => "00000100001000110100010100011101",
			4397 => "11111111110011000100010100011101",
			4398 => "0000000111000000000111010000000100",
			4399 => "00000011011101100100010100011101",
			4400 => "11111110011110000100010100011101",
			4401 => "0000001100000000001000111000000100",
			4402 => "00000011111000010100010100011101",
			4403 => "0000001111000000001000001100000100",
			4404 => "11111110010101100100010100011101",
			4405 => "00000001100011100100010100011101",
			4406 => "0000001001000000001000010100011100",
			4407 => "0000000101000000000111111100001000",
			4408 => "0000001110000000001011111000000100",
			4409 => "11111110011110000100010100011101",
			4410 => "00000011110111100100010100011101",
			4411 => "0000001000000000000110001000010000",
			4412 => "0000000100000000000011110100001000",
			4413 => "0000000001000000000001000100000100",
			4414 => "00001011111111110100010100011101",
			4415 => "11111110100010010100010100011101",
			4416 => "0000001000000000000110001000000100",
			4417 => "00100001011000100100010100011101",
			4418 => "00000101011100110100010100011101",
			4419 => "11111110010110000100010100011101",
			4420 => "0000000011000000000100001100000100",
			4421 => "11111110100000100100010100011101",
			4422 => "00000101101000000100010100011101",
			4423 => "0000001011000000000011011100001100",
			4424 => "0000001010000000001111001000000100",
			4425 => "11111110011010100100011000001001",
			4426 => "0000000000000000000111010000000100",
			4427 => "00000001000000000100011000001001",
			4428 => "00000000000000000100011000001001",
			4429 => "0000001010000000001001101001100100",
			4430 => "0000001000000000001010110000101000",
			4431 => "0000000100000000001111100100010100",
			4432 => "0000000011000000001010000100010000",
			4433 => "0000001111000000000110111100001000",
			4434 => "0000000101000000000110100000000100",
			4435 => "00000000110110110100011000001001",
			4436 => "11111111001000110100011000001001",
			4437 => "0000001011000000001011011100000100",
			4438 => "00000010110101010100011000001001",
			4439 => "11111111110100000100011000001001",
			4440 => "11111110100000110100011000001001",
			4441 => "0000001100000000001001110100010000",
			4442 => "0000001100000000000100011000001000",
			4443 => "0000001100000000001010111000000100",
			4444 => "00000000100100000100011000001001",
			4445 => "11111111101011010100011000001001",
			4446 => "0000001100000000001011000000000100",
			4447 => "00000011000001110100011000001001",
			4448 => "00000001011000000100011000001001",
			4449 => "11111111001000010100011000001001",
			4450 => "0000000100000000000010100100100000",
			4451 => "0000000011000000000000011100010000",
			4452 => "0000000100000000000010111000001000",
			4453 => "0000001111000000001111010000000100",
			4454 => "11111110010010100100011000001001",
			4455 => "11111100110110010100011000001001",
			4456 => "0000001100000000000000101000000100",
			4457 => "00000001101100100100011000001001",
			4458 => "11111111100001110100011000001001",
			4459 => "0000001111000000000010011100001000",
			4460 => "0000000111000000001101100000000100",
			4461 => "00000010001111000100011000001001",
			4462 => "00000000000000000100011000001001",
			4463 => "0000000011000000000101110100000100",
			4464 => "11111111001111010100011000001001",
			4465 => "00000000010000000100011000001001",
			4466 => "0000001011000000000110000100001100",
			4467 => "0000000101000000001010111100000100",
			4468 => "00000000000000000100011000001001",
			4469 => "0000001100000000001000111000000100",
			4470 => "00000001110101100100011000001001",
			4471 => "00000000100001110100011000001001",
			4472 => "0000000011000000001010001100001000",
			4473 => "0000000011000000001010011100000100",
			4474 => "11111101101111110100011000001001",
			4475 => "11111111110001010100011000001001",
			4476 => "0000000100000000001011100000000100",
			4477 => "00000001110010110100011000001001",
			4478 => "00000000010010100100011000001001",
			4479 => "0000001100000000001000111100000100",
			4480 => "00000001010100110100011000001001",
			4481 => "11111110000111010100011000001001",
			4482 => "0000000110000000001011001101100000",
			4483 => "0000001001000000001000010000111000",
			4484 => "0000000110000000001101011000011100",
			4485 => "0000000001000000000110101000000100",
			4486 => "11111110010110100100011110010101",
			4487 => "0000000000000000000001110000001100",
			4488 => "0000001101000000000100010000001000",
			4489 => "0000001011000000000100011000000100",
			4490 => "11111110011011110100011110010101",
			4491 => "00000100000110100100011110010101",
			4492 => "11111110010111100100011110010101",
			4493 => "0000001111000000000010000100001000",
			4494 => "0000000111000000001100101000000100",
			4495 => "11111110100010000100011110010101",
			4496 => "00000110000110110100011110010101",
			4497 => "11111110011010000100011110010101",
			4498 => "0000000011000000001001110100000100",
			4499 => "11111110011000010100011110010101",
			4500 => "0000001111000000000001000000001100",
			4501 => "0000001100000000001000111100001000",
			4502 => "0000000011000000000001101000000100",
			4503 => "00000010001111010100011110010101",
			4504 => "00000101011101100100011110010101",
			4505 => "00000000001110110100011110010101",
			4506 => "0000001001000000001111000000001000",
			4507 => "0000000010000000001110110100000100",
			4508 => "00000000001101100100011110010101",
			4509 => "11111110011000100100011110010101",
			4510 => "00000100100100000100011110010101",
			4511 => "0000000010000000001000001100011000",
			4512 => "0000001010000000001010100000000100",
			4513 => "00000011011001000100011110010101",
			4514 => "0000001100000000000100011000010000",
			4515 => "0000000011000000001100000000001000",
			4516 => "0000000010000000001110110100000100",
			4517 => "00000000000110100100011110010101",
			4518 => "11111110011010110100011110010101",
			4519 => "0000001101000000000101001000000100",
			4520 => "00000101001101000100011110010101",
			4521 => "11111111110100100100011110010101",
			4522 => "11111110011001100100011110010101",
			4523 => "0000000110000000001011001100001100",
			4524 => "0000001100000000001011000000000100",
			4525 => "00000110110010010100011110010101",
			4526 => "0000000110000000001101011000000100",
			4527 => "11111110110010000100011110010101",
			4528 => "00000001001000100100011110010101",
			4529 => "11111110100110100100011110010101",
			4530 => "0000001100000000000001101001000100",
			4531 => "0000001010000000001000010100011100",
			4532 => "0000000001000000001011111100000100",
			4533 => "00000011010011110100011110010101",
			4534 => "0000001110000000001100010000001000",
			4535 => "0000001010000000000011101000000100",
			4536 => "00000001101100100100011110010101",
			4537 => "11111110011000100100011110010101",
			4538 => "0000001011000000000110110100001000",
			4539 => "0000000001000000000111101000000100",
			4540 => "00001000000001010100011110010101",
			4541 => "00000001000000110100011110010101",
			4542 => "0000001101000000001100010100000100",
			4543 => "11111110000101100100011110010101",
			4544 => "00000001000011110100011110010101",
			4545 => "0000000000000000001100101100100000",
			4546 => "0000000110000000001001100100010000",
			4547 => "0000000111000000000101101100001000",
			4548 => "0000000101000000001101010100000100",
			4549 => "11111110011011110100011110010101",
			4550 => "00000010011011100100011110010101",
			4551 => "0000000010000000000011000000000100",
			4552 => "11111110010011010100011110010101",
			4553 => "00000000111111100100011110010101",
			4554 => "0000000111000000000111010000001000",
			4555 => "0000000000000000001010101100000100",
			4556 => "11111111101001110100011110010101",
			4557 => "00000010100001010100011110010101",
			4558 => "0000000011000000000110001100000100",
			4559 => "11111110010111000100011110010101",
			4560 => "00000010100110000100011110010101",
			4561 => "0000000110000000001111000000000100",
			4562 => "11111110011101110100011110010101",
			4563 => "00000000000000000100011110010101",
			4564 => "0000001001000000001000010100011100",
			4565 => "0000000101000000000111111100001000",
			4566 => "0000001111000000001011110000000100",
			4567 => "11111110011110110100011110010101",
			4568 => "00000010101010010100011110010101",
			4569 => "0000000110000000001111000000000100",
			4570 => "00000001001011000100011110010101",
			4571 => "0000001101000000000110111100001000",
			4572 => "0000000111000000000001011000000100",
			4573 => "11111111011101010100011110010101",
			4574 => "11111110010111000100011110010101",
			4575 => "0000001010000000001010110000000100",
			4576 => "00000000001101000100011110010101",
			4577 => "11111110010111010100011110010101",
			4578 => "0000000011000000000100001100000100",
			4579 => "11111110100101100100011110010101",
			4580 => "00000011001110010100011110010101",
			4581 => "0000001001000000000001111001010100",
			4582 => "0000001011000000001100101100101000",
			4583 => "0000000110000000001101011000000100",
			4584 => "11111110101110110100100011010001",
			4585 => "0000001100000000001001110000100000",
			4586 => "0000000010000000001100000000010000",
			4587 => "0000000011000000000100000100001000",
			4588 => "0000000100000000000100001100000100",
			4589 => "11111111011110000100100011010001",
			4590 => "00000000111010010100100011010001",
			4591 => "0000001110000000000101110100000100",
			4592 => "00000001011001000100100011010001",
			4593 => "00000000000000000100100011010001",
			4594 => "0000000010000000000111011000001000",
			4595 => "0000000111000000001000111000000100",
			4596 => "00000000000000000100100011010001",
			4597 => "11111110101111110100100011010001",
			4598 => "0000001101000000001011000000000100",
			4599 => "11111111010000010100100011010001",
			4600 => "00000000100110010100100011010001",
			4601 => "11111110000110100100100011010001",
			4602 => "0000000110000000001000010000100100",
			4603 => "0000000100000000000110001100011000",
			4604 => "0000001100000000001000111100001000",
			4605 => "0000000110000000001011001100000100",
			4606 => "00000000000000000100100011010001",
			4607 => "00000000111111100100100011010001",
			4608 => "0000001100000000000110000100001000",
			4609 => "0000000101000000001001001000000100",
			4610 => "00000000000000000100100011010001",
			4611 => "11111110101110110100100011010001",
			4612 => "0000000110000000000001000100000100",
			4613 => "00000000000000000100100011010001",
			4614 => "00000000101010100100100011010001",
			4615 => "0000000101000000000100011000000100",
			4616 => "00000000000000000100100011010001",
			4617 => "0000000011000000000000110100000100",
			4618 => "11111110010001000100100011010001",
			4619 => "11111111110011010100100011010001",
			4620 => "0000001001000000001110010100000100",
			4621 => "00000000111001100100100011010001",
			4622 => "00000000000000000100100011010001",
			4623 => "0000000101000000001010011100000100",
			4624 => "00000001011101110100100011010001",
			4625 => "0000000011000000000010000000010100",
			4626 => "0000000000000000000000111000001000",
			4627 => "0000000010000000001100010000000100",
			4628 => "00000000000000000100100011010001",
			4629 => "11111110011100010100100011010001",
			4630 => "0000000100000000001100111100001000",
			4631 => "0000000111000000001100101000000100",
			4632 => "00000001001101010100100011010001",
			4633 => "00000000000000000100100011010001",
			4634 => "11111111100111000100100011010001",
			4635 => "0000001101000000001111010000100000",
			4636 => "0000001100000000000100011000010000",
			4637 => "0000001111000000001111010100001000",
			4638 => "0000001000000000000110011000000100",
			4639 => "00000000000000000100100011010001",
			4640 => "11111111011111100100100011010001",
			4641 => "0000001111000000001011110000000100",
			4642 => "00000001010001010100100011010001",
			4643 => "00000000000000000100100011010001",
			4644 => "0000001100000000000100011000001000",
			4645 => "0000000101000000001101000100000100",
			4646 => "11111110110010110100100011010001",
			4647 => "00000000000000000100100011010001",
			4648 => "0000001100000000001000000000000100",
			4649 => "00000000110011000100100011010001",
			4650 => "00000000000000000100100011010001",
			4651 => "0000001100000000000111001000000100",
			4652 => "11111110101011000100100011010001",
			4653 => "0000000110000000001101011000001000",
			4654 => "0000001001000000001000010000000100",
			4655 => "11111111101010100100100011010001",
			4656 => "00000000110100010100100011010001",
			4657 => "0000000011000000001101101100000100",
			4658 => "11111111010110010100100011010001",
			4659 => "00000000001001110100100011010001",
			4660 => "0000001110000000001110101101100000",
			4661 => "0000001011000000001100101100111000",
			4662 => "0000000100000000001000000100001100",
			4663 => "0000001100000000000100000000000100",
			4664 => "00000000000000000100101010101101",
			4665 => "0000001101000000001001110100000100",
			4666 => "11111110100101000100101010101101",
			4667 => "00000000000000000100101010101101",
			4668 => "0000000011000000000100000100011100",
			4669 => "0000000100000000001111100000010000",
			4670 => "0000001011000000000101101100001000",
			4671 => "0000000110000000001011001100000100",
			4672 => "11111111011011110100101010101101",
			4673 => "00000000101001100100101010101101",
			4674 => "0000000111000000001000111100000100",
			4675 => "00000000000000000100101010101101",
			4676 => "11111110111000110100101010101101",
			4677 => "0000000101000000000100001000000100",
			4678 => "11111111110101100100101010101101",
			4679 => "0000000111000000001101100000000100",
			4680 => "00000000110001000100101010101101",
			4681 => "11111111111000100100101010101101",
			4682 => "0000001111000000001110010000001000",
			4683 => "0000001101000000001011000000000100",
			4684 => "00000000000000000100101010101101",
			4685 => "00000001010110110100101010101101",
			4686 => "0000001101000000000110100100000100",
			4687 => "11111110110110110100101010101101",
			4688 => "00000000100000000100101010101101",
			4689 => "0000000010000000000110010000010100",
			4690 => "0000000100000000001011110000001100",
			4691 => "0000001111000000000010110100000100",
			4692 => "00000000000000000100101010101101",
			4693 => "0000000000000000001000101100000100",
			4694 => "11111111101111110100101010101101",
			4695 => "00000000000000000100101010101101",
			4696 => "0000000000000000000010111100000100",
			4697 => "00000000101000010100101010101101",
			4698 => "00000000000000000100101010101101",
			4699 => "0000000110000000001000010000001100",
			4700 => "0000001100000000000100000000000100",
			4701 => "00000000000000000100101010101101",
			4702 => "0000001001000000000111101000000100",
			4703 => "11111110011100010100101010101101",
			4704 => "00000000000000000100101010101101",
			4705 => "0000000101000000001001110100000100",
			4706 => "00000000010001100100101010101101",
			4707 => "00000000000000000100101010101101",
			4708 => "0000000101000000000111100000111100",
			4709 => "0000000110000000000100111100101100",
			4710 => "0000001100000000000100001000010000",
			4711 => "0000000100000000000000010100001100",
			4712 => "0000001011000000000000001100000100",
			4713 => "00000000000000000100101010101101",
			4714 => "0000000111000000000111001000000100",
			4715 => "11111110101001010100101010101101",
			4716 => "00000000000000000100101010101101",
			4717 => "00000000010011000100101010101101",
			4718 => "0000001001000000000100101100001100",
			4719 => "0000001101000000000101110000001000",
			4720 => "0000000000000000001100000100000100",
			4721 => "00000000000000000100101010101101",
			4722 => "00000000111000010100101010101101",
			4723 => "00000000000000000100101010101101",
			4724 => "0000000100000000001011101100001000",
			4725 => "0000001011000000000000011100000100",
			4726 => "00000000000000000100101010101101",
			4727 => "11111111001110100100101010101101",
			4728 => "0000000100000000001011110000000100",
			4729 => "00000000010110110100101010101101",
			4730 => "11111111111101110100101010101101",
			4731 => "0000000000000000000011010000001000",
			4732 => "0000001001000000001101111100000100",
			4733 => "00000000000000000100101010101101",
			4734 => "00000001010110100100101010101101",
			4735 => "0000001100000000000110000100000100",
			4736 => "00000000110111110100101010101101",
			4737 => "11111111001100010100101010101101",
			4738 => "0000000101000000000010011100100000",
			4739 => "0000000111000000001000011000010000",
			4740 => "0000001000000000000001010100001000",
			4741 => "0000001100000000001001110100000100",
			4742 => "11111111100001000100101010101101",
			4743 => "00000000000000000100101010101101",
			4744 => "0000000100000000001001001100000100",
			4745 => "00000000111100000100101010101101",
			4746 => "11111111111101000100101010101101",
			4747 => "0000000011000000000010010100001100",
			4748 => "0000001011000000000110110100000100",
			4749 => "00000000000000000100101010101101",
			4750 => "0000001101000000000111111100000100",
			4751 => "00000000000000000100101010101101",
			4752 => "11111110010100000100101010101101",
			4753 => "00000000000000000100101010101101",
			4754 => "0000001110000000001000101000010100",
			4755 => "0000001101000000000011001000000100",
			4756 => "00000000000000000100101010101101",
			4757 => "0000001100000000000001101000001000",
			4758 => "0000000000000000001011010100000100",
			4759 => "00000000000000000100101010101101",
			4760 => "00000001001000110100101010101101",
			4761 => "0000000011000000000010010100000100",
			4762 => "00000000000000000100101010101101",
			4763 => "00000000000010100100101010101101",
			4764 => "0000000101000000000011001000010000",
			4765 => "0000001110000000001011110000001000",
			4766 => "0000000011000000000010010100000100",
			4767 => "00000000000000000100101010101101",
			4768 => "11111110111011100100101010101101",
			4769 => "0000000101000000001110010000000100",
			4770 => "00000000011000110100101010101101",
			4771 => "11111111100000110100101010101101",
			4772 => "0000000111000000000110110100001000",
			4773 => "0000001101000000001100000000000100",
			4774 => "00000000000000000100101010101101",
			4775 => "00000000110011110100101010101101",
			4776 => "0000001001000000001010100000000100",
			4777 => "00000000011011100100101010101101",
			4778 => "11111111100101100100101010101101",
			4779 => "0000000101000000000100001000001100",
			4780 => "0000000000000000001000011000000100",
			4781 => "11111110101000010100101111111001",
			4782 => "0000000100000000000100100100000100",
			4783 => "00000000000000000100101111111001",
			4784 => "11111111111100000100101111111001",
			4785 => "0000001111000000000010011101001000",
			4786 => "0000000110000000001101011000010100",
			4787 => "0000001110000000001011011100001000",
			4788 => "0000000110000000001001011000000100",
			4789 => "00000000000000000100101111111001",
			4790 => "11111110101110100100101111111001",
			4791 => "0000000001000000001101101000000100",
			4792 => "00000000000000000100101111111001",
			4793 => "0000001000000000000010101100000100",
			4794 => "00000000000000000100101111111001",
			4795 => "00000001001000110100101111111001",
			4796 => "0000000010000000001100010000011100",
			4797 => "0000000100000000001001001100010000",
			4798 => "0000001011000000000101101100001000",
			4799 => "0000001010000000000001010000000100",
			4800 => "00000000000000000100101111111001",
			4801 => "11111110111101000100101111111001",
			4802 => "0000000000000000000000110000000100",
			4803 => "00000000111110010100101111111001",
			4804 => "11111111110010010100101111111001",
			4805 => "0000001100000000001000111000001000",
			4806 => "0000001011000000000011011100000100",
			4807 => "00000000000000000100101111111001",
			4808 => "00000001011100100100101111111001",
			4809 => "00000000000000000100101111111001",
			4810 => "0000000110000000001111000000010000",
			4811 => "0000000001000000000010001100001000",
			4812 => "0000000010000000000111011000000100",
			4813 => "00000000000010110100101111111001",
			4814 => "00000000000000000100101111111001",
			4815 => "0000001001000000001101011100000100",
			4816 => "11111110101101100100101111111001",
			4817 => "00000000000000000100101111111001",
			4818 => "0000001100000000001000111000000100",
			4819 => "00000001000000110100101111111001",
			4820 => "11111111011011100100101111111001",
			4821 => "0000000100000000001110100100101000",
			4822 => "0000000110000000001000010000011000",
			4823 => "0000000001000000000111100100001000",
			4824 => "0000000100000000001000110100000100",
			4825 => "11111110101110110100101111111001",
			4826 => "00000000010101100100101111111001",
			4827 => "0000000101000000000001101000001000",
			4828 => "0000000000000000001000110000000100",
			4829 => "00000000000000000100101111111001",
			4830 => "00000001011010000100101111111001",
			4831 => "0000001100000000000100001000000100",
			4832 => "11111110100000110100101111111001",
			4833 => "00000000001011000100101111111001",
			4834 => "0000000000000000000001110100000100",
			4835 => "00000000000000000100101111111001",
			4836 => "0000001100000000001111011100001000",
			4837 => "0000000001000000001101011000000100",
			4838 => "00000001011001110100101111111001",
			4839 => "00000000000000000100101111111001",
			4840 => "00000000000000000100101111111001",
			4841 => "0000000110000000001000010000011000",
			4842 => "0000001011000000001100101100001100",
			4843 => "0000001101000000001001001000001000",
			4844 => "0000000100000000000010111000000100",
			4845 => "11111110110101110100101111111001",
			4846 => "00000000001001000100101111111001",
			4847 => "00000001011011010100101111111001",
			4848 => "0000001100000000001000111000000100",
			4849 => "11111110000010000100101111111001",
			4850 => "0000000001000000001011111100000100",
			4851 => "00000000011001010100101111111001",
			4852 => "11111101111101000100101111111001",
			4853 => "0000001011000000001010111100000100",
			4854 => "00000001100000100100101111111001",
			4855 => "0000000010000000001011110000001000",
			4856 => "0000000110000000001000010000000100",
			4857 => "11111110010011110100101111111001",
			4858 => "00000000101100000100101111111001",
			4859 => "0000000000000000001111000100000100",
			4860 => "00000000101000110100101111111001",
			4861 => "11111111110011010100101111111001",
			4862 => "0000000011000000001011000000001100",
			4863 => "0000000110000000001001100100000100",
			4864 => "11111110011001110100110100111101",
			4865 => "0000000111000000001000111000000100",
			4866 => "00000001010010010100110100111101",
			4867 => "11111110100100000100110100111101",
			4868 => "0000000110000000000100111101001100",
			4869 => "0000000111000000000101101100100100",
			4870 => "0000000110000000001101011000000100",
			4871 => "11111110011111110100110100111101",
			4872 => "0000000010000000000010000100010000",
			4873 => "0000000011000000000100000100001000",
			4874 => "0000000100000000001111100000000100",
			4875 => "11111111010000010100110100111101",
			4876 => "00000010011000100100110100111101",
			4877 => "0000000010000000001100010100000100",
			4878 => "11111111111111000100110100111101",
			4879 => "00000001101111110100110100111101",
			4880 => "0000000110000000001001100100001000",
			4881 => "0000001001000000001011101000000100",
			4882 => "00000001100100110100110100111101",
			4883 => "11111110010111000100110100111101",
			4884 => "0000001111000000000111111100000100",
			4885 => "00000001100001000100110100111101",
			4886 => "00000000000110100100110100111101",
			4887 => "0000001010000000001001000100011100",
			4888 => "0000001011000000000110110100010000",
			4889 => "0000001110000000001100010000001000",
			4890 => "0000001000000000001010110000000100",
			4891 => "00000000001010000100110100111101",
			4892 => "11111111000001010100110100111101",
			4893 => "0000001010000000000010101100000100",
			4894 => "00000011000010000100110100111101",
			4895 => "00000000100101100100110100111101",
			4896 => "0000001001000000000100101100001000",
			4897 => "0000001111000000001011101100000100",
			4898 => "11111110100100000100110100111101",
			4899 => "00000001010010110100110100111101",
			4900 => "11111110001111000100110100111101",
			4901 => "0000001010000000001001000100000100",
			4902 => "11111011100100000100110100111101",
			4903 => "0000001010000000001001000100000100",
			4904 => "00000001010101100100110100111101",
			4905 => "11111110001000000100110100111101",
			4906 => "0000000101000000000001000000011100",
			4907 => "0000000100000000000111011100010000",
			4908 => "0000001110000000000011001000001000",
			4909 => "0000000111000000000110000100000100",
			4910 => "00000001101100000100110100111101",
			4911 => "11111111001011010100110100111101",
			4912 => "0000001000000000000001010100000100",
			4913 => "00000000010100110100110100111101",
			4914 => "00000001101010100100110100111101",
			4915 => "0000001001000000000001000100000100",
			4916 => "00000001101110110100110100111101",
			4917 => "0000000100000000001100111100000100",
			4918 => "00000000001001010100110100111101",
			4919 => "11111110001010000100110100111101",
			4920 => "0000001111000000001000000100010100",
			4921 => "0000000111000000001000011000000100",
			4922 => "00000000110101000100110100111101",
			4923 => "0000001000000000000101000100001000",
			4924 => "0000000110000000001000010000000100",
			4925 => "11111111101100100100110100111101",
			4926 => "00000010001101010100110100111101",
			4927 => "0000001111000000001110000000000100",
			4928 => "11111110000110010100110100111101",
			4929 => "11111111010101010100110100111101",
			4930 => "0000000011000000000110001100010000",
			4931 => "0000001000000000000001010100001000",
			4932 => "0000000011000000000101000000000100",
			4933 => "00000000000101010100110100111101",
			4934 => "00000110010001000100110100111101",
			4935 => "0000000000000000000000110000000100",
			4936 => "00000001000010110100110100111101",
			4937 => "11111110011100100100110100111101",
			4938 => "0000000000000000001011000100001000",
			4939 => "0000001110000000000010110000000100",
			4940 => "11111110101110010100110100111101",
			4941 => "00000000110000000100110100111101",
			4942 => "11111110011001110100110100111101",
			4943 => "0000000110000000001101011000110100",
			4944 => "0000000000000000000110001000100100",
			4945 => "0000000000000000000101000100000100",
			4946 => "11111110011010100100111011011001",
			4947 => "0000001011000000000101100100010000",
			4948 => "0000001100000000001011000000001100",
			4949 => "0000001100000000001110001100000100",
			4950 => "11111110101100100100111011011001",
			4951 => "0000001101000000001110101100000100",
			4952 => "00000011001011100100111011011001",
			4953 => "00000000010101000100111011011001",
			4954 => "00000101101111010100111011011001",
			4955 => "0000000010000000001000001100001000",
			4956 => "0000001101000000001111010000000100",
			4957 => "00000000000000000100111011011001",
			4958 => "11111110011011100100111011011001",
			4959 => "0000001011000000001011110100000100",
			4960 => "00000011001011000100111011011001",
			4961 => "11111110100101000100111011011001",
			4962 => "0000000011000000001010001100000100",
			4963 => "11111110011000100100111011011001",
			4964 => "0000001111000000001111010000001000",
			4965 => "0000001111000000000111100000000100",
			4966 => "11111110000111100100111011011001",
			4967 => "00000001010101100100111011011001",
			4968 => "11111110011000100100111011011001",
			4969 => "0000001100000000001000011001110100",
			4970 => "0000000110000000001111000001000000",
			4971 => "0000000010000000001100000000100000",
			4972 => "0000001011000000001100101100010000",
			4973 => "0000000011000000000001101000001000",
			4974 => "0000000100000000001111100000000100",
			4975 => "11111110001100000100111011011001",
			4976 => "00000001101001000100111011011001",
			4977 => "0000001101000000000100011000000100",
			4978 => "11111111011000000100111011011001",
			4979 => "00000001111100110100111011011001",
			4980 => "0000000100000000000010010100001000",
			4981 => "0000000110000000001001100100000100",
			4982 => "11111110100100010100111011011001",
			4983 => "00000010001111010100111011011001",
			4984 => "0000000000000000000010011000000100",
			4985 => "11111100100001100100111011011001",
			4986 => "11111111111000000100111011011001",
			4987 => "0000000011000000001100010000010000",
			4988 => "0000001100000000001000111100001000",
			4989 => "0000000010000000001010000100000100",
			4990 => "00000000101101010100111011011001",
			4991 => "11111101111110010100111011011001",
			4992 => "0000001111000000000110100000000100",
			4993 => "00000000000000000100111011011001",
			4994 => "11111110001001000100111011011001",
			4995 => "0000001111000000001010000100001000",
			4996 => "0000001110000000000010000100000100",
			4997 => "00000000100111110100111011011001",
			4998 => "00000100100101010100111011011001",
			4999 => "0000000000000000001011010100000100",
			5000 => "11111110010110010100111011011001",
			5001 => "00000000010101000100111011011001",
			5002 => "0000001000000000000001110000011000",
			5003 => "0000000111000000001000011000001100",
			5004 => "0000000100000000001000011100001000",
			5005 => "0000000000000000000111000100000100",
			5006 => "11111110111101000100111011011001",
			5007 => "00000001111100110100111011011001",
			5008 => "11111111100100010100111011011001",
			5009 => "0000000101000000000001000000000100",
			5010 => "00000001001111000100111011011001",
			5011 => "0000001011000000001010010100000100",
			5012 => "11111101111101100100111011011001",
			5013 => "00000000000111100100111011011001",
			5014 => "0000001110000000000001011100010000",
			5015 => "0000000111000000000110000100001000",
			5016 => "0000001101000000001011000000000100",
			5017 => "00000000110010000100111011011001",
			5018 => "00000010000010000100111011011001",
			5019 => "0000000011000000001110010000000100",
			5020 => "11111111001001110100111011011001",
			5021 => "00000001000010010100111011011001",
			5022 => "0000000110000000001000010000000100",
			5023 => "00000100001001010100111011011001",
			5024 => "0000001011000000001011110100000100",
			5025 => "00000001110101100100111011011001",
			5026 => "00000000101101100100111011011001",
			5027 => "0000001101000000000110111100010000",
			5028 => "0000001100000000000001011000001000",
			5029 => "0000000110000000001111000000000100",
			5030 => "00000000000000000100111011011001",
			5031 => "11111110011001110100111011011001",
			5032 => "0000000011000000001000110100000100",
			5033 => "00000011100111010100111011011001",
			5034 => "11111111011010100100111011011001",
			5035 => "0000000000000000000111000000001000",
			5036 => "0000001110000000001110000000000100",
			5037 => "11111111010010110100111011011001",
			5038 => "00010001100000100100111011011001",
			5039 => "0000000000000000001011000100001100",
			5040 => "0000000100000000001010110100000100",
			5041 => "11111110011100110100111011011001",
			5042 => "0000001010000000000001010000000100",
			5043 => "00000011011010000100111011011001",
			5044 => "00000000011101010100111011011001",
			5045 => "11111110011000100100111011011001",
			5046 => "0000000110000000001101011000111100",
			5047 => "0000001001000000000101010000100000",
			5048 => "0000000001000000000111100100001100",
			5049 => "0000000011000000001010001100000100",
			5050 => "11111110011000110101000001110101",
			5051 => "0000000011000000000100000100000100",
			5052 => "00000000100100010101000001110101",
			5053 => "11111110011111010101000001110101",
			5054 => "0000000111000000000011100000010000",
			5055 => "0000001100000000001110001100000100",
			5056 => "11111110100010010101000001110101",
			5057 => "0000000000000000000001110000000100",
			5058 => "11111110101111100101000001110101",
			5059 => "0000000000000000001101010000000100",
			5060 => "00000011000101100101000001110101",
			5061 => "11111111100100000101000001110101",
			5062 => "11111110010111010101000001110101",
			5063 => "0000001010000000001010100100001000",
			5064 => "0000001011000000000101100100000100",
			5065 => "00000100100111110101000001110101",
			5066 => "11111111100001110101000001110101",
			5067 => "0000001011000000000000011100000100",
			5068 => "11111110100010010101000001110101",
			5069 => "0000000001000000001110010100001100",
			5070 => "0000000111000000000110100100000100",
			5071 => "00000001100001000101000001110101",
			5072 => "0000000001000000000001000100000100",
			5073 => "00000000111100110101000001110101",
			5074 => "11111110011110110101000001110101",
			5075 => "00000010101101010101000001110101",
			5076 => "0000001011000000000000110101101000",
			5077 => "0000000110000000001111000000111000",
			5078 => "0000001011000000001100101100011000",
			5079 => "0000001111000000001110010000010000",
			5080 => "0000000011000000000001011000001000",
			5081 => "0000001111000000001001010000000100",
			5082 => "00000001000000110101000001110101",
			5083 => "11111110001001000101000001110101",
			5084 => "0000000100000000001000000100000100",
			5085 => "00000001011110100101000001110101",
			5086 => "00000010010000100101000001110101",
			5087 => "0000000011000000000111110000000100",
			5088 => "11111101110000000101000001110101",
			5089 => "00000000110000010101000001110101",
			5090 => "0000000100000000000110111000010000",
			5091 => "0000001010000000001000100100001000",
			5092 => "0000001111000000001010000100000100",
			5093 => "00000001010011100101000001110101",
			5094 => "11111111010011110101000001110101",
			5095 => "0000000001000000001101101000000100",
			5096 => "00000001000001100101000001110101",
			5097 => "00000011010100110101000001110101",
			5098 => "0000001011000000001010001100001000",
			5099 => "0000000000000000001111000100000100",
			5100 => "11111101100000100101000001110101",
			5101 => "11111111001111110101000001110101",
			5102 => "0000000001000000000111101000000100",
			5103 => "00000001011010110101000001110101",
			5104 => "11111110110011100101000001110101",
			5105 => "0000001110000000000110111000100000",
			5106 => "0000000101000000000001000000010000",
			5107 => "0000001110000000001111100100001000",
			5108 => "0000000111000000000110000100000100",
			5109 => "00000001110000010101000001110101",
			5110 => "00000000010100100101000001110101",
			5111 => "0000001001000000000010101100000100",
			5112 => "00000001110100000101000001110101",
			5113 => "00000000110001000101000001110101",
			5114 => "0000000111000000001000011000001000",
			5115 => "0000000100000000001011110000000100",
			5116 => "00000000001000010101000001110101",
			5117 => "00000001100011000101000001110101",
			5118 => "0000000011000000001111101000000100",
			5119 => "11111110010001000101000001110101",
			5120 => "00000000000100100101000001110101",
			5121 => "0000000110000000001000010000000100",
			5122 => "00000111100101100101000001110101",
			5123 => "0000000101000000000011001000001000",
			5124 => "0000001100000000001001110100000100",
			5125 => "00000001110100010101000001110101",
			5126 => "00000000010101000101000001110101",
			5127 => "11111110100111000101000001110101",
			5128 => "0000000000000000001011000100101000",
			5129 => "0000001001000000001010100000010100",
			5130 => "0000000110000000001001111100001100",
			5131 => "0000001001000000000000001000001000",
			5132 => "0000000101000000000110010000000100",
			5133 => "00000000000000000101000001110101",
			5134 => "00000010010110100101000001110101",
			5135 => "00000100110011110101000001110101",
			5136 => "0000000001000000000111101000000100",
			5137 => "00000001010110010101000001110101",
			5138 => "11111110101101000101000001110101",
			5139 => "0000000100000000001011100000010000",
			5140 => "0000001011000000000110100000001000",
			5141 => "0000001100000000000100000100000100",
			5142 => "11111110011001000101000001110101",
			5143 => "00000000011100110101000001110101",
			5144 => "0000000000000000001010101100000100",
			5145 => "00000101011100100101000001110101",
			5146 => "11111110011101000101000001110101",
			5147 => "00000001100011000101000001110101",
			5148 => "11111110011001000101000001110101",
			5149 => "0000000100000000000011000001000000",
			5150 => "0000001100000000000100011000100100",
			5151 => "0000000111000000000110100100011000",
			5152 => "0000000001000000001101101000000100",
			5153 => "00000000000000000101001000001001",
			5154 => "0000000001000000001110010100001100",
			5155 => "0000001000000000000010101100000100",
			5156 => "00000000000000000101001000001001",
			5157 => "0000001100000000000100011000000100",
			5158 => "00000000101100000101001000001001",
			5159 => "00000000000000000101001000001001",
			5160 => "0000001110000000001100010000000100",
			5161 => "11111111110101110101001000001001",
			5162 => "00000000000000000101001000001001",
			5163 => "0000000010000000000000010000000100",
			5164 => "11111111001110110101001000001001",
			5165 => "0000001000000000001100011100000100",
			5166 => "00000000001111010101001000001001",
			5167 => "00000000000000000101001000001001",
			5168 => "0000000111000000001000011000011000",
			5169 => "0000001000000000001010110000010000",
			5170 => "0000000100000000001100010000000100",
			5171 => "00000000000000000101001000001001",
			5172 => "0000001011000000001011011100001000",
			5173 => "0000000000000000000101000100000100",
			5174 => "00000000000000000101001000001001",
			5175 => "00000000111001010101001000001001",
			5176 => "00000000000000000101001000001001",
			5177 => "0000001000000000000110011100000100",
			5178 => "11111111111001010101001000001001",
			5179 => "00000000000100010101001000001001",
			5180 => "00000000000000000101001000001001",
			5181 => "0000000000000000000000111000111100",
			5182 => "0000001000000000000111000100111000",
			5183 => "0000000011000000001111101000011100",
			5184 => "0000001100000000001001110000010000",
			5185 => "0000000001000000000110101000001000",
			5186 => "0000001011000000001100101100000100",
			5187 => "00000000000000000101001000001001",
			5188 => "11111110110000010101001000001001",
			5189 => "0000000000000000000011010000000100",
			5190 => "00000000101111010101001000001001",
			5191 => "11111111110000000101001000001001",
			5192 => "0000000001000000001001011000000100",
			5193 => "11111110100110000101001000001001",
			5194 => "0000000111000000001000011000000100",
			5195 => "00000000000101100101001000001001",
			5196 => "11111111001000100101001000001001",
			5197 => "0000000001000000000100110100001100",
			5198 => "0000001100000000000100011000000100",
			5199 => "00000000000000000101001000001001",
			5200 => "0000001010000000001010110000000100",
			5201 => "00000000110000000101001000001001",
			5202 => "00000000000000000101001000001001",
			5203 => "0000001010000000001000010100001000",
			5204 => "0000001100000000001010001100000100",
			5205 => "00000000100011110101001000001001",
			5206 => "00000000000000000101001000001001",
			5207 => "0000001100000000001001110100000100",
			5208 => "00000000000000000101001000001001",
			5209 => "11111111001110100101001000001001",
			5210 => "11111110111011100101001000001001",
			5211 => "0000000000000000001010000000100000",
			5212 => "0000000101000000001110110100011100",
			5213 => "0000000100000000001101001000010000",
			5214 => "0000000000000000000000111000001000",
			5215 => "0000001000000000001111001000000100",
			5216 => "00000000000000000101001000001001",
			5217 => "00000000010101000101001000001001",
			5218 => "0000000000000000000000110000000100",
			5219 => "11111111011100110101001000001001",
			5220 => "00000000000000000101001000001001",
			5221 => "0000001001000000001111001100000100",
			5222 => "00000000000000000101001000001001",
			5223 => "0000001100000000001000000000000100",
			5224 => "00000001011000100101001000001001",
			5225 => "00000000000000000101001000001001",
			5226 => "11111111011111010101001000001001",
			5227 => "0000001010000000000101000100010100",
			5228 => "0000000001000000001001111000001100",
			5229 => "0000000101000000000111001000000100",
			5230 => "11111111101111110101001000001001",
			5231 => "0000000010000000001100010000000100",
			5232 => "00000000101011010101001000001001",
			5233 => "00000000000000000101001000001001",
			5234 => "0000000100000000001010110100000100",
			5235 => "00000000000000000101001000001001",
			5236 => "11111110111110100101001000001001",
			5237 => "0000001000000000001111000100010000",
			5238 => "0000001100000000000011011100001000",
			5239 => "0000000001000000001001111000000100",
			5240 => "00000000000000000101001000001001",
			5241 => "00000001000100000101001000001001",
			5242 => "0000000011000000000101010100000100",
			5243 => "11111111100010110101001000001001",
			5244 => "00000000100000110101001000001001",
			5245 => "0000000100000000000001001100000100",
			5246 => "11111111000000110101001000001001",
			5247 => "0000000101000000000000001100000100",
			5248 => "00000000000000000101001000001001",
			5249 => "00000000001101000101001000001001",
			5250 => "0000000110000000001101011000110100",
			5251 => "0000000001000000000101011100010100",
			5252 => "0000000110000000001001011000001000",
			5253 => "0000000000000000001100000100000100",
			5254 => "11111111110010110101001111011111",
			5255 => "00000000010110010101001111011111",
			5256 => "0000000100000000000101110000001000",
			5257 => "0000001000000000000010101100000100",
			5258 => "11111111001001100101001111011111",
			5259 => "00000000101101000101001111011111",
			5260 => "11111110011010100101001111011111",
			5261 => "0000000011000000001010000100011000",
			5262 => "0000001100000000001011000000010000",
			5263 => "0000000100000000000111010100000100",
			5264 => "11111110110000110101001111011111",
			5265 => "0000001010000000000010101100000100",
			5266 => "00000001110011000101001111011111",
			5267 => "0000001110000000001001011100000100",
			5268 => "00000000011001100101001111011111",
			5269 => "11111111001011100101001111011111",
			5270 => "0000001001000000000101010000000100",
			5271 => "11111111111001100101001111011111",
			5272 => "00000010101011100101001111011111",
			5273 => "0000000001000000000101011100000100",
			5274 => "00000000011000110101001111011111",
			5275 => "11111110011000110101001111011111",
			5276 => "0000000110000000001000010001110000",
			5277 => "0000001111000000001001011100111100",
			5278 => "0000000011000000001000011000011100",
			5279 => "0000001100000000000000101000001100",
			5280 => "0000000111000000000100000000000100",
			5281 => "11111110101100000101001111011111",
			5282 => "0000000100000000001110111000000100",
			5283 => "11111111101100100101001111011111",
			5284 => "00000010001000000101001111011111",
			5285 => "0000001110000000000111001000001000",
			5286 => "0000001101000000001110110000000100",
			5287 => "11111110100101100101001111011111",
			5288 => "00000000100010110101001111011111",
			5289 => "0000001110000000001011000000000100",
			5290 => "11111101101000010101001111011111",
			5291 => "11111111010101010101001111011111",
			5292 => "0000000000000000000011111100010000",
			5293 => "0000000011000000000000011100001000",
			5294 => "0000000000000000000010111100000100",
			5295 => "11111110110000110101001111011111",
			5296 => "11111100111010010101001111011111",
			5297 => "0000001100000000000100000000000100",
			5298 => "00000010001011010101001111011111",
			5299 => "11111111110110010101001111011111",
			5300 => "0000000111000000001001110000001000",
			5301 => "0000001111000000000001000000000100",
			5302 => "00000010101101010101001111011111",
			5303 => "00000001100011010101001111011111",
			5304 => "0000000110000000001001100100000100",
			5305 => "11111110110110100101001111011111",
			5306 => "00000001100010010101001111011111",
			5307 => "0000000100000000001100001100010100",
			5308 => "0000000000000000000010111100010000",
			5309 => "0000000001000000001101101000001000",
			5310 => "0000001110000000001001010100000100",
			5311 => "11111011011001010101001111011111",
			5312 => "11111110010101110101001111011111",
			5313 => "0000000101000000000001101000000100",
			5314 => "00000001100101010101001111011111",
			5315 => "11111111111000010101001111011111",
			5316 => "00000001101010010101001111011111",
			5317 => "0000000100000000000010111000010000",
			5318 => "0000000110000000000100111100001000",
			5319 => "0000000000000000000011111100000100",
			5320 => "11111101101001110101001111011111",
			5321 => "11111111111101100101001111011111",
			5322 => "0000001111000000001000011100000100",
			5323 => "11111011011010100101001111011111",
			5324 => "11111111100111110101001111011111",
			5325 => "0000000110000000001001100100001000",
			5326 => "0000000000000000001111000100000100",
			5327 => "00000000001111110101001111011111",
			5328 => "11111110001011000101001111011111",
			5329 => "0000001001000000000000111100000100",
			5330 => "11111110111010010101001111011111",
			5331 => "00000000100111000101001111011111",
			5332 => "0000001101000000001010001000100000",
			5333 => "0000001000000000000110001000001100",
			5334 => "0000000000000000001010101100000100",
			5335 => "11111111001111010101001111011111",
			5336 => "0000000100000000001001001100000100",
			5337 => "00000001101010000101001111011111",
			5338 => "00000000000000000101001111011111",
			5339 => "0000000111000000000110000100001000",
			5340 => "0000001001000000001100011000000100",
			5341 => "00000001110101110101001111011111",
			5342 => "00000000011110000101001111011111",
			5343 => "0000001001000000001010011000000100",
			5344 => "11111101010110110101001111011111",
			5345 => "0000000111000000001110110000000100",
			5346 => "00000001101001100101001111011111",
			5347 => "11111111001111110101001111011111",
			5348 => "0000001111000000001000000100001100",
			5349 => "0000001111000000000110111000001000",
			5350 => "0000001111000000000010010100000100",
			5351 => "11111111101110010101001111011111",
			5352 => "00000000011101010101001111011111",
			5353 => "11111110010100100101001111011111",
			5354 => "0000000000000000000111000000001100",
			5355 => "0000001111000000001000110100000100",
			5356 => "11111111101001110101001111011111",
			5357 => "0000000111000000000100010000000100",
			5358 => "00000010101100010101001111011111",
			5359 => "00000000010000010101001111011111",
			5360 => "0000000011000000001000000100001000",
			5361 => "0000000011000000001011110000000100",
			5362 => "11111111001101000101001111011111",
			5363 => "00000001110000110101001111011111",
			5364 => "0000001101000000001110110100000100",
			5365 => "00000001000111000101001111011111",
			5366 => "11111111010001010101001111011111",
			5367 => "0000000011000000001001110100100100",
			5368 => "0000001010000000000001010100001000",
			5369 => "0000001011000000000100001000000100",
			5370 => "11111110011100000101010011000001",
			5371 => "00000000000000000101010011000001",
			5372 => "0000001010000000001001101000001100",
			5373 => "0000000101000000001010111100000100",
			5374 => "11111111011111000101010011000001",
			5375 => "0000000110000000001001100100000100",
			5376 => "00000000000000000101010011000001",
			5377 => "00000001001101110101010011000001",
			5378 => "0000000010000000000000010000000100",
			5379 => "11111110100000100101010011000001",
			5380 => "0000000010000000000110101100001000",
			5381 => "0000001110000000000111000000000100",
			5382 => "00000000000000000101010011000001",
			5383 => "00000000101100010101010011000001",
			5384 => "00000000000000000101010011000001",
			5385 => "0000001111000000001100100100011000",
			5386 => "0000001001000000001111001100001000",
			5387 => "0000001000000000000111000100000100",
			5388 => "00000000000000000101010011000001",
			5389 => "00000010001000110101010011000001",
			5390 => "0000000011000000000001101000000100",
			5391 => "11111110101011000101010011000001",
			5392 => "0000000000000000000110011000000100",
			5393 => "00000000000000000101010011000001",
			5394 => "0000000111000000001000111000000100",
			5395 => "00000000000000000101010011000001",
			5396 => "00000001011101010101010011000001",
			5397 => "0000000101000000001010111000010000",
			5398 => "0000001111000000001111010000001100",
			5399 => "0000000011000000001010011100001000",
			5400 => "0000001110000000001000000000000100",
			5401 => "11111110100101000101010011000001",
			5402 => "00000000000000000101010011000001",
			5403 => "00000001001100000101010011000001",
			5404 => "11111110001011010101010011000001",
			5405 => "0000000111000000001000111000001100",
			5406 => "0000000000000000000010011000000100",
			5407 => "11111110110111110101010011000001",
			5408 => "0000001101000000001011000000000100",
			5409 => "00000000000000000101010011000001",
			5410 => "00000001111011110101010011000001",
			5411 => "0000001101000000001000000000010000",
			5412 => "0000000000000000000000110000001000",
			5413 => "0000000010000000001001100000000100",
			5414 => "00000000000000000101010011000001",
			5415 => "11111101001010110101010011000001",
			5416 => "0000001010000000000110011100000100",
			5417 => "11111111001101110101010011000001",
			5418 => "00000000011000100101010011000001",
			5419 => "0000001000000000001111000100001000",
			5420 => "0000000101000000001000000000000100",
			5421 => "00000000101110110101010011000001",
			5422 => "00000000000100010101010011000001",
			5423 => "11111110010011100101010011000001",
			5424 => "0000000011000000001001110100100100",
			5425 => "0000000100000000000010010000001000",
			5426 => "0000001101000000001000011000000100",
			5427 => "11111110100000100101010111000101",
			5428 => "00000000000000000101010111000101",
			5429 => "0000000011000000000100001000010000",
			5430 => "0000000010000000000000010000000100",
			5431 => "11111110101111110101010111000101",
			5432 => "0000000010000000000000010000001000",
			5433 => "0000001011000000000011100000000100",
			5434 => "00000000010100110101010111000101",
			5435 => "00000000000000000101010111000101",
			5436 => "00000000000000000101010111000101",
			5437 => "0000000100000000000101001100001000",
			5438 => "0000000111000000001101100000000100",
			5439 => "00000001000100000101010111000101",
			5440 => "00000000000000000101010111000101",
			5441 => "00000000000000000101010111000101",
			5442 => "0000001111000000001100100100011100",
			5443 => "0000000001000000001001111000001000",
			5444 => "0000001000000000000111000100000100",
			5445 => "00000000000000000101010111000101",
			5446 => "00000010000110000101010111000101",
			5447 => "0000001101000000001011000000000100",
			5448 => "11111110110100010101010111000101",
			5449 => "0000001111000000000000110100000100",
			5450 => "00000000000000000101010111000101",
			5451 => "0000001100000000000100000000000100",
			5452 => "00000000000000000101010111000101",
			5453 => "0000001110000000001000000000000100",
			5454 => "00000000000010000101010111000101",
			5455 => "00000001100101010101010111000101",
			5456 => "0000001101000000001011000000010000",
			5457 => "0000001111000000001111010000001000",
			5458 => "0000000110000000001011001100000100",
			5459 => "11111110101000100101010111000101",
			5460 => "00000000100010010101010111000101",
			5461 => "0000000011000000000000011100000100",
			5462 => "11111101110111000101010111000101",
			5463 => "11111111101011100101010111000101",
			5464 => "0000001111000000000101110000011000",
			5465 => "0000000111000000001001110000001000",
			5466 => "0000000011000000000100000100000100",
			5467 => "00000000011100000101010111000101",
			5468 => "00000010000110000101010111000101",
			5469 => "0000000011000000000010001000001000",
			5470 => "0000001000000000000001110100000100",
			5471 => "11111110100111100101010111000101",
			5472 => "00000000111100100101010111000101",
			5473 => "0000000110000000001010011000000100",
			5474 => "00000000000000000101010111000101",
			5475 => "00000001011011000101010111000101",
			5476 => "0000000001000000000111100100010000",
			5477 => "0000000000000000000010011000001000",
			5478 => "0000001101000000000110100100000100",
			5479 => "11111101011000000101010111000101",
			5480 => "11111111000001010101010111000101",
			5481 => "0000001111000000001001100000000100",
			5482 => "00000000010010000101010111000101",
			5483 => "11111110001000000101010111000101",
			5484 => "0000001011000000000000001100000100",
			5485 => "00000001100011010101010111000101",
			5486 => "0000000001000000000000111100000100",
			5487 => "11111111010100010101010111000101",
			5488 => "00000000010000110101010111000101",
			5489 => "0000000111000000001001110000110100",
			5490 => "0000001110000000000100000100101000",
			5491 => "0000000011000000000000011100100000",
			5492 => "0000000100000000000100001100001000",
			5493 => "0000001101000000001011000000000100",
			5494 => "11111110110111010101011011001001",
			5495 => "00000000000000000101011011001001",
			5496 => "0000000010000000001100010000010000",
			5497 => "0000001011000000000011011100001000",
			5498 => "0000000010000000000010000100000100",
			5499 => "11111111101110110101011011001001",
			5500 => "00000000000000000101011011001001",
			5501 => "0000001100000000000100000000000100",
			5502 => "00000001010010000101011011001001",
			5503 => "00000000000000000101011011001001",
			5504 => "0000000110000000001111000000000100",
			5505 => "11111110111110100101011011001001",
			5506 => "00000000000000000101011011001001",
			5507 => "0000001001000000001001011000000100",
			5508 => "00000000000000000101011011001001",
			5509 => "00000001010111010101011011001001",
			5510 => "0000000011000000000101110100001000",
			5511 => "0000000110000000001001100100000100",
			5512 => "00000000000000000101011011001001",
			5513 => "11111110001101000101011011001001",
			5514 => "00000000111101110101011011001001",
			5515 => "0000000111000000001001110000010100",
			5516 => "0000001100000000001000111100001100",
			5517 => "0000000110000000001101011000000100",
			5518 => "00000000000000000101011011001001",
			5519 => "0000001101000000001110110000000100",
			5520 => "00000000000000000101011011001001",
			5521 => "00000001100011010101011011001001",
			5522 => "0000000111000000001001110000000100",
			5523 => "11111111011101100101011011001001",
			5524 => "00000000100001100101011011001001",
			5525 => "0000001101000000001000000000001000",
			5526 => "0000000100000000000010010000000100",
			5527 => "11111110101011000101011011001001",
			5528 => "00000000000000000101011011001001",
			5529 => "0000001011000000000000001100011000",
			5530 => "0000000110000000001001100100001000",
			5531 => "0000001001000000001101011100000100",
			5532 => "00000000000000000101011011001001",
			5533 => "11111110100100110101011011001001",
			5534 => "0000000000000000000011111100001000",
			5535 => "0000000001000000000111100100000100",
			5536 => "11111111100101110101011011001001",
			5537 => "00000001001011010101011011001001",
			5538 => "0000000111000000000110000100000100",
			5539 => "00000001101010000101011011001001",
			5540 => "00000000000000000101011011001001",
			5541 => "0000000111000000001110001100001100",
			5542 => "0000000110000000001000010000001000",
			5543 => "0000000111000000001101100000000100",
			5544 => "00000000000000000101011011001001",
			5545 => "11111110011010110101011011001001",
			5546 => "00000000001011010101011011001001",
			5547 => "0000000000000000000010011000001000",
			5548 => "0000000011000000001010000100000100",
			5549 => "00000000100011000101011011001001",
			5550 => "00000000000011100101011011001001",
			5551 => "0000001010000000001010110000000100",
			5552 => "11111110011010000101011011001001",
			5553 => "00000000000000000101011011001001",
			5554 => "0000000011000000001001110100011000",
			5555 => "0000001010000000000001010100001000",
			5556 => "0000000001000000000111100100000100",
			5557 => "11111110011011010101011110010101",
			5558 => "00000000000000000101011110010101",
			5559 => "0000000111000000001101100000001100",
			5560 => "0000001011000000001001110000001000",
			5561 => "0000001011000000000100000000000100",
			5562 => "11111110101011100101011110010101",
			5563 => "00000000000000000101011110010101",
			5564 => "00000001011010100101011110010101",
			5565 => "11111110010101110101011110010101",
			5566 => "0000000000000000001001110001001100",
			5567 => "0000000000000000000011010000011100",
			5568 => "0000000011000000000000011100001000",
			5569 => "0000000000000000000011111100000100",
			5570 => "11111110010111110101011110010101",
			5571 => "11111011010001010101011110010101",
			5572 => "0000000101000000000100011000000100",
			5573 => "00000010010111100101011110010101",
			5574 => "0000000001000000000111100100001000",
			5575 => "0000000001000000000111100100000100",
			5576 => "11111111101101000101011110010101",
			5577 => "11111011110111010101011110010101",
			5578 => "0000000101000000000001101000000100",
			5579 => "00000001011111010101011110010101",
			5580 => "00000000000111000101011110010101",
			5581 => "0000000000000000001110111100010000",
			5582 => "0000001010000000001010110000000100",
			5583 => "11111110110001010101011110010101",
			5584 => "0000001100000000001111011100001000",
			5585 => "0000001001000000000000111100000100",
			5586 => "00000000100111000101011110010101",
			5587 => "00000001011010010101011110010101",
			5588 => "11111110110111110101011110010101",
			5589 => "0000001010000000000101000100010000",
			5590 => "0000001111000000001001011100001000",
			5591 => "0000001010000000000110011100000100",
			5592 => "11111110100111010101011110010101",
			5593 => "00000000101101100101011110010101",
			5594 => "0000000000000000000111111000000100",
			5595 => "00000000000011010101011110010101",
			5596 => "11111110010000000101011110010101",
			5597 => "0000001100000000000110000100001000",
			5598 => "0000000100000000000010010000000100",
			5599 => "00000001011011100101011110010101",
			5600 => "11111111110010010101011110010101",
			5601 => "0000001011000000001110101000000100",
			5602 => "11111110011100010101011110010101",
			5603 => "00000001010010100101011110010101",
			5604 => "11111110000101100101011110010101",
			5605 => "0000000011000000001001110100011100",
			5606 => "0000000110000000001011001100001000",
			5607 => "0000000001000000000111100100000100",
			5608 => "11111110011110010101100010101001",
			5609 => "00000000000000000101100010101001",
			5610 => "0000001110000000000001111100010000",
			5611 => "0000000011000000001101010100001000",
			5612 => "0000000010000000000111011000000100",
			5613 => "11111110111100100101100010101001",
			5614 => "00000000000000000101100010101001",
			5615 => "0000001011000000000101101100000100",
			5616 => "00000001010010100101100010101001",
			5617 => "00000000000000000101100010101001",
			5618 => "11111110001111110101100010101001",
			5619 => "0000001111000000000101110000110100",
			5620 => "0000000111000000001001110000011100",
			5621 => "0000001101000000000100011000001100",
			5622 => "0000001111000000001110101000001000",
			5623 => "0000000100000000001000000100000100",
			5624 => "00000000000000000101100010101001",
			5625 => "00000000111111000101100010101001",
			5626 => "11111110111100010101100010101001",
			5627 => "0000000010000000001100010100000100",
			5628 => "11111111010000110101100010101001",
			5629 => "0000001110000000001110110000000100",
			5630 => "00000000000110010101100010101001",
			5631 => "0000000110000000001101011000000100",
			5632 => "00000000000000000101100010101001",
			5633 => "00000001100101100101100010101001",
			5634 => "0000000011000000000100000100001000",
			5635 => "0000000100000000001011100000000100",
			5636 => "11111110100110110101100010101001",
			5637 => "00000000000000000101100010101001",
			5638 => "0000000101000000000110110100001100",
			5639 => "0000001111000000000010011100001000",
			5640 => "0000001111000000000000110100000100",
			5641 => "00000000000000000101100010101001",
			5642 => "00000001000111100101100010101001",
			5643 => "00000000000000000101100010101001",
			5644 => "11111111000011010101100010101001",
			5645 => "0000000011000000000001001000100000",
			5646 => "0000001110000000000111110000011100",
			5647 => "0000000111000000001001110000001100",
			5648 => "0000000011000000000101110100001000",
			5649 => "0000000100000000000010111000000100",
			5650 => "11111101110111010101100010101001",
			5651 => "11111111011111000101100010101001",
			5652 => "00000001001001010101100010101001",
			5653 => "0000001100000000001000111000001000",
			5654 => "0000000110000000001001100100000100",
			5655 => "11111111101111010101100010101001",
			5656 => "00000001101000110101100010101001",
			5657 => "0000000110000000001111000000000100",
			5658 => "11111111000001010101100010101001",
			5659 => "00000001000010010101100010101001",
			5660 => "11111101110011110101100010101001",
			5661 => "0000001101000000001101101100011000",
			5662 => "0000001011000000000000001100001000",
			5663 => "0000000110000000001111000000000100",
			5664 => "00000000000000000101100010101001",
			5665 => "00000001100100100101100010101001",
			5666 => "0000000011000000001001011100001000",
			5667 => "0000000101000000000001101000000100",
			5668 => "00000000001011000101100010101001",
			5669 => "11111110110011100101100010101001",
			5670 => "0000000111000000000100001000000100",
			5671 => "00000001110101000101100010101001",
			5672 => "00000000010000100101100010101001",
			5673 => "11111110011000100101100010101001",
			5674 => "0000000110000000001101011000101100",
			5675 => "0000000001000000000001000100010100",
			5676 => "0000001000000000001001000100010000",
			5677 => "0000000101000000000110110100001100",
			5678 => "0000000111000000001100101000000100",
			5679 => "11111110110001010101100110100101",
			5680 => "0000001000000000000000001000000100",
			5681 => "00000000000000000101100110100101",
			5682 => "00000001110101100101100110100101",
			5683 => "11111110011111100101100110100101",
			5684 => "11111110011001100101100110100101",
			5685 => "0000000011000000001010000100010100",
			5686 => "0000000010000000000110111100010000",
			5687 => "0000000001000000000111101000001100",
			5688 => "0000001010000000001010100000000100",
			5689 => "00000001000001100101100110100101",
			5690 => "0000001101000000000101001000000100",
			5691 => "00000000010000100101100110100101",
			5692 => "11111110101100100101100110100101",
			5693 => "00000001111001100101100110100101",
			5694 => "00000011001110000101100110100101",
			5695 => "11111110111101000101100110100101",
			5696 => "0000001010000000001011010101001100",
			5697 => "0000000110000000001000010000101100",
			5698 => "0000000100000000000010010100011000",
			5699 => "0000001100000000001000000000001100",
			5700 => "0000001001000000001011111100000100",
			5701 => "11111110110111100101100110100101",
			5702 => "0000001001000000001001111100000100",
			5703 => "00000001110111000101100110100101",
			5704 => "00000000101000100101100110100101",
			5705 => "0000001000000000000001010000001000",
			5706 => "0000000010000000000111010100000100",
			5707 => "11111111111010010101100110100101",
			5708 => "00000001111010110101100110100101",
			5709 => "11111110011011100101100110100101",
			5710 => "0000000110000000001011001100000100",
			5711 => "11111110010110110101100110100101",
			5712 => "0000001111000000001001010000001000",
			5713 => "0000000111000000001101100000000100",
			5714 => "00000001000011000101100110100101",
			5715 => "11111101111011110101100110100101",
			5716 => "0000000011000000000001011000000100",
			5717 => "11111110011000100101100110100101",
			5718 => "00000000000110010101100110100101",
			5719 => "0000000111000000001111011100010000",
			5720 => "0000000100000000000111011100001100",
			5721 => "0000001001000000001010011000000100",
			5722 => "00000000001101000101100110100101",
			5723 => "0000001000000000001100000100000100",
			5724 => "00000000011101000101100110100101",
			5725 => "00000001100111100101100110100101",
			5726 => "00000000000000000101100110100101",
			5727 => "0000001110000000000011010100001100",
			5728 => "0000001001000000000111110100001000",
			5729 => "0000001111000000000110001100000100",
			5730 => "11111111001000100101100110100101",
			5731 => "00000001000000010101100110100101",
			5732 => "11111110001101010101100110100101",
			5733 => "00000001011110010101100110100101",
			5734 => "0000000101000000000100011000000100",
			5735 => "00000000011011000101100110100101",
			5736 => "11111110010001010101100110100101",
			5737 => "0000000111000000001001110000101100",
			5738 => "0000000110000000001001100100100000",
			5739 => "0000001110000000000100000100011000",
			5740 => "0000001101000000000100011000000100",
			5741 => "11111111010100110101101011011001",
			5742 => "0000001100000000000100000000001000",
			5743 => "0000000110000000001001100100000100",
			5744 => "11111111100111010101101011011001",
			5745 => "00000000000000000101101011011001",
			5746 => "0000000010000000001100010000001000",
			5747 => "0000000110000000001101011000000100",
			5748 => "00000000000000000101101011011001",
			5749 => "00000000110101000101101011011001",
			5750 => "00000000000000000101101011011001",
			5751 => "0000001000000000001011010100000100",
			5752 => "00000000000000000101101011011001",
			5753 => "11111110110000110101101011011001",
			5754 => "0000001101000000001000000000001000",
			5755 => "0000000111000000001000111000000100",
			5756 => "00000000001011110101101011011001",
			5757 => "11111111100010100101101011011001",
			5758 => "00000000101110110101101011011001",
			5759 => "0000000010000000001111010100101000",
			5760 => "0000000110000000001011001100011000",
			5761 => "0000001100000000001110001100001000",
			5762 => "0000001011000000000101101100000100",
			5763 => "00000000000000000101101011011001",
			5764 => "11111111010111010101101011011001",
			5765 => "0000001011000000000101100100001100",
			5766 => "0000001110000000001011011100000100",
			5767 => "00000000000000000101101011011001",
			5768 => "0000000001000000000001111000000100",
			5769 => "00000000011110010101101011011001",
			5770 => "00000000000000000101101011011001",
			5771 => "00000000000000000101101011011001",
			5772 => "0000001010000000000111110100000100",
			5773 => "00000000000000000101101011011001",
			5774 => "0000001101000000000011100000000100",
			5775 => "00000000000000000101101011011001",
			5776 => "0000001110000000000001101000000100",
			5777 => "00000000000000000101101011011001",
			5778 => "00000001000010110101101011011001",
			5779 => "0000001011000000001011110100100100",
			5780 => "0000001000000000000010101000011100",
			5781 => "0000000010000000001000000100010000",
			5782 => "0000000000000000000011010000001000",
			5783 => "0000000001000000001001011000000100",
			5784 => "11111111001111000101101011011001",
			5785 => "00000000000111000101101011011001",
			5786 => "0000000111000000001101111000000100",
			5787 => "00000000111000000101101011011001",
			5788 => "11111111111010010101101011011001",
			5789 => "0000001111000000000011001100001000",
			5790 => "0000001100000000001001110100000100",
			5791 => "00000001001010100101101011011001",
			5792 => "00000000000000000101101011011001",
			5793 => "00000000000000000101101011011001",
			5794 => "0000000001000000001101101000000100",
			5795 => "00000000000000000101101011011001",
			5796 => "11111111001000000101101011011001",
			5797 => "0000001110000000000011110100011100",
			5798 => "0000000001000000000001111000001100",
			5799 => "0000000111000000000000011100000100",
			5800 => "11111111111000100101101011011001",
			5801 => "0000001110000000001011101100000100",
			5802 => "00000000000000000101101011011001",
			5803 => "00000000011000010101101011011001",
			5804 => "0000000110000000001000010000001000",
			5805 => "0000000000000000001010101100000100",
			5806 => "00000000000000000101101011011001",
			5807 => "00000000001011100101101011011001",
			5808 => "0000000000000000001010101100000100",
			5809 => "00000000000000000101101011011001",
			5810 => "11111111000001110101101011011001",
			5811 => "0000000110000000000000001000000100",
			5812 => "00000000110001000101101011011001",
			5813 => "00000000000000000101101011011001",
			5814 => "0000000101000000001010111000100100",
			5815 => "0000000100000000001111100000001100",
			5816 => "0000000111000000001001110000000100",
			5817 => "11111110010111110101110000001101",
			5818 => "0000000111000000001101100000000100",
			5819 => "00000000000000000101110000001101",
			5820 => "11111111100000010101110000001101",
			5821 => "0000001101000000000001111100000100",
			5822 => "11111110101010000101110000001101",
			5823 => "0000001100000000000000101000001000",
			5824 => "0000000110000000001011001100000100",
			5825 => "00000000000000000101110000001101",
			5826 => "00000001011101110101110000001101",
			5827 => "0000000110000000001001100100001000",
			5828 => "0000000100000000000111011100000100",
			5829 => "11111110110101010101110000001101",
			5830 => "00000000000000000101110000001101",
			5831 => "00000001000101100101110000001101",
			5832 => "0000000101000000000100011000100000",
			5833 => "0000001101000000001011000000010100",
			5834 => "0000000000000000000011010000000100",
			5835 => "11111110101100110101110000001101",
			5836 => "0000000010000000001100010000001000",
			5837 => "0000000110000000001101011000000100",
			5838 => "00000000000000000101110000001101",
			5839 => "00000001011110000101110000001101",
			5840 => "0000001001000000001101011100000100",
			5841 => "00000000000000000101110000001101",
			5842 => "11111111000101010101110000001101",
			5843 => "0000000110000000001101011000000100",
			5844 => "00000000000000000101110000001101",
			5845 => "0000000111000000001101100000000100",
			5846 => "00000001100110000101110000001101",
			5847 => "00000000000000000101110000001101",
			5848 => "0000001101000000001000000000011100",
			5849 => "0000000100000000000010100100010000",
			5850 => "0000000111000000001000111000000100",
			5851 => "11111111010001010101110000001101",
			5852 => "0000000001000000001001111000000100",
			5853 => "00000000000000000101110000001101",
			5854 => "0000000000000000000011111100000100",
			5855 => "00000000000000000101110000001101",
			5856 => "11111101101101100101110000001101",
			5857 => "0000000010000000000111010100001000",
			5858 => "0000001100000000001100110000000100",
			5859 => "00000001000011100101110000001101",
			5860 => "00000000000000000101110000001101",
			5861 => "00000000000000000101110000001101",
			5862 => "0000000010000000000010000100011100",
			5863 => "0000001010000000000001010000010000",
			5864 => "0000000011000000000111110000001000",
			5865 => "0000000100000000000011000000000100",
			5866 => "00000000000000000101110000001101",
			5867 => "11111110111001100101110000001101",
			5868 => "0000000001000000001101101000000100",
			5869 => "11111111111111100101110000001101",
			5870 => "00000001000100100101110000001101",
			5871 => "0000001100000000001001110000001000",
			5872 => "0000000101000000001000000000000100",
			5873 => "00000001110111000101110000001101",
			5874 => "00000000000000000101110000001101",
			5875 => "11111111101001100101110000001101",
			5876 => "0000001110000000000101100100010000",
			5877 => "0000000110000000001001100100001000",
			5878 => "0000001110000000001000000000000100",
			5879 => "00000000000000000101110000001101",
			5880 => "11111101101010110101110000001101",
			5881 => "0000001101000000000001101000000100",
			5882 => "00000001100011110101110000001101",
			5883 => "11111110110110010101110000001101",
			5884 => "0000001101000000001100111000001000",
			5885 => "0000000011000000000110111000000100",
			5886 => "00000000000000010101110000001101",
			5887 => "00000000100110010101110000001101",
			5888 => "0000001100000000000101110100000100",
			5889 => "11111110010000100101110000001101",
			5890 => "00000000000000000101110000001101",
			5891 => "0000000011000000000111110001010100",
			5892 => "0000001010000000000001010000100000",
			5893 => "0000001111000000001001010000010100",
			5894 => "0000001110000000001010001100001000",
			5895 => "0000000110000000001001011000000100",
			5896 => "00000000000000000101110101101001",
			5897 => "11111111001101100101110101101001",
			5898 => "0000000001000000000111100100000100",
			5899 => "00000000000000000101110101101001",
			5900 => "0000001000000000000000001000000100",
			5901 => "00000000000000000101110101101001",
			5902 => "00000000011001000101110101101001",
			5903 => "0000001100000000001100001000000100",
			5904 => "00000000000000000101110101101001",
			5905 => "0000001101000000000001101000000100",
			5906 => "11111110000101000101110101101001",
			5907 => "00000000000000000101110101101001",
			5908 => "0000000100000000000101000000001000",
			5909 => "0000000011000000000000011100000100",
			5910 => "00000000000000000101110101101001",
			5911 => "00000001000110110101110101101001",
			5912 => "0000000100000000000011001100010000",
			5913 => "0000000111000000000100000000000100",
			5914 => "00000000000000000101110101101001",
			5915 => "0000000001000000000110101000001000",
			5916 => "0000001100000000000000101000000100",
			5917 => "00000000000000000101110101101001",
			5918 => "11111110101111100101110101101001",
			5919 => "00000000000000000101110101101001",
			5920 => "0000000110000000001001100100010000",
			5921 => "0000000010000000001110110100001000",
			5922 => "0000000011000000001001110100000100",
			5923 => "11111111010111100101110101101001",
			5924 => "00000000111111000101110101101001",
			5925 => "0000000111000000000100000000000100",
			5926 => "00000000000000000101110101101001",
			5927 => "11111110101000110101110101101001",
			5928 => "0000001101000000000001101000001000",
			5929 => "0000000010000000000110101100000100",
			5930 => "00000000111001000101110101101001",
			5931 => "11111111110110100101110101101001",
			5932 => "11111111000010010101110101101001",
			5933 => "0000001111000000001100010000100000",
			5934 => "0000001101000000001110000100011100",
			5935 => "0000000100000000001101001000010100",
			5936 => "0000000001000000000111100100001000",
			5937 => "0000001100000000001000111000000100",
			5938 => "00000000000000000101110101101001",
			5939 => "11111111111100010101110101101001",
			5940 => "0000001001000000001001111100001000",
			5941 => "0000001000000000000010101100000100",
			5942 => "00000000000000000101110101101001",
			5943 => "00000000111111110101110101101001",
			5944 => "00000000000000000101110101101001",
			5945 => "0000000111000000000101101100000100",
			5946 => "00000000000001110101110101101001",
			5947 => "11111111111011100101110101101001",
			5948 => "00000000000000000101110101101001",
			5949 => "0000001001000000001100011000010000",
			5950 => "0000000010000000001111101000001000",
			5951 => "0000001101000000000111010000000100",
			5952 => "00000000000000000101110101101001",
			5953 => "11111110011111110101110101101001",
			5954 => "0000000000000000001011000100000100",
			5955 => "00000000110011100101110101101001",
			5956 => "00000000000000000101110101101001",
			5957 => "0000001101000000001110101100001100",
			5958 => "0000001100000000000011011100000100",
			5959 => "00000000000000000101110101101001",
			5960 => "0000000010000000001000100000000100",
			5961 => "00000000000000000101110101101001",
			5962 => "00000001010000010101110101101001",
			5963 => "0000000001000000000111101000010000",
			5964 => "0000001111000000001000110100001000",
			5965 => "0000000110000000000100111100000100",
			5966 => "00000000000000000101110101101001",
			5967 => "11111110010011100101110101101001",
			5968 => "0000000000000000000000111000000100",
			5969 => "00000000011101000101110101101001",
			5970 => "00000000000000000101110101101001",
			5971 => "0000000100000000001000001000001000",
			5972 => "0000001010000000001000100100000100",
			5973 => "00000000000000000101110101101001",
			5974 => "00000000100011000101110101101001",
			5975 => "0000001111000000000101000000000100",
			5976 => "11111111000001000101110101101001",
			5977 => "00000000000101010101110101101001",
			5978 => "0000000011000000000010001001000000",
			5979 => "0000001011000000001100101100110100",
			5980 => "0000000000000000000011010000010100",
			5981 => "0000001101000000001000000000001100",
			5982 => "0000001000000000001001101000000100",
			5983 => "00000000000000000101111010011101",
			5984 => "0000000100000000000010110000000100",
			5985 => "11111110100110000101111010011101",
			5986 => "00000000000000000101111010011101",
			5987 => "0000000100000000001000110100000100",
			5988 => "00000000000000000101111010011101",
			5989 => "00000000011000000101111010011101",
			5990 => "0000001111000000001110010000011100",
			5991 => "0000000011000000001010011100010000",
			5992 => "0000000100000000000100001100001000",
			5993 => "0000000011000000000001101000000100",
			5994 => "11111110110010110101111010011101",
			5995 => "00000000000000000101111010011101",
			5996 => "0000001011000000000101101100000100",
			5997 => "00000000011101000101111010011101",
			5998 => "11111111110000110101111010011101",
			5999 => "0000000010000000001100010000000100",
			6000 => "00000001011100110101111010011101",
			6001 => "0000000011000000000001011000000100",
			6002 => "11111111101110110101111010011101",
			6003 => "00000000111111000101111010011101",
			6004 => "11111110110010100101111010011101",
			6005 => "0000001111000000001111010000000100",
			6006 => "00000000000000000101111010011101",
			6007 => "0000000010000000000111010100000100",
			6008 => "11111101111011110101111010011101",
			6009 => "00000000000000000101111010011101",
			6010 => "0000000101000000001001001000001100",
			6011 => "0000000001000000000110101000000100",
			6012 => "11111111010000100101111010011101",
			6013 => "0000000000000000001101010000000100",
			6014 => "00000000000000000101111010011101",
			6015 => "00000001011110010101111010011101",
			6016 => "0000001011000000000111001000011100",
			6017 => "0000000110000000001000010000010100",
			6018 => "0000000111000000001101100000001000",
			6019 => "0000001011000000001110001100000100",
			6020 => "11111111111101000101111010011101",
			6021 => "00000000000000000101111010011101",
			6022 => "0000000000000000000000111000001000",
			6023 => "0000000001000000001111001100000100",
			6024 => "11111110100000110101111010011101",
			6025 => "00000000000000000101111010011101",
			6026 => "00000000000000000101111010011101",
			6027 => "0000001011000000001010111100000100",
			6028 => "00000001000000110101111010011101",
			6029 => "11111111011000000101111010011101",
			6030 => "0000001011000000001011000000010100",
			6031 => "0000000111000000001101111000001000",
			6032 => "0000000010000000000011000000000100",
			6033 => "11111111110010100101111010011101",
			6034 => "00000000000100000101111010011101",
			6035 => "0000000011000000001001010100000100",
			6036 => "00000000000000000101111010011101",
			6037 => "0000000100000000000000100000000100",
			6038 => "00000001011100000101111010011101",
			6039 => "00000000000000000101111010011101",
			6040 => "0000000000000000001111000100010000",
			6041 => "0000001111000000000110111100001000",
			6042 => "0000000101000000000110110100000100",
			6043 => "00000000000000000101111010011101",
			6044 => "11111111011110010101111010011101",
			6045 => "0000000111000000001001001000000100",
			6046 => "00000000000000000101111010011101",
			6047 => "00000000011010110101111010011101",
			6048 => "0000001000000000001001101000001000",
			6049 => "0000000011000000000110111000000100",
			6050 => "11111110010001100101111010011101",
			6051 => "00000000000000000101111010011101",
			6052 => "0000000010000000000011110100000100",
			6053 => "11111111111001110101111010011101",
			6054 => "00000000110011110101111010011101",
			6055 => "0000001011000000000011011100011000",
			6056 => "0000000010000000000111011000010000",
			6057 => "0000000101000000001101010100000100",
			6058 => "11111110011010010101111110011001",
			6059 => "0000001011000000000011011100000100",
			6060 => "11111111010000110101111110011001",
			6061 => "0000000101000000001101010100000100",
			6062 => "00000000000000110101111110011001",
			6063 => "00000000000000000101111110011001",
			6064 => "0000001000000000001111000100000100",
			6065 => "11111110111001100101111110011001",
			6066 => "00000001011011110101111110011001",
			6067 => "0000001010000000001011010101100000",
			6068 => "0000000110000000001000010000111000",
			6069 => "0000001100000000000100000000011000",
			6070 => "0000000110000000001011001100001100",
			6071 => "0000001111000000001100100100001000",
			6072 => "0000001010000000001010110000000100",
			6073 => "11111110111010110101111110011001",
			6074 => "00000001110010000101111110011001",
			6075 => "11111110010001010101111110011001",
			6076 => "0000000010000000001100000000000100",
			6077 => "00000001110110000101111110011001",
			6078 => "0000001101000000001000000000000100",
			6079 => "11111110110110100101111110011001",
			6080 => "00000001101001000101111110011001",
			6081 => "0000000011000000001000011000010000",
			6082 => "0000001011000000001100110000001000",
			6083 => "0000000110000000001011001100000100",
			6084 => "11111110111100110101111110011001",
			6085 => "00000001001000000101111110011001",
			6086 => "0000001000000000001000110000000100",
			6087 => "11111110000110100101111110011001",
			6088 => "00000000001110100101111110011001",
			6089 => "0000001110000000000110100100001000",
			6090 => "0000001011000000001100101100000100",
			6091 => "00000001111110100101111110011001",
			6092 => "11111110111010010101111110011001",
			6093 => "0000000011000000000000011100000100",
			6094 => "11111110011110010101111110011001",
			6095 => "11111111111010100101111110011001",
			6096 => "0000001101000000000111111100010000",
			6097 => "0000001000000000000110001000000100",
			6098 => "00000001101000000101111110011001",
			6099 => "0000001011000000001010111100000100",
			6100 => "00000001101110000101111110011001",
			6101 => "0000000001000000001111001100000100",
			6102 => "11111110010001000101111110011001",
			6103 => "00000000101101000101111110011001",
			6104 => "0000001111000000001000000100001100",
			6105 => "0000001011000000000010001000000100",
			6106 => "00000000011110010101111110011001",
			6107 => "0000001110000000001100111000000100",
			6108 => "00000000000000000101111110011001",
			6109 => "11111110011010010101111110011001",
			6110 => "0000001100000000000100011000000100",
			6111 => "11111110101011110101111110011001",
			6112 => "0000001011000000001011110100000100",
			6113 => "00000001011100100101111110011001",
			6114 => "00000000001001000101111110011001",
			6115 => "0000001100000000001000111100000100",
			6116 => "00000000000000000101111110011001",
			6117 => "11111110010111100101111110011001",
			6118 => "0000001101000000001110110000010100",
			6119 => "0000000100000000000000101100000100",
			6120 => "11111110011110000110000010110101",
			6121 => "0000000000000000000011011100001000",
			6122 => "0000001010000000000001010100000100",
			6123 => "00000000000000000110000010110101",
			6124 => "00000000010101000110000010110101",
			6125 => "0000000010000000000111010100000100",
			6126 => "11111111001101010110000010110101",
			6127 => "00000000000000000110000010110101",
			6128 => "0000000100000000001000001000110000",
			6129 => "0000000001000000000110101000001100",
			6130 => "0000000100000000000110001100000100",
			6131 => "11111110001011010110000010110101",
			6132 => "0000000101000000001110110000000100",
			6133 => "00000000000000000110000010110101",
			6134 => "00000000001010010110000010110101",
			6135 => "0000001100000000000100000000001000",
			6136 => "0000000011000000000010001000000100",
			6137 => "00000000000000000110000010110101",
			6138 => "00000001100100100110000010110101",
			6139 => "0000001100000000000100011000001100",
			6140 => "0000000111000000001000111000000100",
			6141 => "00000001101001010110000010110101",
			6142 => "0000000101000000000001000000000100",
			6143 => "00000000000101000110000010110101",
			6144 => "11111110110000010110000010110101",
			6145 => "0000001001000000000101010000001000",
			6146 => "0000000111000000000101100100000100",
			6147 => "11111110111000110110000010110101",
			6148 => "00000000011001100110000010110101",
			6149 => "0000001001000000001010100100000100",
			6150 => "00000001000010100110000010110101",
			6151 => "00000000010001110110000010110101",
			6152 => "0000000111000000001100101000011000",
			6153 => "0000001010000000001010110000000100",
			6154 => "11111110011001110110000010110101",
			6155 => "0000000011000000001001011100010000",
			6156 => "0000000010000000001111010100001000",
			6157 => "0000000011000000001011011100000100",
			6158 => "00000000010010110110000010110101",
			6159 => "00000001110110000110000010110101",
			6160 => "0000001010000000000101000100000100",
			6161 => "11111111001101010110000010110101",
			6162 => "00000000010100100110000010110101",
			6163 => "00000001101101110110000010110101",
			6164 => "0000000010000000001000000100010100",
			6165 => "0000001010000000001100011100001100",
			6166 => "0000000100000000000000010100000100",
			6167 => "11111101110111010110000010110101",
			6168 => "0000001010000000001001000100000100",
			6169 => "00000000001001000110000010110101",
			6170 => "00000000000000000110000010110101",
			6171 => "0000000100000000001001000000000100",
			6172 => "00000000010001000110000010110101",
			6173 => "11111111101111110110000010110101",
			6174 => "0000001000000000000001110100010000",
			6175 => "0000001100000000000001101000001000",
			6176 => "0000001010000000000001010000000100",
			6177 => "00000000000000000110000010110101",
			6178 => "00000001001110000110000010110101",
			6179 => "0000000101000000001110110100000100",
			6180 => "11111110111110010110000010110101",
			6181 => "00000000100110110110000010110101",
			6182 => "0000001110000000000010100100001000",
			6183 => "0000000010000000001101001000000100",
			6184 => "11111111110001110110000010110101",
			6185 => "11111110000110000110000010110101",
			6186 => "0000001101000000001100111000000100",
			6187 => "00000000111111110110000010110101",
			6188 => "11111111100001110110000010110101",
			6189 => "0000001011000000000011011100011000",
			6190 => "0000000010000000000111011000010000",
			6191 => "0000000101000000001101010100000100",
			6192 => "11111110011001110110000110111001",
			6193 => "0000001011000000000011011100000100",
			6194 => "11111111001110100110000110111001",
			6195 => "0000000101000000001101010100000100",
			6196 => "00000000000000110110000110111001",
			6197 => "00000000000000000110000110111001",
			6198 => "0000001000000000001111000100000100",
			6199 => "11111110110111000110000110111001",
			6200 => "00000001100011100110000110111001",
			6201 => "0000001010000000001011010101100100",
			6202 => "0000000110000000001000010000110100",
			6203 => "0000001100000000000100000000011000",
			6204 => "0000000100000000000010111000001100",
			6205 => "0000000001000000000110101000001000",
			6206 => "0000001111000000000101110000000100",
			6207 => "11111111110000010110000110111001",
			6208 => "11111100110010100110000110111001",
			6209 => "00000001100000110110000110111001",
			6210 => "0000000101000000000111001000001000",
			6211 => "0000001111000000000110100000000100",
			6212 => "00000001100110110110000110111001",
			6213 => "11111110100010100110000110111001",
			6214 => "00000001110110100110000110111001",
			6215 => "0000001101000000001011000000001100",
			6216 => "0000001100000000000100000000000100",
			6217 => "11111100001100000110000110111001",
			6218 => "0000000100000000000010100100000100",
			6219 => "11111110111011110110000110111001",
			6220 => "00000000100001110110000110111001",
			6221 => "0000001011000000000110000100001000",
			6222 => "0000000110000000001011001100000100",
			6223 => "00000000000000000110000110111001",
			6224 => "00000001100100100110000110111001",
			6225 => "0000000100000000001100001100000100",
			6226 => "11111111111101010110000110111001",
			6227 => "11111111000011100110000110111001",
			6228 => "0000001101000000000111111100010100",
			6229 => "0000001000000000000110001000000100",
			6230 => "00000001101001000110000110111001",
			6231 => "0000001100000000000110000100001000",
			6232 => "0000001000000000001111001000000100",
			6233 => "11111111001101100110000110111001",
			6234 => "00000001100100000110000110111001",
			6235 => "0000000001000000000101011100000100",
			6236 => "11111101101111100110000110111001",
			6237 => "00000000101110010110000110111001",
			6238 => "0000001111000000001000000100001100",
			6239 => "0000001011000000000010001000000100",
			6240 => "00000000100001000110000110111001",
			6241 => "0000001110000000001100111000000100",
			6242 => "00000000000000000110000110111001",
			6243 => "11111110010111000110000110111001",
			6244 => "0000000000000000000111000000001000",
			6245 => "0000001111000000001000110100000100",
			6246 => "11111111110001000110000110111001",
			6247 => "00000001111010110110000110111001",
			6248 => "0000001010000000001001000100000100",
			6249 => "11111110110000000110000110111001",
			6250 => "00000000011000100110000110111001",
			6251 => "0000000101000000000100011000000100",
			6252 => "00000000000000000110000110111001",
			6253 => "11111110010101110110000110111001",
			6254 => "0000000100000000001000000101001000",
			6255 => "0000000100000000001111100100011000",
			6256 => "0000000011000000001010000100010100",
			6257 => "0000001010000000000010101100010000",
			6258 => "0000001011000000000101100100001100",
			6259 => "0000000001000000001011111100000100",
			6260 => "00000000000000000110001100001101",
			6261 => "0000001011000000000000011100000100",
			6262 => "00000000000000000110001100001101",
			6263 => "00000000110110010110001100001101",
			6264 => "00000000000000000110001100001101",
			6265 => "00000000000000000110001100001101",
			6266 => "11111111101000000110001100001101",
			6267 => "0000000011000000001100111000100000",
			6268 => "0000000111000000001100101000010000",
			6269 => "0000001100000000001001110000001100",
			6270 => "0000000011000000001011011100000100",
			6271 => "00000000000000000110001100001101",
			6272 => "0000000111000000000101101100000100",
			6273 => "00000000110100000110001100001101",
			6274 => "00000000000000000110001100001101",
			6275 => "11111111100000010110001100001101",
			6276 => "0000001100000000001000000000001100",
			6277 => "0000001001000000001010100100001000",
			6278 => "0000001001000000000111101100000100",
			6279 => "00000001001000100110001100001101",
			6280 => "00000000010111100110001100001101",
			6281 => "00000000000000000110001100001101",
			6282 => "00000000000000000110001100001101",
			6283 => "0000001100000000001001001000001000",
			6284 => "0000000010000000000011000000000100",
			6285 => "11111111010000110110001100001101",
			6286 => "00000000000000000110001100001101",
			6287 => "0000001100000000000001101000000100",
			6288 => "00000000100110000110001100001101",
			6289 => "00000000000000000110001100001101",
			6290 => "0000000100000000001000110100001100",
			6291 => "0000000001000000000001111000001000",
			6292 => "0000000000000000000010011000000100",
			6293 => "11111110110011110110001100001101",
			6294 => "00000000000000000110001100001101",
			6295 => "00000000000000000110001100001101",
			6296 => "0000001111000000001110000000111100",
			6297 => "0000000111000000000101101100011100",
			6298 => "0000000011000000000000011100010000",
			6299 => "0000001011000000000101101100001000",
			6300 => "0000000100000000001001001100000100",
			6301 => "11111111010111110110001100001101",
			6302 => "00000000011111110110001100001101",
			6303 => "0000000010000000000010000000000100",
			6304 => "00000000000000000110001100001101",
			6305 => "11111111000101010110001100001101",
			6306 => "0000001010000000000001010000000100",
			6307 => "11111111011111110110001100001101",
			6308 => "0000000010000000001100000000000100",
			6309 => "00000001000100000110001100001101",
			6310 => "00000000000000000110001100001101",
			6311 => "0000001010000000000101000100010000",
			6312 => "0000001001000000000111101100001000",
			6313 => "0000001010000000001000100100000100",
			6314 => "00000000000000000110001100001101",
			6315 => "11111110111001100110001100001101",
			6316 => "0000001011000000000101110100000100",
			6317 => "00000000001000100110001100001101",
			6318 => "00000000000000000110001100001101",
			6319 => "0000001010000000000001110000001000",
			6320 => "0000001110000000001011011100000100",
			6321 => "00000000000000000110001100001101",
			6322 => "00000000100110110110001100001101",
			6323 => "0000000111000000000101101100000100",
			6324 => "00000000000000000110001100001101",
			6325 => "11111111110001100110001100001101",
			6326 => "0000001010000000000110011100010000",
			6327 => "0000000000000000001010101100000100",
			6328 => "00000000000000000110001100001101",
			6329 => "0000000111000000000111010000000100",
			6330 => "00000000111100000110001100001101",
			6331 => "0000000111000000000000011100000100",
			6332 => "00000000000000000110001100001101",
			6333 => "00000000010100010110001100001101",
			6334 => "0000001110000000000010100100001000",
			6335 => "0000000010000000001101001000000100",
			6336 => "00000000000000000110001100001101",
			6337 => "11111110111001000110001100001101",
			6338 => "00000000000000000110001100001101",
			6339 => "0000000110000000001001100101001000",
			6340 => "0000000101000000000111001000000100",
			6341 => "11111110100111110110010000111001",
			6342 => "0000001111000000001110000100011100",
			6343 => "0000000110000000001101011000001100",
			6344 => "0000000010000000000110100000001000",
			6345 => "0000000000000000000110011000000100",
			6346 => "00000000000000000110010000111001",
			6347 => "00000000100000110110010000111001",
			6348 => "11111110111000100110010000111001",
			6349 => "0000000100000000000010111000000100",
			6350 => "00000000000000000110010000111001",
			6351 => "0000000011000000001001110100000100",
			6352 => "00000000000000000110010000111001",
			6353 => "0000001100000000001001110000000100",
			6354 => "00000001010110000110010000111001",
			6355 => "00000000000000000110010000111001",
			6356 => "0000000100000000001000000100010100",
			6357 => "0000001001000000001110010100001000",
			6358 => "0000000100000000001011110000000100",
			6359 => "00000000000000000110010000111001",
			6360 => "00000001000010110110010000111001",
			6361 => "0000001001000000001000010000000100",
			6362 => "11111110110010010110010000111001",
			6363 => "0000001100000000001011000000000100",
			6364 => "00000000000000110110010000111001",
			6365 => "11111111000001000110010000111001",
			6366 => "0000000010000000001100010000001100",
			6367 => "0000000010000000000110010000000100",
			6368 => "11111111011111000110010000111001",
			6369 => "0000001100000000001000111000000100",
			6370 => "00000000001011010110010000111001",
			6371 => "00000000000000000110010000111001",
			6372 => "0000001100000000000111001000000100",
			6373 => "11111110011011000110010000111001",
			6374 => "00000000000000000110010000111001",
			6375 => "0000000111000000001101100000011100",
			6376 => "0000001011000000001100101100011000",
			6377 => "0000001111000000001110010000010100",
			6378 => "0000001100000000001000111100010000",
			6379 => "0000001101000000001110110000001000",
			6380 => "0000000010000000000010000100000100",
			6381 => "11111111110101010110010000111001",
			6382 => "00000000001000000110010000111001",
			6383 => "0000001001000000001111001100000100",
			6384 => "00000000000000000110010000111001",
			6385 => "00000001011111010110010000111001",
			6386 => "11111111101000110110010000111001",
			6387 => "11111111001001010110010000111001",
			6388 => "00000001100001000110010000111001",
			6389 => "0000001100000000000100000000001000",
			6390 => "0000001000000000001011010100000100",
			6391 => "00000000000000000110010000111001",
			6392 => "11111110011010100110010000111001",
			6393 => "0000000000000000000111111000011100",
			6394 => "0000001010000000001100011100010000",
			6395 => "0000001000000000000111000100001000",
			6396 => "0000001000000000000110001000000100",
			6397 => "11111111111011010110010000111001",
			6398 => "00000000110000110110010000111001",
			6399 => "0000001111000000000110010000000100",
			6400 => "00000000000000000110010000111001",
			6401 => "11111101101011100110010000111001",
			6402 => "0000001100000000001000000000000100",
			6403 => "00000001100001100110010000111001",
			6404 => "0000001111000000000000010100000100",
			6405 => "11111110101010100110010000111001",
			6406 => "00000000110011000110010000111001",
			6407 => "0000000111000000001101100000000100",
			6408 => "00000000000110110110010000111001",
			6409 => "0000000011000000000011011000000100",
			6410 => "11111110100101010110010000111001",
			6411 => "0000001010000000000010101000000100",
			6412 => "00000000001010110110010000111001",
			6413 => "00000000000000000110010000111001",
			6414 => "0000000011000000001011000000010100",
			6415 => "0000000110000000001001100100000100",
			6416 => "11111110011001110110010101111101",
			6417 => "0000001011000000000011011100000100",
			6418 => "11111111011101000110010101111101",
			6419 => "0000000010000000000111011000000100",
			6420 => "00000001110000110110010101111101",
			6421 => "0000001010000000001111001000000100",
			6422 => "11111111100111110110010101111101",
			6423 => "00000000000000000110010101111101",
			6424 => "0000000110000000000100111101000100",
			6425 => "0000001011000000000110110100110000",
			6426 => "0000000110000000001100011000010000",
			6427 => "0000001001000000000101011100001100",
			6428 => "0000000001000000000110101000000100",
			6429 => "11111110110111000110010101111101",
			6430 => "0000000000000000001010100000000100",
			6431 => "00000000000000000110010101111101",
			6432 => "00000001001001010110010101111101",
			6433 => "11111110100010010110010101111101",
			6434 => "0000000100000000000011000000010000",
			6435 => "0000001001000000000111101100001000",
			6436 => "0000001001000000001011111100000100",
			6437 => "11111110101100110110010101111101",
			6438 => "00000001001110110110010101111101",
			6439 => "0000001010000000000111110100000100",
			6440 => "11111110111100110110010101111101",
			6441 => "00000001111010000110010101111101",
			6442 => "0000001111000000001001010000001000",
			6443 => "0000000100000000001111100000000100",
			6444 => "00000000001110010110010101111101",
			6445 => "00000001110011100110010101111101",
			6446 => "0000001101000000001000000000000100",
			6447 => "11111110000010110110010101111101",
			6448 => "00000000000010100110010101111101",
			6449 => "0000000001000000001110010100001100",
			6450 => "0000001111000000001011101100000100",
			6451 => "11111110100110110110010101111101",
			6452 => "0000000001000000000101011100000100",
			6453 => "00000000000000000110010101111101",
			6454 => "00000001101011010110010101111101",
			6455 => "0000001000000000000001010100000100",
			6456 => "11111110011001010110010101111101",
			6457 => "11111100001111000110010101111101",
			6458 => "0000000101000000000001000000011100",
			6459 => "0000000100000000000111011100010000",
			6460 => "0000001110000000000011001000001000",
			6461 => "0000001011000000000001111100000100",
			6462 => "00000001101010110110010101111101",
			6463 => "11111111001110110110010101111101",
			6464 => "0000001000000000000001010100000100",
			6465 => "00000000001111110110010101111101",
			6466 => "00000001101001110110010101111101",
			6467 => "0000001001000000000001000100000100",
			6468 => "00000001101011100110010101111101",
			6469 => "0000000110000000000101010000000100",
			6470 => "11111110001111010110010101111101",
			6471 => "00000000001010110110010101111101",
			6472 => "0000001111000000001000000100010100",
			6473 => "0000001001000000000011101000001100",
			6474 => "0000001101000000000111111100000100",
			6475 => "00000000000000000110010101111101",
			6476 => "0000001111000000001110000000000100",
			6477 => "11111110001011110110010101111101",
			6478 => "11111111111011000110010101111101",
			6479 => "0000001111000000000110111000000100",
			6480 => "00000010000110010110010101111101",
			6481 => "11111110111000110110010101111101",
			6482 => "0000000100000000000000010100010000",
			6483 => "0000000001000000001101011000001000",
			6484 => "0000001111000000001000110100000100",
			6485 => "11111111100110000110010101111101",
			6486 => "00000001110110100110010101111101",
			6487 => "0000001101000000001110110100000100",
			6488 => "00000000010011110110010101111101",
			6489 => "11111110100011010110010101111101",
			6490 => "0000000000000000001011000100001000",
			6491 => "0000000100000000000011101100000100",
			6492 => "11111111000110000110010101111101",
			6493 => "00000000101011010110010101111101",
			6494 => "11111110011010110110010101111101",
			6495 => "0000001011000000000011011100001000",
			6496 => "0000000010000000000111011000000100",
			6497 => "11111110101111100110011001110001",
			6498 => "00000000000000000110011001110001",
			6499 => "0000001100000000001100001000010100",
			6500 => "0000000100000000000010110000001000",
			6501 => "0000000011000000000101110100000100",
			6502 => "11111110110001000110011001110001",
			6503 => "00000000100011000110011001110001",
			6504 => "0000000101000000001010111100000100",
			6505 => "00000000000000000110011001110001",
			6506 => "0000000110000000001011001100000100",
			6507 => "00000000000000000110011001110001",
			6508 => "00000001011101010110011001110001",
			6509 => "0000000100000000001000000100100100",
			6510 => "0000000101000000001000000000001000",
			6511 => "0000000110000000001011001100000100",
			6512 => "00000000000000000110011001110001",
			6513 => "00000001011001000110011001110001",
			6514 => "0000000011000000000001001000001100",
			6515 => "0000001111000000000010110100001000",
			6516 => "0000001100000000000110000100000100",
			6517 => "00000000000000000110011001110001",
			6518 => "00000000001101010110011001110001",
			6519 => "11111110100010000110011001110001",
			6520 => "0000000000000000000111000100001000",
			6521 => "0000000010000000001000100000000100",
			6522 => "00000000000110010110011001110001",
			6523 => "11111110111111100110011001110001",
			6524 => "0000000101000000001100100100000100",
			6525 => "00000000111101110110011001110001",
			6526 => "00000000000000000110011001110001",
			6527 => "0000000110000000000100111100011100",
			6528 => "0000001011000000000110000100001100",
			6529 => "0000001101000000001110110000000100",
			6530 => "11111111001111000110011001110001",
			6531 => "0000000010000000000111011000000100",
			6532 => "00000001000001010110011001110001",
			6533 => "11111111101110110110011001110001",
			6534 => "0000000100000000000110001100001000",
			6535 => "0000000000000000000010111100000100",
			6536 => "11111110001111110110011001110001",
			6537 => "11111111111011000110011001110001",
			6538 => "0000000011000000001001010100000100",
			6539 => "11111111001000100110011001110001",
			6540 => "00000000111110000110011001110001",
			6541 => "0000001100000000000110000100010000",
			6542 => "0000000000000000000011010000001000",
			6543 => "0000000101000000000001101000000100",
			6544 => "00000000011111100110011001110001",
			6545 => "11111111101100010110011001110001",
			6546 => "0000001011000000000110000100000100",
			6547 => "00000000000000000110011001110001",
			6548 => "00000001010100010110011001110001",
			6549 => "0000001110000000001011101100001000",
			6550 => "0000000100000000001000001000000100",
			6551 => "00000000011110110110011001110001",
			6552 => "11111110010111100110011001110001",
			6553 => "0000001101000000001010001000000100",
			6554 => "00000000111110010110011001110001",
			6555 => "11111111110101010110011001110001",
			6556 => "0000000101000000000111100010001000",
			6557 => "0000000111000000001110110001001100",
			6558 => "0000001000000000000110001000011000",
			6559 => "0000001100000000000100000000001000",
			6560 => "0000000110000000001011001100000100",
			6561 => "00000000000000000110100000011101",
			6562 => "00000000000011110110100000011101",
			6563 => "0000001111000000001001010000000100",
			6564 => "00000000000000000110100000011101",
			6565 => "0000000010000000001100010100000100",
			6566 => "00000000000000000110100000011101",
			6567 => "0000000110000000001000010000000100",
			6568 => "11111110111100010110100000011101",
			6569 => "00000000000000000110100000011101",
			6570 => "0000000011000000001011011100011100",
			6571 => "0000001111000000001111010000010000",
			6572 => "0000000011000000001001110100001000",
			6573 => "0000001111000000000110100000000100",
			6574 => "00000000000000000110100000011101",
			6575 => "11111111010000000110100000011101",
			6576 => "0000000001000000000110101000000100",
			6577 => "00000000101011110110100000011101",
			6578 => "11111111111101100110100000011101",
			6579 => "0000000111000000001000111000000100",
			6580 => "00000000000000000110100000011101",
			6581 => "0000000110000000001111000000000100",
			6582 => "11111110110001110110100000011101",
			6583 => "00000000000000000110100000011101",
			6584 => "0000000010000000000110111100001000",
			6585 => "0000000000000000000000111000000100",
			6586 => "00000001000100000110100000011101",
			6587 => "00000000000000000110100000011101",
			6588 => "0000001010000000001100011100001000",
			6589 => "0000001100000000001000111100000100",
			6590 => "00000000000000000110100000011101",
			6591 => "11111111010100110110100000011101",
			6592 => "0000001000000000001101010000000100",
			6593 => "00000000101100100110100000011101",
			6594 => "11111111101011110110100000011101",
			6595 => "0000001111000000001111010100011000",
			6596 => "0000001100000000001010111000010000",
			6597 => "0000001010000000000011101000001100",
			6598 => "0000000111000000001001001000001000",
			6599 => "0000000001000000000111101000000100",
			6600 => "00000000011100000110100000011101",
			6601 => "00000000000000000110100000011101",
			6602 => "00000000000000000110100000011101",
			6603 => "00000000000000000110100000011101",
			6604 => "0000000111000000001000011000000100",
			6605 => "11111111010001100110100000011101",
			6606 => "00000000000000000110100000011101",
			6607 => "0000000111000000000001101000011000",
			6608 => "0000000111000000001001001000001100",
			6609 => "0000001100000000000100011000001000",
			6610 => "0000001100000000000100001000000100",
			6611 => "00000000000000000110100000011101",
			6612 => "00000000101111010110100000011101",
			6613 => "00000000000000000110100000011101",
			6614 => "0000001111000000001010000100000100",
			6615 => "00000000000000000110100000011101",
			6616 => "0000000111000000000110100100000100",
			6617 => "11111111011010100110100000011101",
			6618 => "00000000000000000110100000011101",
			6619 => "0000001100000000000111001000000100",
			6620 => "00000000000000000110100000011101",
			6621 => "0000001101000000001110000100000100",
			6622 => "00000000000000000110100000011101",
			6623 => "00000000111010100110100000011101",
			6624 => "0000000011000000000110111000011000",
			6625 => "0000000001000000000100110100001100",
			6626 => "0000000111000000000101100100001000",
			6627 => "0000001001000000001010100100000100",
			6628 => "11111110110000100110100000011101",
			6629 => "00000000000000000110100000011101",
			6630 => "00000000000000000110100000011101",
			6631 => "0000000111000000001000011000000100",
			6632 => "00000000010011100110100000011101",
			6633 => "0000000111000000001111011100000100",
			6634 => "11111111101101100110100000011101",
			6635 => "00000000000000000110100000011101",
			6636 => "0000001101000000001100010100001100",
			6637 => "0000001100000000000100011000000100",
			6638 => "00000000000000000110100000011101",
			6639 => "0000001111000000001000011100000100",
			6640 => "00000000000000000110100000011101",
			6641 => "00000000101110000110100000011101",
			6642 => "0000001110000000000010110000011000",
			6643 => "0000000110000000001000010000001100",
			6644 => "0000001100000000001111011100000100",
			6645 => "00000000000000000110100000011101",
			6646 => "0000000111000000001011011100000100",
			6647 => "00000000000000000110100000011101",
			6648 => "00000000011011000110100000011101",
			6649 => "0000001010000000001000010100000100",
			6650 => "00000000000000000110100000011101",
			6651 => "0000000101000000001100010000000100",
			6652 => "11111110111011000110100000011101",
			6653 => "00000000000000000110100000011101",
			6654 => "0000001101000000001101101100001100",
			6655 => "0000000001000000001101111100000100",
			6656 => "00000000000000000110100000011101",
			6657 => "0000000010000000001101001000000100",
			6658 => "00000000000000000110100000011101",
			6659 => "00000000101110110110100000011101",
			6660 => "0000001100000000000101110100000100",
			6661 => "11111111101001010110100000011101",
			6662 => "00000000000000000110100000011101",
			6663 => "0000000101000000001010111100010100",
			6664 => "0000000010000000001100000000000100",
			6665 => "11111110011110000110100100001001",
			6666 => "0000000100000000000000101100000100",
			6667 => "11111111001110100110100100001001",
			6668 => "0000000010000000000000010000001000",
			6669 => "0000000000000000000100000000000100",
			6670 => "00000000000000000110100100001001",
			6671 => "00000000101111110110100100001001",
			6672 => "11111111100000110110100100001001",
			6673 => "0000001101000000001101101101100000",
			6674 => "0000000100000000000011001100111100",
			6675 => "0000000001000000000101011100011100",
			6676 => "0000000010000000001100000000010000",
			6677 => "0000000000000000000010011000001000",
			6678 => "0000000001000000000111100100000100",
			6679 => "11111110100000110110100100001001",
			6680 => "00000000001110100110100100001001",
			6681 => "0000001100000000001001110000000100",
			6682 => "00000000101110010110100100001001",
			6683 => "11111101111100010110100100001001",
			6684 => "0000001000000000000111000100001000",
			6685 => "0000001010000000001010110000000100",
			6686 => "11111110100100100110100100001001",
			6687 => "00000000100000110110100100001001",
			6688 => "11111101011100100110100100001001",
			6689 => "0000000101000000000111100000010000",
			6690 => "0000001100000000000100011000001000",
			6691 => "0000000010000000000000010000000100",
			6692 => "11111111111111110110100100001001",
			6693 => "00000000111101000110100100001001",
			6694 => "0000001011000000001011011100000100",
			6695 => "00000001011101110110100100001001",
			6696 => "00000000000011110110100100001001",
			6697 => "0000000001000000000100110100001000",
			6698 => "0000000001000000000101011100000100",
			6699 => "00000001001010010110100100001001",
			6700 => "11111111000100010110100100001001",
			6701 => "0000000111000000000110110100000100",
			6702 => "00000000110011110110100100001001",
			6703 => "11111111100100100110100100001001",
			6704 => "0000001100000000000000101000001000",
			6705 => "0000000110000000001011001100000100",
			6706 => "00000000000000000110100100001001",
			6707 => "00000001110010110110100100001001",
			6708 => "0000001110000000000011100000001100",
			6709 => "0000000111000000001101100000001000",
			6710 => "0000000100000000000010100100000100",
			6711 => "11111111000001000110100100001001",
			6712 => "00000001000111110110100100001001",
			6713 => "11111110001101010110100100001001",
			6714 => "0000001100000000001100110000001000",
			6715 => "0000000101000000001010111000000100",
			6716 => "11111111010110000110100100001001",
			6717 => "00000001000111010110100100001001",
			6718 => "0000000010000000001000000100000100",
			6719 => "11111110110011000110100100001001",
			6720 => "00000000011100110110100100001001",
			6721 => "11111110010101000110100100001001",
			6722 => "0000001001000000001011111101010000",
			6723 => "0000000111000000001000111000100000",
			6724 => "0000000110000000001101011000000100",
			6725 => "11111110110001000110101001111101",
			6726 => "0000000011000000001001110100010000",
			6727 => "0000000111000000001000111000001100",
			6728 => "0000001011000000001000111100000100",
			6729 => "00000000000000000110101001111101",
			6730 => "0000000110000000001001100100000100",
			6731 => "00000000000000000110101001111101",
			6732 => "00000001000000010110101001111101",
			6733 => "11111111010111000110101001111101",
			6734 => "0000000010000000001111010100001000",
			6735 => "0000000111000000001000111100000100",
			6736 => "00000000000000000110101001111101",
			6737 => "00000001011111000110101001111101",
			6738 => "00000000000000000110101001111101",
			6739 => "0000000100000000000010010000100000",
			6740 => "0000001111000000000010000000011000",
			6741 => "0000000110000000000100111100010000",
			6742 => "0000000010000000001100000000001000",
			6743 => "0000001100000000001001110000000100",
			6744 => "00000000000000100110101001111101",
			6745 => "11111110100001010110101001111101",
			6746 => "0000001101000000001001001000000100",
			6747 => "11111110100011010110101001111101",
			6748 => "11111111110101010110101001111101",
			6749 => "0000000110000000000100111100000100",
			6750 => "00000001001010010110101001111101",
			6751 => "00000000000000000110101001111101",
			6752 => "0000000110000000001000010000000100",
			6753 => "11111110000010010110101001111101",
			6754 => "00000000000000000110101001111101",
			6755 => "0000001100000000000011011100001100",
			6756 => "0000000110000000001001100100000100",
			6757 => "00000000000000000110101001111101",
			6758 => "0000000100000000000000000100000100",
			6759 => "00000001001000110110101001111101",
			6760 => "00000000000000000110101001111101",
			6761 => "00000000000000000110101001111101",
			6762 => "0000001111000000001111100100110000",
			6763 => "0000001011000000001011011100101100",
			6764 => "0000001011000000000000011100011000",
			6765 => "0000001000000000000101000100001100",
			6766 => "0000000011000000000101110100000100",
			6767 => "00000000000000000110101001111101",
			6768 => "0000001111000000000000010000000100",
			6769 => "11111110101100100110101001111101",
			6770 => "00000000000000000110101001111101",
			6771 => "0000001111000000000000010000001000",
			6772 => "0000000101000000000001101000000100",
			6773 => "00000000111000100110101001111101",
			6774 => "11111111110100000110101001111101",
			6775 => "00000001011110110110101001111101",
			6776 => "0000000111000000001001001000000100",
			6777 => "11111111110111100110101001111101",
			6778 => "0000000111000000000110100100001000",
			6779 => "0000000010000000001000001100000100",
			6780 => "00000010001110010110101001111101",
			6781 => "00000000000000000110101001111101",
			6782 => "0000000111000000000110100100000100",
			6783 => "00000000000000000110101001111101",
			6784 => "00000000111000110110101001111101",
			6785 => "11111111001011000110101001111101",
			6786 => "0000001001000000000100111100001100",
			6787 => "0000000111000000001100101000000100",
			6788 => "00000000000000000110101001111101",
			6789 => "0000000000000000000010111100000100",
			6790 => "00000000000000000110101001111101",
			6791 => "11111110011001000110101001111101",
			6792 => "0000000101000000001110101000010000",
			6793 => "0000000000000000000001110100000100",
			6794 => "00000000000000000110101001111101",
			6795 => "0000001111000000001110000000001000",
			6796 => "0000001001000000001010100000000100",
			6797 => "00000001011000110110101001111101",
			6798 => "00000000000000000110101001111101",
			6799 => "00000000000000000110101001111101",
			6800 => "0000000101000000000010011100010000",
			6801 => "0000000011000000000110111000001000",
			6802 => "0000000100000000001101001000000100",
			6803 => "11111111100011010110101001111101",
			6804 => "11111110001011000110101001111101",
			6805 => "0000001111000000000011001100000100",
			6806 => "00000001000001010110101001111101",
			6807 => "00000000000000000110101001111101",
			6808 => "0000001011000000001011110100001000",
			6809 => "0000001011000000000101110100000100",
			6810 => "00000000000000000110101001111101",
			6811 => "00000001010110000110101001111101",
			6812 => "0000001100000000001001110100000100",
			6813 => "11111110111001100110101001111101",
			6814 => "00000000001111000110101001111101",
			6815 => "0000000110000000001011001101011000",
			6816 => "0000000001000000000101011100110000",
			6817 => "0000000110000000001011001100011100",
			6818 => "0000000110000000001001011000001000",
			6819 => "0000001100000000001100110000000100",
			6820 => "11111110011110100110110000011001",
			6821 => "00000100010011100110110000011001",
			6822 => "0000000011000000001010001100000100",
			6823 => "11111110010111000110110000011001",
			6824 => "0000001110000000000110100100001000",
			6825 => "0000000110000000001101011000000100",
			6826 => "11111110111100000110110000011001",
			6827 => "00000100001101000110110000011001",
			6828 => "0000001101000000000100010000000100",
			6829 => "11111111010000010110110000011001",
			6830 => "11111110010111100110110000011001",
			6831 => "0000000010000000000010000100010000",
			6832 => "0000001110000000001010111000000100",
			6833 => "11111110011100110110110000011001",
			6834 => "0000001010000000001010110000001000",
			6835 => "0000000000000000000010011000000100",
			6836 => "00000000110001100110110000011001",
			6837 => "11111110011101100110110000011001",
			6838 => "00000011010110010110110000011001",
			6839 => "11111110011001110110110000011001",
			6840 => "0000000011000000001100000000001000",
			6841 => "0000000001000000000101011100000100",
			6842 => "00000000111011100110110000011001",
			6843 => "11111110011001100110110000011001",
			6844 => "0000000000000000001001101000010000",
			6845 => "0000000111000000000110100100000100",
			6846 => "00000010110010010110110000011001",
			6847 => "0000000001000000000111101000001000",
			6848 => "0000001011000000000101100100000100",
			6849 => "00000000110000010110110000011001",
			6850 => "11111110011100000110110000011001",
			6851 => "00000001101010110110110000011001",
			6852 => "0000001010000000000011101000001100",
			6853 => "0000000001000000001110010100000100",
			6854 => "00001000001100010110110000011001",
			6855 => "0000001101000000001001010000000100",
			6856 => "00000011111101010110110000011001",
			6857 => "11111111111011110110110000011001",
			6858 => "11111110010001010110110000011001",
			6859 => "0000001011000000000001001001001100",
			6860 => "0000001000000000000001010100100100",
			6861 => "0000000100000000001000000100011100",
			6862 => "0000000000000000000001110100010000",
			6863 => "0000000101000000001101000100001000",
			6864 => "0000001110000000001111010100000100",
			6865 => "00000000001101110110110000011001",
			6866 => "00000100110000000110110000011001",
			6867 => "0000000010000000001000101000000100",
			6868 => "11111110111000110110110000011001",
			6869 => "00000001000110000110110000011001",
			6870 => "0000000000000000000010101000001000",
			6871 => "0000001110000000000111010100000100",
			6872 => "00000000000110100110110000011001",
			6873 => "00000100011011010110110000011001",
			6874 => "00000001010100000110110000011001",
			6875 => "0000000101000000000111111100000100",
			6876 => "11111110001111010110110000011001",
			6877 => "00000000011010010110110000011001",
			6878 => "0000000100000000000100001100010000",
			6879 => "0000001101000000001110110000000100",
			6880 => "11111110001000010110110000011001",
			6881 => "0000000111000000000101100100001000",
			6882 => "0000000000000000001010101100000100",
			6883 => "00000000010010010110110000011001",
			6884 => "00000010010000010110110000011001",
			6885 => "00000111100011000110110000011001",
			6886 => "0000001100000000001000111000001100",
			6887 => "0000000101000000000100001000000100",
			6888 => "11111110011101100110110000011001",
			6889 => "0000000100000000001110001000000100",
			6890 => "00000010100010100110110000011001",
			6891 => "11111111010100000110110000011001",
			6892 => "0000000110000000001111000000000100",
			6893 => "11111110011000010110110000011001",
			6894 => "0000000111000000001100101000000100",
			6895 => "00000001101101100110110000011001",
			6896 => "11111110111110010110110000011001",
			6897 => "0000000001000000001111000000100100",
			6898 => "0000000111000000000101100100001100",
			6899 => "0000000010000000000011001100001000",
			6900 => "0000001011000000000000110100000100",
			6901 => "00000001110001000110110000011001",
			6902 => "11111110011001100110110000011001",
			6903 => "00000010110110110110110000011001",
			6904 => "0000000001000000000001111000001100",
			6905 => "0000001010000000001010110000001000",
			6906 => "0000001101000000000111010100000100",
			6907 => "00000001011100010110110000011001",
			6908 => "00010000000001010110110000011001",
			6909 => "11111110010111110110110000011001",
			6910 => "0000001101000000001010000100000100",
			6911 => "11111110010111010110110000011001",
			6912 => "0000000101000000001110110100000100",
			6913 => "00000111101001100110110000011001",
			6914 => "11111110011100100110110000011001",
			6915 => "0000000010000000000011110100000100",
			6916 => "11111110011100010110110000011001",
			6917 => "00000010101100110110110000011001",
			6918 => "0000001110000000001110101101101100",
			6919 => "0000001011000000001110001101001000",
			6920 => "0000001101000000001001001000110000",
			6921 => "0000000100000000000011001100010100",
			6922 => "0000000010000000001100010100001000",
			6923 => "0000000011000000000100000100000100",
			6924 => "11111111101101000110110111011101",
			6925 => "00000000011101010110110111011101",
			6926 => "0000001000000000001001101000000100",
			6927 => "00000000000000000110110111011101",
			6928 => "0000000000000000000011010000000100",
			6929 => "11111110100010110110110111011101",
			6930 => "00000000000000000110110111011101",
			6931 => "0000000011000000001001110100001100",
			6932 => "0000001010000000000001010100000100",
			6933 => "11111110111010000110110111011101",
			6934 => "0000001011000000001001110000000100",
			6935 => "00000000000000000110110111011101",
			6936 => "00000000100111000110110111011101",
			6937 => "0000001100000000000100000000001000",
			6938 => "0000001101000000001110110000000100",
			6939 => "00000000000000000110110111011101",
			6940 => "00000000111110010110110111011101",
			6941 => "0000001000000000001010101100000100",
			6942 => "11111111010000100110110111011101",
			6943 => "00000000000011110110110111011101",
			6944 => "0000000000000000000011010000001000",
			6945 => "0000000110000000001011001100000100",
			6946 => "00000000000000000110110111011101",
			6947 => "00000001011010000110110111011101",
			6948 => "0000001110000000000100000100001000",
			6949 => "0000000011000000000100000100000100",
			6950 => "00000000000000000110110111011101",
			6951 => "00000001001001010110110111011101",
			6952 => "0000000110000000000100111100000100",
			6953 => "11111110111111000110110111011101",
			6954 => "00000000010001100110110111011101",
			6955 => "0000000000000000000011010000010000",
			6956 => "0000001100000000000100000000000100",
			6957 => "00000000000000000110110111011101",
			6958 => "0000000011000000000001001000001000",
			6959 => "0000000100000000001000101000000100",
			6960 => "00000000000000000110110111011101",
			6961 => "11111101111101000110110111011101",
			6962 => "00000000000000000110110111011101",
			6963 => "0000001101000000000001101000001000",
			6964 => "0000000011000000000010001000000100",
			6965 => "00000000000000000110110111011101",
			6966 => "00000001000110000110110111011101",
			6967 => "0000001010000000000110011100000100",
			6968 => "11111110110111010110110111011101",
			6969 => "0000000011000000000010110100000100",
			6970 => "00000000000000000110110111011101",
			6971 => "11111111110001110110110111011101",
			6972 => "0000000100000000001000001001000000",
			6973 => "0000000110000000000100111100100000",
			6974 => "0000001100000000000000001100001000",
			6975 => "0000000101000000000001101000000100",
			6976 => "00000000000000000110110111011101",
			6977 => "11111110110000110110110111011101",
			6978 => "0000001001000000001010100100001100",
			6979 => "0000001000000000000101000100001000",
			6980 => "0000001001000000000101010000000100",
			6981 => "00000000100101100110110111011101",
			6982 => "00000000000000110110110111011101",
			6983 => "00000001001101100110110111011101",
			6984 => "0000000100000000000110111000000100",
			6985 => "00000000000000000110110111011101",
			6986 => "0000001001000000001010100100000100",
			6987 => "00000000000000000110110111011101",
			6988 => "11111111001101100110110111011101",
			6989 => "0000001101000000000111111100000100",
			6990 => "00000001011011100110110111011101",
			6991 => "0000001111000000001000110100001100",
			6992 => "0000000010000000000011000000000100",
			6993 => "00000000010011000110110111011101",
			6994 => "0000001011000000000100010000000100",
			6995 => "00000000000000000110110111011101",
			6996 => "11111111000101010110110111011101",
			6997 => "0000001011000000001110101100001000",
			6998 => "0000001001000000000011101000000100",
			6999 => "00000001001100100110110111011101",
			7000 => "00000000000000000110110111011101",
			7001 => "0000001001000000000011101000000100",
			7002 => "11111111110110110110110111011101",
			7003 => "00000000010011000110110111011101",
			7004 => "0000001000000000001011010100011100",
			7005 => "0000000011000000000010010100001100",
			7006 => "0000000110000000000100111100000100",
			7007 => "00000000000000000110110111011101",
			7008 => "0000001110000000000110111000000100",
			7009 => "11111110010001010110110111011101",
			7010 => "00000000000000000110110111011101",
			7011 => "0000000101000000001110010000001000",
			7012 => "0000000000000000001101010000000100",
			7013 => "00000000000000000110110111011101",
			7014 => "00000000110100110110110111011101",
			7015 => "0000001001000000000100101100000100",
			7016 => "00000000000000000110110111011101",
			7017 => "11111111110111000110110111011101",
			7018 => "0000001100000000000011011100000100",
			7019 => "11111111010000100110110111011101",
			7020 => "0000001100000000000000001100001000",
			7021 => "0000000100000000000010111000000100",
			7022 => "00000000000000000110110111011101",
			7023 => "00000001001110000110110111011101",
			7024 => "0000001110000000000011010100001000",
			7025 => "0000001000000000001111001000000100",
			7026 => "00000000100000110110110111011101",
			7027 => "11111111010100010110110111011101",
			7028 => "0000000000000000001100001000000100",
			7029 => "00000001000010000110110111011101",
			7030 => "00000000000000000110110111011101",
			7031 => "0000001011000000000011011100010100",
			7032 => "0000000010000000000111011000000100",
			7033 => "11111110100001000110111100010001",
			7034 => "0000000010000000000000010000001100",
			7035 => "0000001001000000001101101000001000",
			7036 => "0000001001000000001100110100000100",
			7037 => "00000000000000000110111100010001",
			7038 => "00000000010001000110111100010001",
			7039 => "00000000000000000110111100010001",
			7040 => "11111111100111010110111100010001",
			7041 => "0000000111000000001000111000100100",
			7042 => "0000001111000000000101001000010100",
			7043 => "0000000010000000001100010100000100",
			7044 => "11111111001001000110111100010001",
			7045 => "0000001100000000001000111000001100",
			7046 => "0000001011000000000011011100000100",
			7047 => "00000000000000000110111100010001",
			7048 => "0000001010000000000001010000000100",
			7049 => "00000000000000000110111100010001",
			7050 => "00000001100010000110111100010001",
			7051 => "00000000000000000110111100010001",
			7052 => "0000000010000000001111010100001100",
			7053 => "0000000011000000000000011100000100",
			7054 => "11111111010110000110111100010001",
			7055 => "0000000000000000000010011000000100",
			7056 => "11111111111110100110111100010001",
			7057 => "00000001010101100110111100010001",
			7058 => "11111110101110110110111100010001",
			7059 => "0000001001000000000111101001000000",
			7060 => "0000000010000000000010000000100000",
			7061 => "0000000010000000000011001000010000",
			7062 => "0000001001000000001011111100001000",
			7063 => "0000001010000000001010100000000100",
			7064 => "00000000000000000110111100010001",
			7065 => "11111111001000110110111100010001",
			7066 => "0000000101000000001000011000000100",
			7067 => "00000000000011110110111100010001",
			7068 => "00000000000000000110111100010001",
			7069 => "0000000111000000001001110000001000",
			7070 => "0000000011000000001001110100000100",
			7071 => "00000000000000000110111100010001",
			7072 => "00000001011010010110111100010001",
			7073 => "0000000101000000000111010000000100",
			7074 => "11111111001100100110111100010001",
			7075 => "00000000111111110110111100010001",
			7076 => "0000000101000000001001001000010000",
			7077 => "0000001101000000001001001000001000",
			7078 => "0000000100000000001110111000000100",
			7079 => "11111110101010110110111100010001",
			7080 => "11111111111000100110111100010001",
			7081 => "0000000000000000000010111100000100",
			7082 => "11111110110101010110111100010001",
			7083 => "00000000101100100110111100010001",
			7084 => "0000000010000000001010000100001000",
			7085 => "0000001101000000000110100100000100",
			7086 => "00000000000000000110111100010001",
			7087 => "11111101111101000110111100010001",
			7088 => "0000001100000000001001110000000100",
			7089 => "00000000101110010110111100010001",
			7090 => "11111111001010100110111100010001",
			7091 => "0000000101000000001010011100001000",
			7092 => "0000001110000000000010011100000100",
			7093 => "00000001101101110110111100010001",
			7094 => "11111111011100110110111100010001",
			7095 => "0000000011000000001001011100001100",
			7096 => "0000000010000000001101000100001000",
			7097 => "0000001111000000000101110100000100",
			7098 => "00000000000000000110111100010001",
			7099 => "00000000101011010110111100010001",
			7100 => "11111110011001010110111100010001",
			7101 => "0000000111000000001100101000001000",
			7102 => "0000000000000000000011111100000100",
			7103 => "00000000000000000110111100010001",
			7104 => "00000001101110110110111100010001",
			7105 => "0000000111000000000111001000000100",
			7106 => "11111110010011010110111100010001",
			7107 => "00000000000001000110111100010001",
			7108 => "0000000110000000001001100101010000",
			7109 => "0000000101000000000111001000000100",
			7110 => "11111110100101010111000001101101",
			7111 => "0000000001000000001001111000010000",
			7112 => "0000001111000000000001000000001100",
			7113 => "0000001000000000000111000100000100",
			7114 => "00000000000000000111000001101101",
			7115 => "0000000011000000001001110100000100",
			7116 => "00000000000000000111000001101101",
			7117 => "00000001100011100111000001101101",
			7118 => "11111111101000000111000001101101",
			7119 => "0000001000000000001010110000011100",
			7120 => "0000000100000000001011101100010000",
			7121 => "0000001101000000001111010000001000",
			7122 => "0000000000000000001011010100000100",
			7123 => "00000000100010110111000001101101",
			7124 => "11111111000101110111000001101101",
			7125 => "0000001101000000000100101000000100",
			7126 => "11111110101000100111000001101101",
			7127 => "00000000000000000111000001101101",
			7128 => "0000000110000000001101011000000100",
			7129 => "00000000000000000111000001101101",
			7130 => "0000000011000000001111010100000100",
			7131 => "00000000000000000111000001101101",
			7132 => "00000001100100100111000001101101",
			7133 => "0000001111000000000101110000010000",
			7134 => "0000001110000000001010001100001000",
			7135 => "0000001001000000001101011100000100",
			7136 => "00000000000000000111000001101101",
			7137 => "11111111001001010111000001101101",
			7138 => "0000000100000000000110111000000100",
			7139 => "00000000000000000111000001101101",
			7140 => "00000000110100100111000001101101",
			7141 => "0000001100000000001010111000001000",
			7142 => "0000001100000000000100000000000100",
			7143 => "11111111111101110111000001101101",
			7144 => "11111110011110110111000001101101",
			7145 => "0000001101000000000010011100000100",
			7146 => "11111111001010000111000001101101",
			7147 => "00000000011101100111000001101101",
			7148 => "0000001101000000000110100100110000",
			7149 => "0000001011000000001100101100100100",
			7150 => "0000001101000000001001001000011100",
			7151 => "0000001011000000000101101100010000",
			7152 => "0000001001000000001111001100001000",
			7153 => "0000001011000000001000111000000100",
			7154 => "00000000000000000111000001101101",
			7155 => "00000001010100110111000001101101",
			7156 => "0000000000000000000000110000000100",
			7157 => "00000000001110100111000001101101",
			7158 => "11111110110110010111000001101101",
			7159 => "0000001101000000001000000000001000",
			7160 => "0000000101000000000100011000000100",
			7161 => "11111111100110000111000001101101",
			7162 => "11111110010101000111000001101101",
			7163 => "00000000000000000111000001101101",
			7164 => "0000000000000000000010111100000100",
			7165 => "00000000000000000111000001101101",
			7166 => "00000001011100010111000001101101",
			7167 => "0000000000000000000010011000000100",
			7168 => "00000000000000000111000001101101",
			7169 => "0000001111000000001110000100000100",
			7170 => "00000000000000000111000001101101",
			7171 => "00000001110011110111000001101101",
			7172 => "0000001001000000001011111100010000",
			7173 => "0000001010000000001100011100000100",
			7174 => "11111110000000110111000001101101",
			7175 => "0000001101000000001000011000001000",
			7176 => "0000000011000000000101110100000100",
			7177 => "00000000000000000111000001101101",
			7178 => "00000000110001010111000001101101",
			7179 => "00000000000000000111000001101101",
			7180 => "0000000101000000000001101000001000",
			7181 => "0000000110000000001111000000000100",
			7182 => "00000000010100010111000001101101",
			7183 => "00000001100100000111000001101101",
			7184 => "0000001110000000001110101000001000",
			7185 => "0000000110000000001001100100000100",
			7186 => "00000000000000000111000001101101",
			7187 => "11111110011001010111000001101101",
			7188 => "0000001100000000000110000100001000",
			7189 => "0000001000000000001111001000000100",
			7190 => "11111111101100010111000001101101",
			7191 => "00000001011110000111000001101101",
			7192 => "0000000100000000001000001000000100",
			7193 => "00000000010100000111000001101101",
			7194 => "11111111011111000111000001101101",
			7195 => "0000001011000000000011011100010000",
			7196 => "0000000010000000000111011000000100",
			7197 => "11111110011010110111000110110001",
			7198 => "0000001101000000000001111100000100",
			7199 => "11111110110001010111000110110001",
			7200 => "0000001101000000001101010100000100",
			7201 => "00000000110011100111000110110001",
			7202 => "00000000000000000111000110110001",
			7203 => "0000000100000000000011000001000000",
			7204 => "0000000010000000000111010100100000",
			7205 => "0000001111000000001010000100011100",
			7206 => "0000001111000000001111010100001100",
			7207 => "0000001010000000001001000100001000",
			7208 => "0000001101000000001111010000000100",
			7209 => "00000000001001110111000110110001",
			7210 => "11111110101000000111000110110001",
			7211 => "00000001011100100111000110110001",
			7212 => "0000000010000000001111010100001000",
			7213 => "0000000011000000001010000100000100",
			7214 => "00000010001010000111000110110001",
			7215 => "00000000000000000111000110110001",
			7216 => "0000001100000000001011000000000100",
			7217 => "11111111010000110111000110110001",
			7218 => "00000000011011100111000110110001",
			7219 => "11111110011101100111000110110001",
			7220 => "0000001110000000000111010100001100",
			7221 => "0000001111000000001000001100000100",
			7222 => "11111111001110110111000110110001",
			7223 => "0000000111000000000001101000000100",
			7224 => "00000001100101100111000110110001",
			7225 => "00000011111100110111000110110001",
			7226 => "0000000010000000000110101100001100",
			7227 => "0000000111000000000001101000000100",
			7228 => "11111110100001010111000110110001",
			7229 => "0000000001000000000001111000000100",
			7230 => "11111111100100100111000110110001",
			7231 => "00000000010001110111000110110001",
			7232 => "0000001010000000000011101000000100",
			7233 => "00000010000100000111000110110001",
			7234 => "11111111010011000111000110110001",
			7235 => "0000001100000000001000111100100100",
			7236 => "0000000000000000001111000100001100",
			7237 => "0000000000000000001111000100001000",
			7238 => "0000001000000000001001101000000100",
			7239 => "11111111010111110111000110110001",
			7240 => "00000000110110100111000110110001",
			7241 => "11111011011011010111000110110001",
			7242 => "0000000100000000001011100000010000",
			7243 => "0000000011000000000001101000001000",
			7244 => "0000001100000000000000101000000100",
			7245 => "00000000001100000111000110110001",
			7246 => "11111110001111010111000110110001",
			7247 => "0000000010000000000010000100000100",
			7248 => "00000001011100110111000110110001",
			7249 => "00000000000011000111000110110001",
			7250 => "0000000111000000001101100000000100",
			7251 => "00000001101101110111000110110001",
			7252 => "00000000000000000111000110110001",
			7253 => "0000000011000000000010000000011100",
			7254 => "0000001000000000000110001000010000",
			7255 => "0000000000000000001000101100001000",
			7256 => "0000001010000000001000100100000100",
			7257 => "11111111001110000111000110110001",
			7258 => "00000001010010110111000110110001",
			7259 => "0000000000000000000010111100000100",
			7260 => "11111110001100100111000110110001",
			7261 => "11111111101010010111000110110001",
			7262 => "0000000100000000001100001100000100",
			7263 => "00000001110011100111000110110001",
			7264 => "0000001100000000001100110000000100",
			7265 => "11111111110101010111000110110001",
			7266 => "11111110001010000111000110110001",
			7267 => "0000000111000000000001111100000100",
			7268 => "00000010000010100111000110110001",
			7269 => "0000000000000000001111000100001000",
			7270 => "0000000000000000000111000100000100",
			7271 => "11111111000111000111000110110001",
			7272 => "00000000100100000111000110110001",
			7273 => "0000001000000000001001101000000100",
			7274 => "11111100110011010111000110110001",
			7275 => "11111111101110100111000110110001",
			7276 => "0000000101000000000111100010001000",
			7277 => "0000000111000000001110110001001100",
			7278 => "0000001000000000000110001000011000",
			7279 => "0000001100000000000100000000001000",
			7280 => "0000000110000000001011001100000100",
			7281 => "00000000000000000111001101011101",
			7282 => "00000000000100010111001101011101",
			7283 => "0000001101000000001000000000000100",
			7284 => "00000000000000000111001101011101",
			7285 => "0000001000000000001001000100000100",
			7286 => "00000000000000000111001101011101",
			7287 => "0000000110000000001000010000000100",
			7288 => "11111111000011010111001101011101",
			7289 => "00000000000000000111001101011101",
			7290 => "0000000011000000001011011100011100",
			7291 => "0000001111000000001111010000010000",
			7292 => "0000000011000000001001110100001000",
			7293 => "0000001111000000000110100000000100",
			7294 => "00000000000000000111001101011101",
			7295 => "11111111010101010111001101011101",
			7296 => "0000000001000000000110101000000100",
			7297 => "00000000101000010111001101011101",
			7298 => "11111111111111100111001101011101",
			7299 => "0000000111000000001000111000000100",
			7300 => "00000000000000000111001101011101",
			7301 => "0000000110000000001111000000000100",
			7302 => "11111110110110000111001101011101",
			7303 => "00000000000000000111001101011101",
			7304 => "0000001111000000001001011100001000",
			7305 => "0000000101000000000110100100000100",
			7306 => "00000001001001100111001101011101",
			7307 => "00000000000000000111001101011101",
			7308 => "0000000110000000000100111100001000",
			7309 => "0000000010000000001100000000000100",
			7310 => "00000000000000000111001101011101",
			7311 => "11111111011101010111001101011101",
			7312 => "0000000010000000000101000000000100",
			7313 => "00000000100110110111001101011101",
			7314 => "00000000000000000111001101011101",
			7315 => "0000001111000000000110111100010100",
			7316 => "0000001100000000001010111000010000",
			7317 => "0000000010000000001110110100001100",
			7318 => "0000001101000000000111100000001000",
			7319 => "0000001111000000001110101000000100",
			7320 => "00000000000000000111001101011101",
			7321 => "00000000001110010111001101011101",
			7322 => "00000000000000000111001101011101",
			7323 => "00000000000000000111001101011101",
			7324 => "11111111010101110111001101011101",
			7325 => "0000000111000000000001101000011000",
			7326 => "0000000111000000001001001000001100",
			7327 => "0000001100000000000100011000001000",
			7328 => "0000001100000000000100001000000100",
			7329 => "00000000000000000111001101011101",
			7330 => "00000000101010010111001101011101",
			7331 => "00000000000000000111001101011101",
			7332 => "0000001111000000001010000100000100",
			7333 => "00000000000000000111001101011101",
			7334 => "0000000111000000000110100100000100",
			7335 => "11111111011110010111001101011101",
			7336 => "00000000000000000111001101011101",
			7337 => "0000001111000000001010000100000100",
			7338 => "00000000000000000111001101011101",
			7339 => "0000001011000000000101100100000100",
			7340 => "00000000000000000111001101011101",
			7341 => "0000001011000000000010001000000100",
			7342 => "00000000110111000111001101011101",
			7343 => "00000000000000000111001101011101",
			7344 => "0000000011000000000110111000011000",
			7345 => "0000000001000000000100110100001100",
			7346 => "0000000111000000000101100100001000",
			7347 => "0000001001000000001010100100000100",
			7348 => "11111110110101000111001101011101",
			7349 => "00000000000000000111001101011101",
			7350 => "00000000000000000111001101011101",
			7351 => "0000000111000000001000011000000100",
			7352 => "00000000001110100111001101011101",
			7353 => "0000000111000000001111011100000100",
			7354 => "11111111110100000111001101011101",
			7355 => "00000000000000000111001101011101",
			7356 => "0000000101000000000111111100001000",
			7357 => "0000000001000000000100110100000100",
			7358 => "00000000000000000111001101011101",
			7359 => "00000000101111000111001101011101",
			7360 => "0000000011000000000010111000011000",
			7361 => "0000000110000000001000010000001100",
			7362 => "0000001100000000001111011100000100",
			7363 => "00000000000000000111001101011101",
			7364 => "0000000111000000001011011100000100",
			7365 => "00000000000000000111001101011101",
			7366 => "00000000010111110111001101011101",
			7367 => "0000001010000000001000010100000100",
			7368 => "00000000000000000111001101011101",
			7369 => "0000000101000000001100010000000100",
			7370 => "11111110110100000111001101011101",
			7371 => "00000000000000000111001101011101",
			7372 => "0000001100000000000111010000001100",
			7373 => "0000000001000000001010011000000100",
			7374 => "00000000000000000111001101011101",
			7375 => "0000001000000000001001101000000100",
			7376 => "00000000000000000111001101011101",
			7377 => "00000000101110000111001101011101",
			7378 => "0000000111000000000000110100000100",
			7379 => "11111111010010100111001101011101",
			7380 => "0000000110000000000100101100000100",
			7381 => "00000000100001010111001101011101",
			7382 => "00000000000000000111001101011101",
			7383 => "0000001110000000001110101101101100",
			7384 => "0000001111000000001001010000110100",
			7385 => "0000000011000000001010001100100100",
			7386 => "0000000010000000001110110100001100",
			7387 => "0000000100000000001110111000001000",
			7388 => "0000001101000000000111010000000100",
			7389 => "11111110110100110111010100110001",
			7390 => "00000000000000000111010100110001",
			7391 => "00000000000000000111010100110001",
			7392 => "0000000110000000001011001100001100",
			7393 => "0000000001000000000010001100001000",
			7394 => "0000000101000000001010111000000100",
			7395 => "00000000000000000111010100110001",
			7396 => "00000000000011110111010100110001",
			7397 => "11111111000001000111010100110001",
			7398 => "0000000011000000001001110100001000",
			7399 => "0000000101000000001110110000000100",
			7400 => "00000000000010110111010100110001",
			7401 => "11111111110001010111010100110001",
			7402 => "00000001001101000111010100110001",
			7403 => "0000000010000000001100010100000100",
			7404 => "00000000000000000111010100110001",
			7405 => "0000001100000000000100000000000100",
			7406 => "00000000000000000111010100110001",
			7407 => "0000000000000000001100001000000100",
			7408 => "00000001010000000111010100110001",
			7409 => "00000000000000000111010100110001",
			7410 => "0000000100000000000010111000011000",
			7411 => "0000001100000000000100000000001000",
			7412 => "0000000110000000001001100100000100",
			7413 => "00000000000000000111010100110001",
			7414 => "00000000100110110111010100110001",
			7415 => "0000000001000000000111100100001000",
			7416 => "0000000110000000001011001100000100",
			7417 => "00000000000000000111010100110001",
			7418 => "11111110110000000111010100110001",
			7419 => "0000000110000000001001100100000100",
			7420 => "11111111111110010111010100110001",
			7421 => "00000000001110000111010100110001",
			7422 => "0000000000000000000000110000001100",
			7423 => "0000000110000000001001100100000100",
			7424 => "00000000000000000111010100110001",
			7425 => "0000000101000000000110100100000100",
			7426 => "00000001001010010111010100110001",
			7427 => "00000000000000000111010100110001",
			7428 => "0000000110000000001111000000001000",
			7429 => "0000001010000000000001010100000100",
			7430 => "11111110111000000111010100110001",
			7431 => "00000000000000000111010100110001",
			7432 => "0000001010000000001100000100001000",
			7433 => "0000000011000000000010001000000100",
			7434 => "00000000000000000111010100110001",
			7435 => "00000000100101000111010100110001",
			7436 => "00000000000000000111010100110001",
			7437 => "0000000101000000000111100000110100",
			7438 => "0000000011000000000010000100011100",
			7439 => "0000001111000000001111100100011000",
			7440 => "0000001010000000000001010000001100",
			7441 => "0000000010000000000111011000001000",
			7442 => "0000001110000000000101001000000100",
			7443 => "00000000110110000111010100110001",
			7444 => "11111111110000100111010100110001",
			7445 => "11111110111001110111010100110001",
			7446 => "0000001001000000000001111000000100",
			7447 => "00000000000000000111010100110001",
			7448 => "0000001110000000000111111100000100",
			7449 => "00000001011010010111010100110001",
			7450 => "00000000000000000111010100110001",
			7451 => "11111110110110110111010100110001",
			7452 => "0000001000000000000111000000010100",
			7453 => "0000000010000000001000101000010000",
			7454 => "0000001001000000000111101100001000",
			7455 => "0000001111000000000110111100000100",
			7456 => "00000000000000000111010100110001",
			7457 => "00000000110000110111010100110001",
			7458 => "0000000001000000000001111000000100",
			7459 => "11111111010010010111010100110001",
			7460 => "00000000001011000111010100110001",
			7461 => "00000001001110000111010100110001",
			7462 => "11111111111110010111010100110001",
			7463 => "0000000101000000000010011100011000",
			7464 => "0000000101000000001111010000001100",
			7465 => "0000000000000000001010101100000100",
			7466 => "11111111000000010111010100110001",
			7467 => "0000000100000000001001001100000100",
			7468 => "00000001000100110111010100110001",
			7469 => "00000000000000000111010100110001",
			7470 => "0000001001000000000010101100001000",
			7471 => "0000000011000000000110111000000100",
			7472 => "11111110001110000111010100110001",
			7473 => "00000000000000000111010100110001",
			7474 => "00000000000000000111010100110001",
			7475 => "0000001110000000001000101000010100",
			7476 => "0000001101000000000011001000000100",
			7477 => "00000000000000000111010100110001",
			7478 => "0000001100000000000001101000001000",
			7479 => "0000000000000000001011010100000100",
			7480 => "00000000000000000111010100110001",
			7481 => "00000001001110110111010100110001",
			7482 => "0000000001000000000101011100000100",
			7483 => "00000000010000110111010100110001",
			7484 => "11111111111000010111010100110001",
			7485 => "0000000101000000000011001000010000",
			7486 => "0000001110000000001011110000001000",
			7487 => "0000000011000000000010010100000100",
			7488 => "00000000000000000111010100110001",
			7489 => "11111110110111110111010100110001",
			7490 => "0000000101000000001110010000000100",
			7491 => "00000000011011110111010100110001",
			7492 => "11111111010111010111010100110001",
			7493 => "0000000011000000000100001100001000",
			7494 => "0000000001000000001101011000000100",
			7495 => "00000000100011010111010100110001",
			7496 => "00000000000000000111010100110001",
			7497 => "0000001110000000001011100000000100",
			7498 => "11111111010100010111010100110001",
			7499 => "00000000000000000111010100110001",
			7500 => "0000001011000000000011011100001000",
			7501 => "0000000110000000001001100100000100",
			7502 => "11111110011011000111011001010101",
			7503 => "11111111111110110111011001010101",
			7504 => "0000000100000000000011000000110000",
			7505 => "0000000011000000000111110000010000",
			7506 => "0000001001000000001011111100001000",
			7507 => "0000000111000000001101111000000100",
			7508 => "11111110101101100111011001010101",
			7509 => "00000000000000000111011001010101",
			7510 => "0000001101000000001010001100000100",
			7511 => "00000000001101110111011001010101",
			7512 => "00000000000000000111011001010101",
			7513 => "0000001010000000001000100100011100",
			7514 => "0000001011000000000000011100010000",
			7515 => "0000001101000000000101110100001000",
			7516 => "0000000111000000001100101000000100",
			7517 => "00000000000000000111011001010101",
			7518 => "00000001111001010111011001010101",
			7519 => "0000000011000000001100000000000100",
			7520 => "11111110101110000111011001010101",
			7521 => "00000000000000000111011001010101",
			7522 => "0000000001000000000101011100000100",
			7523 => "11111110110011010111011001010101",
			7524 => "0000000110000000001001100100000100",
			7525 => "00000001001110010111011001010101",
			7526 => "11111111101000010111011001010101",
			7527 => "00000001101011000111011001010101",
			7528 => "0000000110000000001001100100111100",
			7529 => "0000000001000000000110101000011100",
			7530 => "0000000011000000001010011100010000",
			7531 => "0000000100000000001111100000001000",
			7532 => "0000001110000000001000000000000100",
			7533 => "11111110001111100111011001010101",
			7534 => "00000000000000000111011001010101",
			7535 => "0000001100000000000100000000000100",
			7536 => "00000001001001000111011001010101",
			7537 => "11111110111110110111011001010101",
			7538 => "0000000010000000001100000000001000",
			7539 => "0000000000000000000011010000000100",
			7540 => "11111111000111110111011001010101",
			7541 => "00000010000001100111011001010101",
			7542 => "11111110101011110111011001010101",
			7543 => "0000000100000000000011110000010000",
			7544 => "0000000000000000000010111100001000",
			7545 => "0000001101000000000110100100000100",
			7546 => "11111101110100100111011001010101",
			7547 => "00000000000000000111011001010101",
			7548 => "0000000111000000001001110000000100",
			7549 => "00000000000000000111011001010101",
			7550 => "00000001101000110111011001010101",
			7551 => "0000001011000000000110000100001000",
			7552 => "0000001001000000001001011000000100",
			7553 => "11111110011011000111011001010101",
			7554 => "00000000000000000111011001010101",
			7555 => "0000000000000000001101010000000100",
			7556 => "00000000000000000111011001010101",
			7557 => "11111101100011110111011001010101",
			7558 => "0000001100000000001000111100001100",
			7559 => "0000001100000000000000101000001000",
			7560 => "0000000001000000000110101000000100",
			7561 => "00000001101011010111011001010101",
			7562 => "11111110011011010111011001010101",
			7563 => "00000001100111100111011001010101",
			7564 => "0000000000000000001001110000010000",
			7565 => "0000000001000000001101011000001000",
			7566 => "0000001001000000000111101100000100",
			7567 => "11111111111011000111011001010101",
			7568 => "00000000100011110111011001010101",
			7569 => "0000000000000000000000111000000100",
			7570 => "11111110101001110111011001010101",
			7571 => "00000000100000100111011001010101",
			7572 => "11111110001001110111011001010101",
			7573 => "0000001110000000001110101101100000",
			7574 => "0000001011000000001110001101000100",
			7575 => "0000001101000000001001001000101100",
			7576 => "0000000101000000000100011000011100",
			7577 => "0000001101000000001110110000001100",
			7578 => "0000000100000000000001101100000100",
			7579 => "11111110111100110111100000101001",
			7580 => "0000001011000000001001110000000100",
			7581 => "00000000000000000111100000101001",
			7582 => "00000000100001000111100000101001",
			7583 => "0000001111000000001001010000001000",
			7584 => "0000000111000000001000111000000100",
			7585 => "00000000000000000111100000101001",
			7586 => "00000000111101000111100000101001",
			7587 => "0000000111000000001000111000000100",
			7588 => "00000000000000000111100000101001",
			7589 => "11111111001111000111100000101001",
			7590 => "0000000010000000000111011000001000",
			7591 => "0000001100000000000100000000000100",
			7592 => "00000000000000000111100000101001",
			7593 => "11111110101010010111100000101001",
			7594 => "0000000010000000001111010100000100",
			7595 => "00000000000000000111100000101001",
			7596 => "11111111111110000111100000101001",
			7597 => "0000000000000000000011010000001000",
			7598 => "0000001111000000001111010000000100",
			7599 => "00000000000000000111100000101001",
			7600 => "00000001011011110111100000101001",
			7601 => "0000001110000000000100000100001000",
			7602 => "0000000111000000001101100000000100",
			7603 => "00000001001110010111100000101001",
			7604 => "00000000000000000111100000101001",
			7605 => "0000000111000000001101100000000100",
			7606 => "11111110101100100111100000101001",
			7607 => "00000000101100000111100000101001",
			7608 => "0000000001000000000110101000001000",
			7609 => "0000001010000000000110011100000100",
			7610 => "11111101110100000111100000101001",
			7611 => "00000000000000000111100000101001",
			7612 => "0000000101000000001001001000001000",
			7613 => "0000001111000000000100101000000100",
			7614 => "11111111011010100111100000101001",
			7615 => "00000001010101000111100000101001",
			7616 => "0000001001000000000101011100000100",
			7617 => "00000000000000000111100000101001",
			7618 => "0000000100000000001000001100000100",
			7619 => "00000000000000000111100000101001",
			7620 => "11111110100011010111100000101001",
			7621 => "0000000100000000001000001001001100",
			7622 => "0000001100000000001110001100010000",
			7623 => "0000001011000000000100001000001000",
			7624 => "0000001010000000000110011000000100",
			7625 => "00000000000000000111100000101001",
			7626 => "00000000101010110111100000101001",
			7627 => "0000000001000000001001011000000100",
			7628 => "11111110110111100111100000101001",
			7629 => "00000000000000000111100000101001",
			7630 => "0000001000000000000101000100100000",
			7631 => "0000001010000000000010101100010000",
			7632 => "0000000010000000000111011000001000",
			7633 => "0000001100000000001010111000000100",
			7634 => "00000000110001000111100000101001",
			7635 => "11111111010110010111100000101001",
			7636 => "0000000001000000000001000100000100",
			7637 => "00000000000000000111100000101001",
			7638 => "00000001000110000111100000101001",
			7639 => "0000000100000000001011101100001000",
			7640 => "0000000101000000000010110100000100",
			7641 => "00000000000000000111100000101001",
			7642 => "11111110111110000111100000101001",
			7643 => "0000000100000000000011000000000100",
			7644 => "00000000011011010111100000101001",
			7645 => "11111111101010110111100000101001",
			7646 => "0000000111000000000110110100001100",
			7647 => "0000000001000000001101011000001000",
			7648 => "0000000000000000000001110100000100",
			7649 => "00000000000000000111100000101001",
			7650 => "00000000111011100111100000101001",
			7651 => "00000000000000000111100000101001",
			7652 => "0000001111000000000110001100001000",
			7653 => "0000001001000000000011101000000100",
			7654 => "11111111100100110111100000101001",
			7655 => "00000000000000000111100000101001",
			7656 => "0000001110000000001110100100000100",
			7657 => "00000000000110100111100000101001",
			7658 => "00000000000000000111100000101001",
			7659 => "0000001000000000001011010100101000",
			7660 => "0000000000000000001111000100011100",
			7661 => "0000001001000000000100101100001100",
			7662 => "0000001010000000000110011000001000",
			7663 => "0000000100000000000010111000000100",
			7664 => "00000000000000000111100000101001",
			7665 => "00000001000000110111100000101001",
			7666 => "00000000000000000111100000101001",
			7667 => "0000000000000000001101010000001000",
			7668 => "0000001100000000001011000000000100",
			7669 => "00000000000000000111100000101001",
			7670 => "11111111010110110111100000101001",
			7671 => "0000001001000000000000001000000100",
			7672 => "00000000000000000111100000101001",
			7673 => "00000000010101000111100000101001",
			7674 => "0000001110000000001011110000000100",
			7675 => "11111110001010110111100000101001",
			7676 => "0000000111000000000001011000000100",
			7677 => "00000000000111110111100000101001",
			7678 => "00000000000000000111100000101001",
			7679 => "0000001100000000000011011100000100",
			7680 => "11111111001101010111100000101001",
			7681 => "0000000111000000000100001000000100",
			7682 => "00000001011001110111100000101001",
			7683 => "0000001110000000000011010100001000",
			7684 => "0000001010000000000110011100000100",
			7685 => "00000000001101110111100000101001",
			7686 => "11111111000111000111100000101001",
			7687 => "0000000000000000001100001000000100",
			7688 => "00000001000101010111100000101001",
			7689 => "00000000000000000111100000101001",
			7690 => "0000000011000000001001110100100000",
			7691 => "0000000001000000000111100100011100",
			7692 => "0000000010000000001001100000000100",
			7693 => "11111110011001000111100101111101",
			7694 => "0000001100000000000100000000001100",
			7695 => "0000001000000000001000110000000100",
			7696 => "11111110011010100111100101111101",
			7697 => "0000000101000000000000001100000100",
			7698 => "11111110100111100111100101111101",
			7699 => "00000010000010100111100101111101",
			7700 => "0000000111000000001000111000001000",
			7701 => "0000000111000000001000111000000100",
			7702 => "11111110110010000111100101111101",
			7703 => "00000000000000000111100101111101",
			7704 => "11111110010110100111100101111101",
			7705 => "00000001110101110111100101111101",
			7706 => "0000001100000000001000011001100100",
			7707 => "0000001000000000000001110000110000",
			7708 => "0000000000000000001100000100010000",
			7709 => "0000001001000000000101010000001100",
			7710 => "0000001101000000000100010000001000",
			7711 => "0000000001000000001011101000000100",
			7712 => "11111110100100100111100101111101",
			7713 => "00000011000010110111100101111101",
			7714 => "11111110011010000111100101111101",
			7715 => "00000001000110100111100101111101",
			7716 => "0000000101000000000111100000010000",
			7717 => "0000001011000000000100000100001000",
			7718 => "0000001110000000000110111100000100",
			7719 => "11111111001001000111100101111101",
			7720 => "00000001010011110111100101111101",
			7721 => "0000000111000000001001001000000100",
			7722 => "11111111011001100111100101111101",
			7723 => "00000001100101110111100101111101",
			7724 => "0000001001000000001001111100001000",
			7725 => "0000000101000000000101110000000100",
			7726 => "11111110011111000111100101111101",
			7727 => "00000001110101010111100101111101",
			7728 => "0000000000000000001010101100000100",
			7729 => "11111110100100100111100101111101",
			7730 => "00000000001010100111100101111101",
			7731 => "0000001001000000000111101100100000",
			7732 => "0000001100000000001000111000010000",
			7733 => "0000000101000000000111001000001000",
			7734 => "0000000100000000000011110100000100",
			7735 => "11111110010011100111100101111101",
			7736 => "00000000001001010111100101111101",
			7737 => "0000000001000000000111100100000100",
			7738 => "00000001000000100111100101111101",
			7739 => "00000001110111010111100101111101",
			7740 => "0000000011000000001110010000001000",
			7741 => "0000000111000000000101101100000100",
			7742 => "00000000010000010111100101111101",
			7743 => "11111110011111010111100101111101",
			7744 => "0000001100000000000110000100000100",
			7745 => "00000010000010100111100101111101",
			7746 => "00000000000000000111100101111101",
			7747 => "0000001011000000001011110100001000",
			7748 => "0000000100000000001110111000000100",
			7749 => "00000001110111110111100101111101",
			7750 => "00000000000000000111100101111101",
			7751 => "0000001110000000001011110000000100",
			7752 => "11111110000110100111100101111101",
			7753 => "0000001100000000001001110100000100",
			7754 => "11111110110101110111100101111101",
			7755 => "00000001111000110111100101111101",
			7756 => "0000001001000000001000010100100000",
			7757 => "0000001000000000001011010100011100",
			7758 => "0000001101000000001010000100010000",
			7759 => "0000000001000000000001111000001000",
			7760 => "0000000001000000000001111000000100",
			7761 => "11111111111001100111100101111101",
			7762 => "00000110010111010111100101111101",
			7763 => "0000001101000000000110111100000100",
			7764 => "11111110011001100111100101111101",
			7765 => "11111111011111110111100101111101",
			7766 => "0000001110000000001000011100000100",
			7767 => "00000011111010000111100101111101",
			7768 => "0000000111000000000111110000000100",
			7769 => "11111110100011010111100101111101",
			7770 => "00000011111010100111100101111101",
			7771 => "11111110011001110111100101111101",
			7772 => "0000000000000000000010111100000100",
			7773 => "11111111001100100111100101111101",
			7774 => "00000001100100100111100101111101",
			7775 => "0000000110000000001011001101001100",
			7776 => "0000001001000000001000010000100100",
			7777 => "0000000110000000001101011000011000",
			7778 => "0000000110000000001001011000001000",
			7779 => "0000000101000000000110100100000100",
			7780 => "11111110100010110111101100111001",
			7781 => "00000010011111010111101100111001",
			7782 => "0000000100000000000101110000001100",
			7783 => "0000001010000000001001111100000100",
			7784 => "11111110011110100111101100111001",
			7785 => "0000000101000000001110101100000100",
			7786 => "00000011011111000111101100111001",
			7787 => "11111111011011000111101100111001",
			7788 => "11111110011000110111101100111001",
			7789 => "0000000011000000001010001100000100",
			7790 => "11111110011100000111101100111001",
			7791 => "0000000010000000000010000100000100",
			7792 => "00000011010010000111101100111001",
			7793 => "11111110101100010111101100111001",
			7794 => "0000000111000000001001001000001000",
			7795 => "0000001110000000000111111100000100",
			7796 => "00000001001101010111101100111001",
			7797 => "11111110010111100111101100111001",
			7798 => "0000000111000000000110100100010000",
			7799 => "0000001110000000000010000000000100",
			7800 => "11111110110100000111101100111001",
			7801 => "0000000001000000000001000100000100",
			7802 => "11111111001010100111101100111001",
			7803 => "0000000111000000000110100100000100",
			7804 => "00000100010111110111101100111001",
			7805 => "00000010100110010111101100111001",
			7806 => "0000000000000000001001101000001000",
			7807 => "0000001011000000000101100100000100",
			7808 => "00000001011000110111101100111001",
			7809 => "11111110011101000111101100111001",
			7810 => "0000001100000000001001110100000100",
			7811 => "00000011101000100111101100111001",
			7812 => "11111110100111010111101100111001",
			7813 => "0000001100000000001000011001101000",
			7814 => "0000000110000000001000010000111100",
			7815 => "0000000111000000001101100000011100",
			7816 => "0000000001000000000110101000010000",
			7817 => "0000001111000000000111111100001000",
			7818 => "0000000101000000000111001000000100",
			7819 => "11111111111011000111101100111001",
			7820 => "00000001110010000111101100111001",
			7821 => "0000000000000000000000111000000100",
			7822 => "11111101000111000111101100111001",
			7823 => "11111111111100100111101100111001",
			7824 => "0000000110000000001001100100000100",
			7825 => "11111111111100100111101100111001",
			7826 => "0000000001000000000111100100000100",
			7827 => "00000001100101110111101100111001",
			7828 => "00000010001010100111101100111001",
			7829 => "0000000011000000001100010000010000",
			7830 => "0000001011000000001101111000001000",
			7831 => "0000000001000000000111100100000100",
			7832 => "11111110110110000111101100111001",
			7833 => "00000010001111100111101100111001",
			7834 => "0000000110000000001000010000000100",
			7835 => "11111110011000100111101100111001",
			7836 => "00000000000000000111101100111001",
			7837 => "0000000101000000000001000000001000",
			7838 => "0000001010000000000111110100000100",
			7839 => "00000000001100010111101100111001",
			7840 => "00000001101100010111101100111001",
			7841 => "0000001001000000001001111100000100",
			7842 => "00000010110001000111101100111001",
			7843 => "11111110110110000111101100111001",
			7844 => "0000001011000000001011110100011000",
			7845 => "0000000100000000000011010100001100",
			7846 => "0000001010000000001001000100000100",
			7847 => "00000000000000000111101100111001",
			7848 => "0000001001000000001010011000000100",
			7849 => "00000001001100110111101100111001",
			7850 => "00000010000001010111101100111001",
			7851 => "0000000111000000000001111100000100",
			7852 => "00000001111010010111101100111001",
			7853 => "0000000110000000001001111100000100",
			7854 => "11111110001111010111101100111001",
			7855 => "11111111011111110111101100111001",
			7856 => "0000001111000000000010110000001000",
			7857 => "0000001100000000001000011000000100",
			7858 => "11111110000101010111101100111001",
			7859 => "00000000110110100111101100111001",
			7860 => "0000001010000000000001010000000100",
			7861 => "11111110111110000111101100111001",
			7862 => "0000000100000000001011100000000100",
			7863 => "00000001001011000111101100111001",
			7864 => "00000010001101110111101100111001",
			7865 => "0000001001000000001000010100100100",
			7866 => "0000001010000000001010110000100000",
			7867 => "0000001001000000001010100000010000",
			7868 => "0000000111000000000100010000001000",
			7869 => "0000000110000000001000010000000100",
			7870 => "00000001001101010111101100111001",
			7871 => "11111110100101110111101100111001",
			7872 => "0000001010000000000001010000000100",
			7873 => "00000110010001100111101100111001",
			7874 => "00000001001101110111101100111001",
			7875 => "0000001011000000000110100000001000",
			7876 => "0000001100000000001000011000000100",
			7877 => "00000000001011110111101100111001",
			7878 => "11111110011100110111101100111001",
			7879 => "0000000100000000000110001100000100",
			7880 => "00000110010101010111101100111001",
			7881 => "11111110011100010111101100111001",
			7882 => "11111110011000110111101100111001",
			7883 => "0000000000000000000010111100000100",
			7884 => "11111110111111110111101100111001",
			7885 => "00000010001011110111101100111001",
			7886 => "0000000001000000000110101001001100",
			7887 => "0000000100000000000010111000010100",
			7888 => "0000001001000000000101011100010000",
			7889 => "0000001111000000001110000100000100",
			7890 => "00000000000000000111110011111101",
			7891 => "0000000111000000001101100000001000",
			7892 => "0000000111000000001000111000000100",
			7893 => "00000000000000000111110011111101",
			7894 => "11111110101101110111110011111101",
			7895 => "00000000000000000111110011111101",
			7896 => "00000000000000000111110011111101",
			7897 => "0000001100000000000100000000100000",
			7898 => "0000000101000000001010111000010100",
			7899 => "0000000110000000001001100100001100",
			7900 => "0000001100000000000100010100000100",
			7901 => "00000000000000000111110011111101",
			7902 => "0000000100000000000111011100000100",
			7903 => "11111111001111000111110011111101",
			7904 => "00000000000000000111110011111101",
			7905 => "0000001011000000000011011100000100",
			7906 => "00000000000000000111110011111101",
			7907 => "00000000011001000111110011111101",
			7908 => "0000001101000000000100011000000100",
			7909 => "00000000000000000111110011111101",
			7910 => "0000000111000000001001110000000100",
			7911 => "00000001000100000111110011111101",
			7912 => "00000000000000000111110011111101",
			7913 => "0000000100000000000010010000010000",
			7914 => "0000000001000000000110101000001100",
			7915 => "0000001001000000001011101000000100",
			7916 => "00000000000000000111110011111101",
			7917 => "0000000111000000001000111000000100",
			7918 => "00000000000000000111110011111101",
			7919 => "11111110111100000111110011111101",
			7920 => "00000000000000000111110011111101",
			7921 => "0000000110000000001111000000000100",
			7922 => "00000000000000000111110011111101",
			7923 => "00000000010001110111110011111101",
			7924 => "0000000010000000000110111100110100",
			7925 => "0000000110000000001001100100100100",
			7926 => "0000000100000000001100001100100000",
			7927 => "0000000111000000000110100100010000",
			7928 => "0000001100000000001110001100001000",
			7929 => "0000000111000000001101100000000100",
			7930 => "00000000011010010111110011111101",
			7931 => "11111111100110110111110011111101",
			7932 => "0000000001000000000111101000000100",
			7933 => "00000000101101000111110011111101",
			7934 => "00000000000000000111110011111101",
			7935 => "0000001000000000001000100100001000",
			7936 => "0000000001000000000000111100000100",
			7937 => "00000000000000000111110011111101",
			7938 => "00000000001000000111110011111101",
			7939 => "0000000001000000001110010100000100",
			7940 => "11111111011111010111110011111101",
			7941 => "00000000000000000111110011111101",
			7942 => "11111111100100110111110011111101",
			7943 => "0000000100000000001011110000001000",
			7944 => "0000000100000000001111101000000100",
			7945 => "00000000010110010111110011111101",
			7946 => "00000000000000000111110011111101",
			7947 => "0000001010000000000001010000000100",
			7948 => "00000000000000000111110011111101",
			7949 => "00000001010110000111110011111101",
			7950 => "0000001111000000001011110000110100",
			7951 => "0000000010000000000010010100100000",
			7952 => "0000001111000000000000010000010000",
			7953 => "0000000110000000001111000000001000",
			7954 => "0000001100000000001011000000000100",
			7955 => "11111110110011100111110011111101",
			7956 => "00000000000000000111110011111101",
			7957 => "0000001011000000001101111000000100",
			7958 => "00000000110101000111110011111101",
			7959 => "11111111110011110111110011111101",
			7960 => "0000000111000000000110100100001000",
			7961 => "0000001101000000001110000100000100",
			7962 => "00000000010000110111110011111101",
			7963 => "11111111011111100111110011111101",
			7964 => "0000000001000000000101011100000100",
			7965 => "00000000000000000111110011111101",
			7966 => "00000000011101100111110011111101",
			7967 => "0000000110000000000101010000001100",
			7968 => "0000000110000000001111000000000100",
			7969 => "00000000000000000111110011111101",
			7970 => "0000000100000000001000110100000100",
			7971 => "00000000000000000111110011111101",
			7972 => "11111110100110010111110011111101",
			7973 => "0000000111000000000110100100000100",
			7974 => "00000000011010100111110011111101",
			7975 => "00000000000000000111110011111101",
			7976 => "0000001011000000001011110100010000",
			7977 => "0000000001000000000111101000000100",
			7978 => "00000000000000000111110011111101",
			7979 => "0000001111000000000011001100001000",
			7980 => "0000001001000000000010101100000100",
			7981 => "00000001001100000111110011111101",
			7982 => "00000000000000000111110011111101",
			7983 => "00000000000000000111110011111101",
			7984 => "0000000110000000001001111100010000",
			7985 => "0000000111000000000000011100001000",
			7986 => "0000001001000000000011101000000100",
			7987 => "11111111110100110111110011111101",
			7988 => "00000000000000000111110011111101",
			7989 => "0000000001000000001100011000000100",
			7990 => "00000000011111010111110011111101",
			7991 => "00000000000000000111110011111101",
			7992 => "0000000011000000000011011000001000",
			7993 => "0000000111000000000010001000000100",
			7994 => "00000000000000000111110011111101",
			7995 => "11111111000011010111110011111101",
			7996 => "0000000010000000000011111000000100",
			7997 => "00000000000000010111110011111101",
			7998 => "00000000000000000111110011111101",
			7999 => "0000000110000000001101011001000100",
			8000 => "0000001001000000000101010000100000",
			8001 => "0000000001000000000111100100001100",
			8002 => "0000000011000000001010001100000100",
			8003 => "11111110011000110111111011001011",
			8004 => "0000001110000000000110100100000100",
			8005 => "00000000111001010111111011001011",
			8006 => "11111110100000000111111011001011",
			8007 => "0000000111000000000011100000010000",
			8008 => "0000001100000000001110001100000100",
			8009 => "11111110100100100111111011001011",
			8010 => "0000000000000000000001110000000100",
			8011 => "11111110110011100111111011001011",
			8012 => "0000000000000000001101010000000100",
			8013 => "00000010101100100111111011001011",
			8014 => "11111111101001110111111011001011",
			8015 => "11111110010111100111111011001011",
			8016 => "0000001010000000001010100100001000",
			8017 => "0000001001000000000101010000000100",
			8018 => "11111111100001000111111011001011",
			8019 => "00000011101100000111111011001011",
			8020 => "0000000111000000001001001000000100",
			8021 => "11111110100101010111111011001011",
			8022 => "0000001000000000000001010000010000",
			8023 => "0000000001000000001011111100001000",
			8024 => "0000000001000000000001000100000100",
			8025 => "00000000000010110111111011001011",
			8026 => "11111110111001110111111011001011",
			8027 => "0000001000000000000110011000000100",
			8028 => "00000000110001100111111011001011",
			8029 => "00000011011000000111111011001011",
			8030 => "0000001010000000000011101000000100",
			8031 => "11111110110010010111111011001011",
			8032 => "00000000001100110111111011001011",
			8033 => "0000001100000000001000011001110100",
			8034 => "0000000110000000001001100100111000",
			8035 => "0000000010000000001001100000011000",
			8036 => "0000000011000000000100000100001100",
			8037 => "0000000100000000001001001100000100",
			8038 => "11111110010011110111111011001011",
			8039 => "0000000011000000001010111100000100",
			8040 => "11111110101000000111111011001011",
			8041 => "00000010001010110111111011001011",
			8042 => "0000000000000000000011111100001000",
			8043 => "0000000110000000001011001100000100",
			8044 => "00000000010010110111111011001011",
			8045 => "00000001111010010111111011001011",
			8046 => "00000010011110000111111011001011",
			8047 => "0000000011000000001100010000010000",
			8048 => "0000001111000000001110010000001000",
			8049 => "0000001000000000001001101000000100",
			8050 => "11111011100100110111111011001011",
			8051 => "00000000010000110111111011001011",
			8052 => "0000000010000000001100010000000100",
			8053 => "11111111101000000111111011001011",
			8054 => "11111110001000000111111011001011",
			8055 => "0000001111000000001010000100001000",
			8056 => "0000000001000000000001111000000100",
			8057 => "00000011001011010111111011001011",
			8058 => "11111110110000000111111011001011",
			8059 => "0000000000000000001011010100000100",
			8060 => "11111110011000000111111011001011",
			8061 => "00000000100011000111111011001011",
			8062 => "0000001000000000000001110000100000",
			8063 => "0000000111000000001000011000010000",
			8064 => "0000000100000000001000000100001000",
			8065 => "0000000000000000000111000100000100",
			8066 => "11111110100100100111111011001011",
			8067 => "00000001111000010111111011001011",
			8068 => "0000000011000000001100111000000100",
			8069 => "11111101100001010111111011001011",
			8070 => "00000001110000000111111011001011",
			8071 => "0000001101000000000110010000001000",
			8072 => "0000001101000000000100101000000100",
			8073 => "00000000100100110111111011001011",
			8074 => "11111110001011010111111011001011",
			8075 => "0000000111000000000001011000000100",
			8076 => "00000010111101010111111011001011",
			8077 => "11111111010101000111111011001011",
			8078 => "0000001110000000000001011100010000",
			8079 => "0000000111000000001101100000001000",
			8080 => "0000000001000000000110101000000100",
			8081 => "00000001000101010111111011001011",
			8082 => "00000001110010000111111011001011",
			8083 => "0000001000000000001001101000000100",
			8084 => "00000001111001110111111011001011",
			8085 => "00000000000010010111111011001011",
			8086 => "0000001000000000000111000100001000",
			8087 => "0000000110000000001000010000000100",
			8088 => "00000011010010010111111011001011",
			8089 => "00000001101010110111111011001011",
			8090 => "00000000011000110111111011001011",
			8091 => "0000001101000000000110111100010100",
			8092 => "0000000001000000000001111000010000",
			8093 => "0000000001000000000001111000001100",
			8094 => "0000001101000000001100000000000100",
			8095 => "11111110100111000111111011001011",
			8096 => "0000000000000000001101010000000100",
			8097 => "00000001101011100111111011001011",
			8098 => "11111111011010010111111011001011",
			8099 => "00000011001111010111111011001011",
			8100 => "11111110011010100111111011001011",
			8101 => "0000000000000000000111000000001100",
			8102 => "0000000011000000001100001100001000",
			8103 => "0000001100000000000111010000000100",
			8104 => "11111111001110000111111011001011",
			8105 => "00000001111000100111111011001011",
			8106 => "00000111111111010111111011001011",
			8107 => "0000000000000000001011000100001100",
			8108 => "0000000100000000001010110100000100",
			8109 => "11111110011111010111111011001011",
			8110 => "0000001010000000000001010000000100",
			8111 => "00000010100101100111111011001011",
			8112 => "00000000010111110111111011001011",
			8113 => "11111110011001010111111011001011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(2750, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(5367, initial_addr_3'length));
	end generate gen_rom_9;

	gen_rom_10: if SELECT_ROM = 10 generate
		bank <= (
			0 => "00000000000000000000000000000101",
			1 => "00000000000000000000000000001001",
			2 => "00000000000000000000000000001101",
			3 => "00000000000000000000000000010001",
			4 => "00000000000000000000000000010101",
			5 => "00000000000000000000000000011001",
			6 => "00000000000000000000000000011101",
			7 => "00000000000000000000000000100001",
			8 => "00000000000000000000000000100101",
			9 => "00000000000000000000000000101001",
			10 => "00000000000000000000000000101101",
			11 => "00000000000000000000000000110001",
			12 => "00000000000000000000000000110101",
			13 => "00000000000000000000000000111001",
			14 => "00000000000000000000000000111101",
			15 => "00000000000000000000000001000001",
			16 => "00000000000000000000000001000101",
			17 => "00000000000000000000000001001001",
			18 => "00000000000000000000000001001101",
			19 => "00000000000000000000000001010001",
			20 => "0000000100000000001111100100000100",
			21 => "00000000000000000000000001100101",
			22 => "0000000001000000001100011000000100",
			23 => "11111111101111010000000001100101",
			24 => "00000000000000000000000001100101",
			25 => "0000000110000000000100111100000100",
			26 => "00000000000000000000000001111001",
			27 => "0000000110000000001001111100000100",
			28 => "00000000000100010000000001111001",
			29 => "00000000000000000000000001111001",
			30 => "0000000001000000000100110100001000",
			31 => "0000001001000000000111101100000100",
			32 => "00000000000000000000000010001101",
			33 => "00000000010010010000000010001101",
			34 => "00000000000000000000000010001101",
			35 => "0000000001000000001100011000001000",
			36 => "0000000000000000000001110000000100",
			37 => "00000000000000000000000010100001",
			38 => "11111111111010010000000010100001",
			39 => "00000000000000000000000010100001",
			40 => "0000001001000000001010100100001000",
			41 => "0000001110000000001011110000000100",
			42 => "11111111110100100000000010110101",
			43 => "00000000000000000000000010110101",
			44 => "00000000000000000000000010110101",
			45 => "0000000000000000000010101000001100",
			46 => "0000000000000000000010101000000100",
			47 => "00000000000000000000000011010001",
			48 => "0000001000000000000101000100000100",
			49 => "00000000000000000000000011010001",
			50 => "00000000001100000000000011010001",
			51 => "11111111111101100000000011010001",
			52 => "0000001110000000001100001100001100",
			53 => "0000000001000000001100011000001000",
			54 => "0000001110000000001011111000000100",
			55 => "00000000000000000000000011101101",
			56 => "11111111111001100000000011101101",
			57 => "00000000000000000000000011101101",
			58 => "00000000000000000000000011101101",
			59 => "0000000100000000001000011100000100",
			60 => "00000000000000000000000100001001",
			61 => "0000000100000000001011100000001000",
			62 => "0000001001000000000100101100000100",
			63 => "00000000000000000000000100001001",
			64 => "11111111110110110000000100001001",
			65 => "00000000000000000000000100001001",
			66 => "0000001001000000001010100000000100",
			67 => "00000000000000000000000100100101",
			68 => "0000000101000000000111011000001000",
			69 => "0000001001000000000011101000000100",
			70 => "00000000010001010000000100100101",
			71 => "00000000000000000000000100100101",
			72 => "00000000000000000000000100100101",
			73 => "0000000000000000000010101000001100",
			74 => "0000001001000000001010100100000100",
			75 => "00000000000000000000000101010001",
			76 => "0000001111000000000011000000000100",
			77 => "00000000010100110000000101010001",
			78 => "00000000000000000000000101010001",
			79 => "0000001111000000000101000000001000",
			80 => "0000000000000000001010101100000100",
			81 => "00000000000000000000000101010001",
			82 => "11111111110110110000000101010001",
			83 => "00000000000000000000000101010001",
			84 => "0000001011000000001011011100000100",
			85 => "00000000000000000000000101110101",
			86 => "0000000110000000001001111100001100",
			87 => "0000000110000000000100111100000100",
			88 => "00000000000000000000000101110101",
			89 => "0000001011000000000110100000000100",
			90 => "00000000001101000000000101110101",
			91 => "00000000000000000000000101110101",
			92 => "00000000000000000000000101110101",
			93 => "0000000111000000000110100100001000",
			94 => "0000001100000000001101010100000100",
			95 => "00000000000000000000000110100001",
			96 => "00000000000001000000000110100001",
			97 => "0000000001000000000111101000000100",
			98 => "00000000000000000000000110100001",
			99 => "0000001001000000001010100100001000",
			100 => "0000001001000000000100101100000100",
			101 => "00000000000000000000000110100001",
			102 => "11111111100111010000000110100001",
			103 => "00000000000000000000000110100001",
			104 => "0000000111000000000001101000010000",
			105 => "0000000000000000000010101000001100",
			106 => "0000000111000000001000000000000100",
			107 => "00000000000000000000000111001101",
			108 => "0000000000000000000001010100000100",
			109 => "00000000000000000000000111001101",
			110 => "00000000001011110000000111001101",
			111 => "00000000000000000000000111001101",
			112 => "0000000111000000000111010000000100",
			113 => "11111111110000100000000111001101",
			114 => "00000000000000000000000111001101",
			115 => "0000000000000000001010101100001100",
			116 => "0000001001000000001010100100000100",
			117 => "00000000000000000000001000001001",
			118 => "0000000011000000000001011100000100",
			119 => "00000000100010110000001000001001",
			120 => "00000000000000000000001000001001",
			121 => "0000001110000000001110000000001000",
			122 => "0000000001000000001100011000000100",
			123 => "11111111011101000000001000001001",
			124 => "00000000000000000000001000001001",
			125 => "0000001101000000001111100100001000",
			126 => "0000000111000000000111010000000100",
			127 => "00000000000000000000001000001001",
			128 => "00000000010001010000001000001001",
			129 => "00000000000000000000001000001001",
			130 => "0000000100000000001011110000010100",
			131 => "0000000011000000001101101100010000",
			132 => "0000001100000000001000000000001100",
			133 => "0000001100000000001101010100000100",
			134 => "00000000000000000000001000111101",
			135 => "0000000100000000000010000100000100",
			136 => "00000000000000000000001000111101",
			137 => "00000000001101000000001000111101",
			138 => "00000000000000000000001000111101",
			139 => "00000000000000000000001000111101",
			140 => "0000000011000000001000000100000100",
			141 => "11111111111010110000001000111101",
			142 => "00000000000000000000001000111101",
			143 => "0000001011000000001011011100000100",
			144 => "00000000000000000000001001101001",
			145 => "0000000110000000001001111100010000",
			146 => "0000000110000000000100111100000100",
			147 => "00000000000000000000001001101001",
			148 => "0000000101000000000111011000001000",
			149 => "0000000101000000001100100100000100",
			150 => "00000000000000000000001001101001",
			151 => "00000000001111110000001001101001",
			152 => "00000000000000000000001001101001",
			153 => "00000000000000000000001001101001",
			154 => "0000001001000000000111101100010000",
			155 => "0000000111000000000111010000001100",
			156 => "0000001110000000001000101000001000",
			157 => "0000000110000000000100110100000100",
			158 => "00000000000000000000001010101101",
			159 => "11111111110101000000001010101101",
			160 => "00000000000000000000001010101101",
			161 => "00000000000000000000001010101101",
			162 => "0000001001000000000011101000010000",
			163 => "0000000110000000001001111100001100",
			164 => "0000001010000000000011101000000100",
			165 => "00000000000000000000001010101101",
			166 => "0000001110000000000110010000000100",
			167 => "00000000000000000000001010101101",
			168 => "00000000001011110000001010101101",
			169 => "00000000000000000000001010101101",
			170 => "00000000000000000000001010101101",
			171 => "0000000111000000000110100100010100",
			172 => "0000001100000000001101010100000100",
			173 => "00000000000000000000001011110001",
			174 => "0000001000000000000001010100001100",
			175 => "0000001000000000001000010100000100",
			176 => "00000000000000000000001011110001",
			177 => "0000000111000000000011100000000100",
			178 => "00000000000000000000001011110001",
			179 => "00000000000111010000001011110001",
			180 => "00000000000000000000001011110001",
			181 => "0000000001000000000111101000000100",
			182 => "00000000000000000000001011110001",
			183 => "0000001001000000001010100100001000",
			184 => "0000001001000000000100101100000100",
			185 => "00000000000000000000001011110001",
			186 => "11111111100100110000001011110001",
			187 => "00000000000000000000001011110001",
			188 => "0000000100000000001011110000010100",
			189 => "0000001110000000001011101100010000",
			190 => "0000001000000000001010110000000100",
			191 => "00000000000000000000001101000101",
			192 => "0000001110000000000110010000000100",
			193 => "00000000000000000000001101000101",
			194 => "0000000000000000000010101000000100",
			195 => "00000000010100100000001101000101",
			196 => "00000000000000000000001101000101",
			197 => "00000000000000000000001101000101",
			198 => "0000001110000000001110000000001100",
			199 => "0000001001000000001001111100000100",
			200 => "00000000000000000000001101000101",
			201 => "0000001001000000000010101100000100",
			202 => "11111111101110100000001101000101",
			203 => "00000000000000000000001101000101",
			204 => "0000000101000000001111010100001000",
			205 => "0000001011000000001011110100000100",
			206 => "00000000000000000000001101000101",
			207 => "00000000001100000000001101000101",
			208 => "00000000000000000000001101000101",
			209 => "0000000100000000001011110000011000",
			210 => "0000001110000000001011101100010100",
			211 => "0000001101000000001110101100000100",
			212 => "00000000000000000000001110000001",
			213 => "0000001101000000001100010100001100",
			214 => "0000001000000000001000100100000100",
			215 => "00000000000000000000001110000001",
			216 => "0000000000000000001010101100000100",
			217 => "00000000010100010000001110000001",
			218 => "00000000000000000000001110000001",
			219 => "00000000000000000000001110000001",
			220 => "00000000000000000000001110000001",
			221 => "0000001110000000000010010100000100",
			222 => "11111111110100110000001110000001",
			223 => "00000000000000000000001110000001",
			224 => "0000001101000000001111100100011000",
			225 => "0000000110000000001011001100000100",
			226 => "00000000000000000000001110110101",
			227 => "0000000110000000001001111100010000",
			228 => "0000001100000000001101010100000100",
			229 => "00000000000000000000001110110101",
			230 => "0000000000000000000000111000001000",
			231 => "0000001010000000000011101000000100",
			232 => "00000000000000000000001110110101",
			233 => "00000000001100010000001110110101",
			234 => "00000000000000000000001110110101",
			235 => "00000000000000000000001110110101",
			236 => "00000000000000000000001110110101",
			237 => "0000000101000000001001010000000100",
			238 => "00000000000000000000001111101001",
			239 => "0000001101000000001011111000010100",
			240 => "0000001001000000000010101100010000",
			241 => "0000000000000000000010101000000100",
			242 => "00000000000000000000001111101001",
			243 => "0000001110000000001100111000000100",
			244 => "00000000000000000000001111101001",
			245 => "0000000100000000000111011100000100",
			246 => "00000000011011000000001111101001",
			247 => "00000000000000000000001111101001",
			248 => "00000000000000000000001111101001",
			249 => "00000000000000000000001111101001",
			250 => "0000001101000000001110010000011000",
			251 => "0000001001000000000000001000000100",
			252 => "00000000000000000000010000110101",
			253 => "0000001110000000001111101000010000",
			254 => "0000000111000000001000011000001100",
			255 => "0000001010000000001001000100001000",
			256 => "0000001000000000001010110000000100",
			257 => "00000000000000000000010000110101",
			258 => "00000000101101100000010000110101",
			259 => "00000000000000000000010000110101",
			260 => "00000000000000000000010000110101",
			261 => "00000000000000000000010000110101",
			262 => "0000000001000000000111101000000100",
			263 => "00000000000000000000010000110101",
			264 => "0000000010000000000011110100001000",
			265 => "0000001001000000000100101100000100",
			266 => "00000000000000000000010000110101",
			267 => "11111111110000110000010000110101",
			268 => "00000000000000000000010000110101",
			269 => "0000000000000000000001110100010100",
			270 => "0000000011000000001111100100010000",
			271 => "0000000110000000000100110100000100",
			272 => "00000000000000000000010010010001",
			273 => "0000001101000000001110010000001000",
			274 => "0000001100000000001101010100000100",
			275 => "00000000000000000000010010010001",
			276 => "00000000100100100000010010010001",
			277 => "00000000000000000000010010010001",
			278 => "00000000000000000000010010010001",
			279 => "0000000111000000001111011100001100",
			280 => "0000001001000000001010100100001000",
			281 => "0000000001000000001100011000000100",
			282 => "11111111010010110000010010010001",
			283 => "00000000000000000000010010010001",
			284 => "00000000000000000000010010010001",
			285 => "0000000001000000000100110100001100",
			286 => "0000001101000000001111100100001000",
			287 => "0000001001000000001111000000000100",
			288 => "00000000000000000000010010010001",
			289 => "00000000011110100000010010010001",
			290 => "00000000000000000000010010010001",
			291 => "00000000000000000000010010010001",
			292 => "0000001001000000000111101100001100",
			293 => "0000000110000000001000010000001000",
			294 => "0000001100000000001000011000000100",
			295 => "11111111110010110000010011011101",
			296 => "00000000000000000000010011011101",
			297 => "00000000000000000000010011011101",
			298 => "0000001101000000001110010000011000",
			299 => "0000001110000000001111101000010100",
			300 => "0000000101000000001100100100000100",
			301 => "00000000000000000000010011011101",
			302 => "0000000000000000000111000100000100",
			303 => "00000000000000000000010011011101",
			304 => "0000001100000000001001001000001000",
			305 => "0000001000000000000001110000000100",
			306 => "00000000110100110000010011011101",
			307 => "00000000000000000000010011011101",
			308 => "00000000000000000000010011011101",
			309 => "00000000000000000000010011011101",
			310 => "00000000000000000000010011011101",
			311 => "0000000110000000000100111100001100",
			312 => "0000000100000000001011101100000100",
			313 => "00000000000000000000010100101001",
			314 => "0000000001000000001010011000000100",
			315 => "11111111100000110000010100101001",
			316 => "00000000000000000000010100101001",
			317 => "0000001100000000000001011000011000",
			318 => "0000000000000000000010101000000100",
			319 => "00000000000000000000010100101001",
			320 => "0000000000000000000010111100010000",
			321 => "0000001011000000000010001000000100",
			322 => "00000000000000000000010100101001",
			323 => "0000001100000000000100011000000100",
			324 => "00000000000000000000010100101001",
			325 => "0000001101000000000111010100000100",
			326 => "00000000011100100000010100101001",
			327 => "00000000000000000000010100101001",
			328 => "00000000000000000000010100101001",
			329 => "00000000000000000000010100101001",
			330 => "0000000000000000001010101100011100",
			331 => "0000001011000000000101110100011000",
			332 => "0000001001000000000000001000000100",
			333 => "00000000000000000000010101101101",
			334 => "0000000111000000001000011000010000",
			335 => "0000000010000000001000101000001100",
			336 => "0000000101000000001100100100000100",
			337 => "00000000000000000000010101101101",
			338 => "0000000000000000000111000100000100",
			339 => "00000000000000000000010101101101",
			340 => "00000000101011010000010101101101",
			341 => "00000000000000000000010101101101",
			342 => "00000000000000000000010101101101",
			343 => "00000000000000000000010101101101",
			344 => "0000000110000000001000010000000100",
			345 => "11111111110010010000010101101101",
			346 => "00000000000000000000010101101101",
			347 => "0000001001000000000111101100010100",
			348 => "0000000110000000001000010000001000",
			349 => "0000000000000000000111000100000100",
			350 => "00000000000000000000010111011001",
			351 => "11111111001001010000010111011001",
			352 => "0000000100000000000000010100001000",
			353 => "0000000101000000000111111100000100",
			354 => "00000000000000000000010111011001",
			355 => "00000000010011000000010111011001",
			356 => "00000000000000000000010111011001",
			357 => "0000001011000000000001000000100000",
			358 => "0000000001000000000100110100010000",
			359 => "0000001010000000000011101000000100",
			360 => "00000000000000000000010111011001",
			361 => "0000000000000000001011010100000100",
			362 => "00000000000000000000010111011001",
			363 => "0000001110000000000110010000000100",
			364 => "00000000000000000000010111011001",
			365 => "00000000101000110000010111011001",
			366 => "0000000000000000000111000000001000",
			367 => "0000000000000000000001110100000100",
			368 => "00000000000000000000010111011001",
			369 => "11111111101011000000010111011001",
			370 => "0000000000000000000010011000000100",
			371 => "00000000001011110000010111011001",
			372 => "00000000000000000000010111011001",
			373 => "11111111111001110000010111011001",
			374 => "0000000110000000000100111100000100",
			375 => "00000000000000000000011000010101",
			376 => "0000001101000000001111100100011000",
			377 => "0000000110000000001001111100010100",
			378 => "0000001101000000000111111100000100",
			379 => "00000000000000000000011000010101",
			380 => "0000001010000000000110011100001100",
			381 => "0000001011000000000110110100000100",
			382 => "00000000000000000000011000010101",
			383 => "0000001010000000001000010100000100",
			384 => "00000000000000000000011000010101",
			385 => "00000000010001100000011000010101",
			386 => "00000000000000000000011000010101",
			387 => "00000000000000000000011000010101",
			388 => "00000000000000000000011000010101",
			389 => "0000001011000000001011011100001000",
			390 => "0000000100000000001011101100000100",
			391 => "00000000000000000000011001110001",
			392 => "11111111101111100000011001110001",
			393 => "0000001011000000000010110100011000",
			394 => "0000000110000000001001100100000100",
			395 => "00000000000000000000011001110001",
			396 => "0000001000000000001011010100010000",
			397 => "0000001001000000000011101000001100",
			398 => "0000001100000000000100011000000100",
			399 => "00000000000000000000011001110001",
			400 => "0000000111000000000001101000000100",
			401 => "00000000000000000000011001110001",
			402 => "00000000100001100000011001110001",
			403 => "00000000000000000000011001110001",
			404 => "00000000000000000000011001110001",
			405 => "0000001000000000001111001000001100",
			406 => "0000001100000000001111011100000100",
			407 => "00000000000000000000011001110001",
			408 => "0000000111000000000010001000000100",
			409 => "00000000000000000000011001110001",
			410 => "11111111110011010000011001110001",
			411 => "00000000000000000000011001110001",
			412 => "0000000000000000000010101000010100",
			413 => "0000001001000000000000001000000100",
			414 => "00000000000000000000011011010101",
			415 => "0000000111000000001000011000001100",
			416 => "0000000010000000001000101000001000",
			417 => "0000001110000000000110010000000100",
			418 => "00000000000000000000011011010101",
			419 => "00000000110011110000011011010101",
			420 => "00000000000000000000011011010101",
			421 => "00000000000000000000011011010101",
			422 => "0000000111000000001111011100000100",
			423 => "11111111001010010000011011010101",
			424 => "0000000110000000001000010000001000",
			425 => "0000000111000000000101100100000100",
			426 => "00000000000000000000011011010101",
			427 => "11111111110010100000011011010101",
			428 => "0000001101000000001011111000010000",
			429 => "0000001001000000000010101100001100",
			430 => "0000000110000000001001111100001000",
			431 => "0000001110000000001100111000000100",
			432 => "00000000000000000000011011010101",
			433 => "00000000100110110000011011010101",
			434 => "00000000000000000000011011010101",
			435 => "00000000000000000000011011010101",
			436 => "00000000000000000000011011010101",
			437 => "0000001001000000000111101100011100",
			438 => "0000001110000000000001011100001100",
			439 => "0000000100000000001100010000000100",
			440 => "00000000000000000000011101100001",
			441 => "0000001100000000001111011100000100",
			442 => "11111111001111010000011101100001",
			443 => "00000000000000000000011101100001",
			444 => "0000000101000000000010000100001100",
			445 => "0000000111000000000111010000000100",
			446 => "00000000000000000000011101100001",
			447 => "0000000100000000000011010100000100",
			448 => "00000000001011100000011101100001",
			449 => "00000000000000000000011101100001",
			450 => "00000000000000000000011101100001",
			451 => "0000001110000000001011101100010000",
			452 => "0000000101000000001100100100000100",
			453 => "00000000000000000000011101100001",
			454 => "0000000000000000001010101100001000",
			455 => "0000000000000000000111000100000100",
			456 => "00000000000000000000011101100001",
			457 => "00000000101010110000011101100001",
			458 => "00000000000000000000011101100001",
			459 => "0000000000000000000111000000001000",
			460 => "0000001000000000000001010100000100",
			461 => "00000000000000000000011101100001",
			462 => "11111111101001000000011101100001",
			463 => "0000000101000000000110111100010000",
			464 => "0000000110000000001000010000000100",
			465 => "00000000000000000000011101100001",
			466 => "0000000101000000001001010000000100",
			467 => "00000000000000000000011101100001",
			468 => "0000000110000000001001111100000100",
			469 => "00000000100010000000011101100001",
			470 => "00000000000000000000011101100001",
			471 => "00000000000000000000011101100001",
			472 => "0000000100000000001000110100011100",
			473 => "0000001101000000001100010100011000",
			474 => "0000000110000000001000010000010100",
			475 => "0000000000000000000010101000010000",
			476 => "0000000110000000000100110100000100",
			477 => "00000000000000000000011111010101",
			478 => "0000000010000000001000101000001000",
			479 => "0000000111000000000011100000000100",
			480 => "00000000000000000000011111010101",
			481 => "00000000011110100000011111010101",
			482 => "00000000000000000000011111010101",
			483 => "00000000000000000000011111010101",
			484 => "00000000000000000000011111010101",
			485 => "00000000000000000000011111010101",
			486 => "0000000101000000000111111100001000",
			487 => "0000000000000000001010101100000100",
			488 => "00000000000000000000011111010101",
			489 => "11111111001101100000011111010101",
			490 => "0000000111000000000100010000010000",
			491 => "0000000100000000001110111000001100",
			492 => "0000001010000000001000010100000100",
			493 => "00000000000000000000011111010101",
			494 => "0000001001000000000010101100000100",
			495 => "00000000101100110000011111010101",
			496 => "00000000000000000000011111010101",
			497 => "00000000000000000000011111010101",
			498 => "0000001110000000001110100100000100",
			499 => "11111111101111100000011111010101",
			500 => "00000000000000000000011111010101",
			501 => "0000000000000000001101010000101100",
			502 => "0000001100000000000100011000010000",
			503 => "0000000100000000001000100000001100",
			504 => "0000001010000000000011101000000100",
			505 => "00000000000000000000100001011001",
			506 => "0000001110000000000110010000000100",
			507 => "00000000000000000000100001011001",
			508 => "00000000000111000000100001011001",
			509 => "11111111110001000000100001011001",
			510 => "0000000111000000000101100100010100",
			511 => "0000001001000000000011101000010000",
			512 => "0000001101000000000101110000000100",
			513 => "00000000000000000000100001011001",
			514 => "0000001000000000001100000100001000",
			515 => "0000001010000000001000100100000100",
			516 => "00000000000000000000100001011001",
			517 => "00000000101010100000100001011001",
			518 => "00000000000000000000100001011001",
			519 => "00000000000000000000100001011001",
			520 => "0000001000000000000001110000000100",
			521 => "11111111111110010000100001011001",
			522 => "00000000000000000000100001011001",
			523 => "0000001110000000001100001100000100",
			524 => "11111111001011000000100001011001",
			525 => "0000001001000000001010100100010000",
			526 => "0000001101000000001011111000001100",
			527 => "0000000011000000000101000000000100",
			528 => "00000000000000000000100001011001",
			529 => "0000000000000000001000111100000100",
			530 => "00000000100101000000100001011001",
			531 => "00000000000000000000100001011001",
			532 => "00000000000000000000100001011001",
			533 => "00000000000000000000100001011001",
			534 => "0000000100000000001000110100011100",
			535 => "0000001101000000001100010100011000",
			536 => "0000000110000000001000010000010100",
			537 => "0000000110000000000100110100000100",
			538 => "00000000000000000000100011010101",
			539 => "0000000010000000001000101000001100",
			540 => "0000001010000000001000010100001000",
			541 => "0000000111000000000011100000000100",
			542 => "00000000000000000000100011010101",
			543 => "00000000011011100000100011010101",
			544 => "00000000000000000000100011010101",
			545 => "00000000000000000000100011010101",
			546 => "00000000000000000000100011010101",
			547 => "00000000000000000000100011010101",
			548 => "0000001110000000001000110100001100",
			549 => "0000000001000000001110010100000100",
			550 => "00000000000000000000100011010101",
			551 => "0000001001000000001001111100000100",
			552 => "00000000000000000000100011010101",
			553 => "11111111011001100000100011010101",
			554 => "0000001101000000001111100100010100",
			555 => "0000000111000000000111010000000100",
			556 => "00000000000000000000100011010101",
			557 => "0000000001000000000001000100000100",
			558 => "00000000000000000000100011010101",
			559 => "0000000001000000001100011000001000",
			560 => "0000001110000000001000011100000100",
			561 => "00000000000000000000100011010101",
			562 => "00000000101100000000100011010101",
			563 => "00000000000000000000100011010101",
			564 => "00000000000000000000100011010101",
			565 => "0000000111000000001000011000100100",
			566 => "0000001100000000000100011000001100",
			567 => "0000000100000000001000100000000100",
			568 => "00000000000000000000100101100001",
			569 => "0000000001000000001100011000000100",
			570 => "11111111110001010000100101100001",
			571 => "00000000000000000000100101100001",
			572 => "0000001100000000001000000000010100",
			573 => "0000001101000000001110010000010000",
			574 => "0000001010000000001001000100001100",
			575 => "0000000111000000000110100100000100",
			576 => "00000000000000000000100101100001",
			577 => "0000000110000000000100110100000100",
			578 => "00000000000000000000100101100001",
			579 => "00000000101101000000100101100001",
			580 => "00000000000000000000100101100001",
			581 => "00000000000000000000100101100001",
			582 => "00000000000000000000100101100001",
			583 => "0000000111000000001111011100000100",
			584 => "11111111010011000000100101100001",
			585 => "0000000101000000000110111100011000",
			586 => "0000000001000000000100110100010000",
			587 => "0000000001000000000101011100000100",
			588 => "00000000000000000000100101100001",
			589 => "0000001100000000001001110100000100",
			590 => "00000000000000000000100101100001",
			591 => "0000000101000000000101110000000100",
			592 => "00000000000000000000100101100001",
			593 => "00000000100100110000100101100001",
			594 => "0000000111000000001111011100000100",
			595 => "00000000000000000000100101100001",
			596 => "11111111110000010000100101100001",
			597 => "0000001100000000000100000100000100",
			598 => "00000000000000000000100101100001",
			599 => "11111111101001000000100101100001",
			600 => "0000001001000000001010100000101000",
			601 => "0000000111000000001111011100001000",
			602 => "0000000100000000000110101100000100",
			603 => "00000000000000000000101000001101",
			604 => "11111110110010100000101000001101",
			605 => "0000000111000000000010001000010100",
			606 => "0000000100000000000011001100010000",
			607 => "0000001111000000000000010000000100",
			608 => "00000000000000000000101000001101",
			609 => "0000000000000000000110001000000100",
			610 => "00000000000000000000101000001101",
			611 => "0000000101000000001100010100000100",
			612 => "00000000100111100000101000001101",
			613 => "00000000000000000000101000001101",
			614 => "00000000000000000000101000001101",
			615 => "0000001111000000001000001000001000",
			616 => "0000001100000000001111011100000100",
			617 => "00000000000000000000101000001101",
			618 => "11111111100110010000101000001101",
			619 => "00000000000000000000101000001101",
			620 => "0000001100000000001001110100011100",
			621 => "0000000000000000001000101100011000",
			622 => "0000000101000000001100100100001000",
			623 => "0000001100000000001010111000000100",
			624 => "00000000001011010000101000001101",
			625 => "00000000000000000000101000001101",
			626 => "0000001100000000000100011000000100",
			627 => "00000000000000000000101000001101",
			628 => "0000000001000000001101111100000100",
			629 => "00000000000000000000101000001101",
			630 => "0000001001000000001010100000000100",
			631 => "00000000000000000000101000001101",
			632 => "00000001001011000000101000001101",
			633 => "00000000000000000000101000001101",
			634 => "0000000001000000000100110100001100",
			635 => "0000000110000000001000010000000100",
			636 => "00000000000000000000101000001101",
			637 => "0000000101000000000111111100000100",
			638 => "00000000000000000000101000001101",
			639 => "00000000100010100000101000001101",
			640 => "0000000100000000000110111000000100",
			641 => "00000000000000000000101000001101",
			642 => "11111111010100100000101000001101",
			643 => "0000000100000000001000000100100100",
			644 => "0000001001000000001010100100011000",
			645 => "0000000110000000001001100100010100",
			646 => "0000000110000000000100110100000100",
			647 => "00000000000000000000101010110001",
			648 => "0000000001000000001101111100001100",
			649 => "0000000101000000000101110000001000",
			650 => "0000000111000000001000000000000100",
			651 => "00000000000000000000101010110001",
			652 => "00000000101110100000101010110001",
			653 => "00000000000000000000101010110001",
			654 => "00000000000000000000101010110001",
			655 => "11111111100000110000101010110001",
			656 => "0000000111000000001111011100001000",
			657 => "0000000010000000001000101000000100",
			658 => "00000001001110100000101010110001",
			659 => "00000000000000000000101010110001",
			660 => "00000000000000000000101010110001",
			661 => "0000001110000000001100001100011100",
			662 => "0000000100000000001010110100011000",
			663 => "0000000101000000000111111100001000",
			664 => "0000000001000000001100011000000100",
			665 => "11111111011110000000101010110001",
			666 => "00000000000000000000101010110001",
			667 => "0000000100000000000110001100000100",
			668 => "00000000000000000000101010110001",
			669 => "0000001101000000000111011000001000",
			670 => "0000000001000000001100011000000100",
			671 => "00000000101101100000101010110001",
			672 => "00000000000000000000101010110001",
			673 => "00000000000000000000101010110001",
			674 => "11111110111110110000101010110001",
			675 => "0000001011000000000001000000010000",
			676 => "0000001011000000000000110100000100",
			677 => "00000000000000000000101010110001",
			678 => "0000001001000000000010101100001000",
			679 => "0000000001000000001011111100000100",
			680 => "00000000000000000000101010110001",
			681 => "00000001001111010000101010110001",
			682 => "00000000000000000000101010110001",
			683 => "11111111101110100000101010110001",
			684 => "0000000001000000000101011100011000",
			685 => "0000000000000000000111000100010000",
			686 => "0000001010000000000011101000001100",
			687 => "0000001001000000001011111100001000",
			688 => "0000000101000000001111011100000100",
			689 => "11111110100000110000101101010101",
			690 => "00000110010100100000101101010101",
			691 => "11111110011010010000101101010101",
			692 => "00000110110000110000101101010101",
			693 => "0000000001000000001001011000000100",
			694 => "11111110011001000000101101010101",
			695 => "11111101101000110000101101010101",
			696 => "0000001001000000000010101100110100",
			697 => "0000000101000000001001010000011100",
			698 => "0000001001000000001010100000001100",
			699 => "0000000100000000001111100100001000",
			700 => "0000000110000000001011001100000100",
			701 => "11111110100010100000101101010101",
			702 => "00000110011011000000101101010101",
			703 => "11111110010001110000101101010101",
			704 => "0000000010000000001111100100000100",
			705 => "00000100000101010000101101010101",
			706 => "0000000001000000001100011000001000",
			707 => "0000000001000000001100011000000100",
			708 => "11111110010011000000101101010101",
			709 => "00000000001110000000101101010101",
			710 => "00000110000000010000101101010101",
			711 => "0000001000000000000101000100001000",
			712 => "0000001001000000000101010000000100",
			713 => "00000000111100000000101101010101",
			714 => "11111110011011100000101101010101",
			715 => "0000000010000000000010010100000100",
			716 => "00000110010001100000101101010101",
			717 => "0000000101000000000111011000001000",
			718 => "0000000110000000000100111100000100",
			719 => "11111101110000110000101101010101",
			720 => "00000001101101000000101101010101",
			721 => "11111110101010100000101101010101",
			722 => "0000000111000000000001101000000100",
			723 => "00000000011101100000101101010101",
			724 => "11111110011001110000101101010101",
			725 => "0000000000000000000010111101000100",
			726 => "0000001110000000001000110100110100",
			727 => "0000000000000000001000101100101000",
			728 => "0000001011000000001011110100011000",
			729 => "0000000101000000001001010000001100",
			730 => "0000000011000000001111100100001000",
			731 => "0000001001000000000000001000000100",
			732 => "00000000000000000000101111101001",
			733 => "00000000011101010000101111101001",
			734 => "11111111011000110000101111101001",
			735 => "0000000111000000001000011000000100",
			736 => "00000000000000000000101111101001",
			737 => "0000000100000000001111101000000100",
			738 => "00000000000000000000101111101001",
			739 => "00000001001011100000101111101001",
			740 => "0000000000000000000111000000001000",
			741 => "0000000011000000001111101000000100",
			742 => "00000000000000000000101111101001",
			743 => "11111111001001010000101111101001",
			744 => "0000001101000000001110110100000100",
			745 => "00000000011000000000101111101001",
			746 => "00000000000000000000101111101001",
			747 => "0000001110000000001110000000001000",
			748 => "0000001001000000001010100100000100",
			749 => "11111111000000000000101111101001",
			750 => "00000000000000000000101111101001",
			751 => "00000000000000000000101111101001",
			752 => "0000000101000000000111111100000100",
			753 => "00000000000000000000101111101001",
			754 => "0000001010000000000110011000000100",
			755 => "00000000000000000000101111101001",
			756 => "0000000001000000001010011000000100",
			757 => "00000001000111110000101111101001",
			758 => "00000000000000000000101111101001",
			759 => "0000001110000000000010110000000100",
			760 => "11111110111010000000101111101001",
			761 => "00000000000000000000101111101001",
			762 => "0000001100000000001101010100000100",
			763 => "11111110011101110000110001101101",
			764 => "0000000010000000001000100000100000",
			765 => "0000000110000000001011001100001100",
			766 => "0000000001000000001011101000001000",
			767 => "0000000111000000001001001000000100",
			768 => "00000000000000000000110001101101",
			769 => "00000001000111000000110001101101",
			770 => "11111110111100100000110001101101",
			771 => "0000001000000000000101000100010000",
			772 => "0000001110000000001011111000001100",
			773 => "0000001110000000000110010000000100",
			774 => "00000000000000000000110001101101",
			775 => "0000001010000000000011101000000100",
			776 => "00000000000000000000110001101101",
			777 => "00000001010001110000110001101101",
			778 => "00000000000000000000110001101101",
			779 => "11111111101001010000110001101101",
			780 => "0000001011000000000010001000000100",
			781 => "11111110100000010000110001101101",
			782 => "0000001100000000001000000000001100",
			783 => "0000001100000000001011000000000100",
			784 => "00000000000000000000110001101101",
			785 => "0000000001000000000100110100000100",
			786 => "00000000000000000000110001101101",
			787 => "00000001100011000000110001101101",
			788 => "0000001001000000001010100100001100",
			789 => "0000000111000000001111011100000100",
			790 => "11111110100000010000110001101101",
			791 => "0000001101000000001111100100000100",
			792 => "00000000010111100000110001101101",
			793 => "11111110111000010000110001101101",
			794 => "11111110011011000000110001101101",
			795 => "0000000101000000001001010100000100",
			796 => "11111110011010100000110011001001",
			797 => "0000001101000000001111100100101000",
			798 => "0000001001000000000010101100100000",
			799 => "0000000110000000000100110100000100",
			800 => "11111110101011110000110011001001",
			801 => "0000001110000000001100001100010000",
			802 => "0000000000000000001101010000001000",
			803 => "0000000110000000001000010000000100",
			804 => "00000000011000010000110011001001",
			805 => "00000001100011000000110011001001",
			806 => "0000001110000000001000011100000100",
			807 => "11111110001011000000110011001001",
			808 => "00000000000000000000110011001001",
			809 => "0000000000000000000000110000001000",
			810 => "0000000101000000000011001000000100",
			811 => "11111111111010010000110011001001",
			812 => "00000001101110110000110011001001",
			813 => "11111111101011110000110011001001",
			814 => "0000000101000000001110000100000100",
			815 => "00000000100101000000110011001001",
			816 => "11111110100101000000110011001001",
			817 => "11111110001111110000110011001001",
			818 => "0000000101000000000110111100111100",
			819 => "0000000011000000000011110000110000",
			820 => "0000001000000000001100000100101000",
			821 => "0000000110000000001000010000011100",
			822 => "0000001110000000001011111000001100",
			823 => "0000000011000000000000010000000100",
			824 => "00000000000000000000110101000101",
			825 => "0000000110000000001111000000000100",
			826 => "00000000101000110000110101000101",
			827 => "00000000000000000000110101000101",
			828 => "0000000110000000000100111100001000",
			829 => "0000000001000000000001000100000100",
			830 => "00000000000000000000110101000101",
			831 => "11111111001100100000110101000101",
			832 => "0000001111000000001000000100000100",
			833 => "00000000000000000000110101000101",
			834 => "11111111111110010000110101000101",
			835 => "0000000111000000001000011000000100",
			836 => "00000000000000000000110101000101",
			837 => "0000001001000000000010101100000100",
			838 => "00000000101010110000110101000101",
			839 => "00000000000000000000110101000101",
			840 => "0000001110000000001000110100000100",
			841 => "11111111011001110000110101000101",
			842 => "00000000000000000000110101000101",
			843 => "0000001001000000000010101100001000",
			844 => "0000000100000000000001100100000100",
			845 => "00000000110100010000110101000101",
			846 => "00000000000000000000110101000101",
			847 => "00000000000000000000110101000101",
			848 => "11111111100010110000110101000101",
			849 => "0000000111000000000110100100001100",
			850 => "0000001001000000001010100100000100",
			851 => "11111110011001010000110111001001",
			852 => "0000000001000000001100011000000100",
			853 => "00000010001110010000110111001001",
			854 => "00000000000000000000110111001001",
			855 => "0000001101000000001111100100110100",
			856 => "0000001001000000000010101100101100",
			857 => "0000001101000000001001011100010000",
			858 => "0000001101000000000110100000000100",
			859 => "00000010101111100000110111001001",
			860 => "0000001001000000001010100000000100",
			861 => "11111110011100010000110111001001",
			862 => "0000000110000000000100111100000100",
			863 => "00000001110110000000110111001001",
			864 => "11111110101100000000110111001001",
			865 => "0000000010000000001110000000010000",
			866 => "0000001011000000001010010100001000",
			867 => "0000000000000000000110001000000100",
			868 => "11111110111010010000110111001001",
			869 => "00000011010110100000110111001001",
			870 => "0000000001000000001011111100000100",
			871 => "00000001000001100000110111001001",
			872 => "11111110100111110000110111001001",
			873 => "0000001011000000001011110100000100",
			874 => "11111101111101110000110111001001",
			875 => "0000000110000000001000010000000100",
			876 => "11111110111110000000110111001001",
			877 => "00000001010101100000110111001001",
			878 => "0000001011000000000110110100000100",
			879 => "00000001010010000000110111001001",
			880 => "11111110011101000000110111001001",
			881 => "11111110001110000000110111001001",
			882 => "0000001001000000001010100001000000",
			883 => "0000000111000000001111011100011000",
			884 => "0000000000000000000110001000010100",
			885 => "0000001011000000000100000100010000",
			886 => "0000000111000000001000000000000100",
			887 => "00000000000000000000111010100101",
			888 => "0000001100000000001101010100000100",
			889 => "00000000000000000000111010100101",
			890 => "0000000111000000000110100100000100",
			891 => "00000001001010100000111010100101",
			892 => "00000000000000000000111010100101",
			893 => "11111111011110100000111010100101",
			894 => "11111110011101010000111010100101",
			895 => "0000000101000000001110110100011000",
			896 => "0000000011000000001110000000010000",
			897 => "0000001111000000001000110100001100",
			898 => "0000000110000000001001100100000100",
			899 => "11111111110110100000111010100101",
			900 => "0000000111000000000101100100000100",
			901 => "00000000110010110000111010100101",
			902 => "00000000000000000000111010100101",
			903 => "11111111000101110000111010100101",
			904 => "0000000000000000000000110000000100",
			905 => "00000001001000000000111010100101",
			906 => "00000000000000000000111010100101",
			907 => "0000001010000000000001010000000100",
			908 => "11111110101111100000111010100101",
			909 => "0000001101000000001000001100001000",
			910 => "0000001111000000001111100000000100",
			911 => "00000000010100100000111010100101",
			912 => "00000000000000000000111010100101",
			913 => "00000000000000000000111010100101",
			914 => "0000000011000000001101101100010000",
			915 => "0000000000000000001010101100001100",
			916 => "0000001011000000001011011100001000",
			917 => "0000001011000000000000011100000100",
			918 => "00000000101111000000111010100101",
			919 => "00000000000000000000111010100101",
			920 => "00000001110001010000111010100101",
			921 => "00000000000000000000111010100101",
			922 => "0000000000000000000010101000000100",
			923 => "11111111000111000000111010100101",
			924 => "0000000000000000001101010000010100",
			925 => "0000001001000000000010101100001100",
			926 => "0000001101000000001010001000000100",
			927 => "00000000000000000000111010100101",
			928 => "0000000111000000001011011100000100",
			929 => "00000001011100010000111010100101",
			930 => "00000000000000000000111010100101",
			931 => "0000001100000000001000000000000100",
			932 => "00000000000010100000111010100101",
			933 => "11111111000111100000111010100101",
			934 => "0000001110000000000011110000000100",
			935 => "11111111000110000000111010100101",
			936 => "00000000000000000000111010100101",
			937 => "0000000000000000000010101000101100",
			938 => "0000001010000000001000100100100000",
			939 => "0000001110000000001011111000011000",
			940 => "0000000110000000001011001100001000",
			941 => "0000001001000000000000001000000100",
			942 => "11111111110001110000111101110001",
			943 => "00000000000000000000111101110001",
			944 => "0000001000000000000101000100001100",
			945 => "0000001000000000001100011100000100",
			946 => "00000000000000000000111101110001",
			947 => "0000000011000000000111011000000100",
			948 => "00000000000000000000111101110001",
			949 => "00000001000100000000111101110001",
			950 => "00000000000000000000111101110001",
			951 => "0000000000000000000010101000000100",
			952 => "11111111010001010000111101110001",
			953 => "00000000000000000000111101110001",
			954 => "0000000110000000001000010000001000",
			955 => "0000000011000000000001011100000100",
			956 => "00000001011010100000111101110001",
			957 => "00000000000000000000111101110001",
			958 => "00000000000000000000111101110001",
			959 => "0000001110000000000001011100000100",
			960 => "11111110101001010000111101110001",
			961 => "0000001011000000000110100000100100",
			962 => "0000001101000000001100010100010100",
			963 => "0000000110000000001000010000001100",
			964 => "0000001100000000001011000000000100",
			965 => "00000000000000000000111101110001",
			966 => "0000001011000000000100010000000100",
			967 => "00000000000000000000111101110001",
			968 => "00000000011001000000111101110001",
			969 => "0000000111000000001000011000000100",
			970 => "00000000000000000000111101110001",
			971 => "11111111000110100000111101110001",
			972 => "0000001001000000000010101100001100",
			973 => "0000000110000000001000010000000100",
			974 => "00000000000000000000111101110001",
			975 => "0000001000000000000110001000000100",
			976 => "00000001000110010000111101110001",
			977 => "00000000000000000000111101110001",
			978 => "00000000000000000000111101110001",
			979 => "0000000110000000001001111100001000",
			980 => "0000001101000000001111010100000100",
			981 => "00000000000000000000111101110001",
			982 => "11111111001100100000111101110001",
			983 => "0000001001000000001010100100001000",
			984 => "0000001001000000000100101100000100",
			985 => "00000000000000000000111101110001",
			986 => "00000000000111000000111101110001",
			987 => "00000000000000000000111101110001",
			988 => "0000000000000000000010011001001000",
			989 => "0000000011000000001000110100110100",
			990 => "0000000000000000001000110000101100",
			991 => "0000001011000000001011110100011000",
			992 => "0000000101000000001001010000001100",
			993 => "0000000011000000001111100100001000",
			994 => "0000001001000000000000001000000100",
			995 => "11111111111100110001000000001101",
			996 => "00000000011110110001000000001101",
			997 => "11111111001010110001000000001101",
			998 => "0000000111000000001000011000000100",
			999 => "00000000000000000001000000001101",
			1000 => "0000000100000000001111101000000100",
			1001 => "00000000000000000001000000001101",
			1002 => "00000001001111000001000000001101",
			1003 => "0000000000000000000111000000001100",
			1004 => "0000000011000000001111101000000100",
			1005 => "00000000000000000001000000001101",
			1006 => "0000000100000000001100001100000100",
			1007 => "11111111000001010001000000001101",
			1008 => "00000000000000000001000000001101",
			1009 => "0000000101000000000011001000000100",
			1010 => "00000000100011000001000000001101",
			1011 => "00000000000000000001000000001101",
			1012 => "0000000011000000001110000000000100",
			1013 => "11111110111101100001000000001101",
			1014 => "00000000000000000001000000001101",
			1015 => "0000001010000000000110011000000100",
			1016 => "00000000000000000001000000001101",
			1017 => "0000000001000000001100011000001100",
			1018 => "0000000100000000000100001100001000",
			1019 => "0000000000000000000010011000000100",
			1020 => "00000001000111110001000000001101",
			1021 => "00000000000000000001000000001101",
			1022 => "00000000000000000001000000001101",
			1023 => "00000000000000000001000000001101",
			1024 => "0000001110000000000011110000000100",
			1025 => "11111110110011010001000000001101",
			1026 => "00000000000000000001000000001101",
			1027 => "0000000100000000001011110000101100",
			1028 => "0000000110000000001011001100001000",
			1029 => "0000000001000000001101111100000100",
			1030 => "11111111011110000001000011011001",
			1031 => "00000000000000000001000011011001",
			1032 => "0000001110000000001011101100011100",
			1033 => "0000000101000000001100100100010000",
			1034 => "0000000010000000000110111100001000",
			1035 => "0000000011000000000010000100000100",
			1036 => "00000000000000000001000011011001",
			1037 => "00000000000000110001000011011001",
			1038 => "0000001100000000000111001000000100",
			1039 => "00000000000000000001000011011001",
			1040 => "11111111111001010001000011011001",
			1041 => "0000001010000000000011101000000100",
			1042 => "00000000000000000001000011011001",
			1043 => "0000000000000000000110001000000100",
			1044 => "00000000000000000001000011011001",
			1045 => "00000001100001000001000011011001",
			1046 => "0000001100000000001000000000000100",
			1047 => "11111111110101010001000011011001",
			1048 => "00000000000000000001000011011001",
			1049 => "0000001110000000000001011100001000",
			1050 => "0000001001000000000010101100000100",
			1051 => "11111110100111000001000011011001",
			1052 => "00000000000000000001000011011001",
			1053 => "0000000000000000000111000000001000",
			1054 => "0000001110000000001000101000000100",
			1055 => "00000000000000000001000011011001",
			1056 => "11111111001011000001000011011001",
			1057 => "0000001011000000000110100000010100",
			1058 => "0000001011000000001011110100001000",
			1059 => "0000001010000000001001000100000100",
			1060 => "00000000001001100001000011011001",
			1061 => "11111111010001100001000011011001",
			1062 => "0000000100000000001110111000001000",
			1063 => "0000000110000000001000010000000100",
			1064 => "00000000000000000001000011011001",
			1065 => "00000001001100100001000011011001",
			1066 => "00000000000000000001000011011001",
			1067 => "0000000110000000001001111100001100",
			1068 => "0000001101000000001111010100000100",
			1069 => "00000000000000000001000011011001",
			1070 => "0000000100000000001010110100000100",
			1071 => "00000000000000000001000011011001",
			1072 => "11111111001100000001000011011001",
			1073 => "0000000001000000000100110100001000",
			1074 => "0000000001000000001110010100000100",
			1075 => "00000000000000000001000011011001",
			1076 => "00000000001011000001000011011001",
			1077 => "00000000000000000001000011011001",
			1078 => "0000000001000000000101011100011000",
			1079 => "0000000000000000000111000000010000",
			1080 => "0000000011000000001000100000001100",
			1081 => "0000001100000000001011000000000100",
			1082 => "11111110011010000001000110011101",
			1083 => "0000001001000000001101011000000100",
			1084 => "00000110100001000001000110011101",
			1085 => "11111110011101010001000110011101",
			1086 => "00000101011001000001000110011101",
			1087 => "0000001001000000001001100100000100",
			1088 => "11111110011000110001000110011101",
			1089 => "11111100111111100001000110011101",
			1090 => "0000001001000000000010101101000100",
			1091 => "0000000101000000001001010000100000",
			1092 => "0000000100000000000110111000011000",
			1093 => "0000001001000000001010100000001100",
			1094 => "0000001001000000000000001000000100",
			1095 => "11111110011100010001000110011101",
			1096 => "0000000001000000000001111000000100",
			1097 => "00000111101101100001000110011101",
			1098 => "11111111100010100001000110011101",
			1099 => "0000001110000000001000001100000100",
			1100 => "00000110010000000001000110011101",
			1101 => "0000000011000000001011101100000100",
			1102 => "00000001011101110001000110011101",
			1103 => "11111101111010110001000110011101",
			1104 => "0000000001000000001100011000000100",
			1105 => "11111110010011000001000110011101",
			1106 => "00000000011001110001000110011101",
			1107 => "0000001000000000000001010100010000",
			1108 => "0000001001000000000101010000001000",
			1109 => "0000001011000000001011110100000100",
			1110 => "11111111110100000001000110011101",
			1111 => "00000001000100110001000110011101",
			1112 => "0000000111000000000101110100000100",
			1113 => "11111110011100010001000110011101",
			1114 => "11111100110011000001000110011101",
			1115 => "0000000101000000000111011000010000",
			1116 => "0000000100000000000110001100001000",
			1117 => "0000001100000000001001110100000100",
			1118 => "00000110111001100001000110011101",
			1119 => "00000001011100100001000110011101",
			1120 => "0000001110000000001011110000000100",
			1121 => "00000000001010000001000110011101",
			1122 => "00000001111011000001000110011101",
			1123 => "11111110001010000001000110011101",
			1124 => "0000000100000000001011110000000100",
			1125 => "00000001001111010001000110011101",
			1126 => "11111110011001100001000110011101",
			1127 => "0000001011000000001010011100000100",
			1128 => "11111110011010010001001000000001",
			1129 => "0000000101000000001111010100101100",
			1130 => "0000001001000000000010101100100100",
			1131 => "0000000110000000000100110100000100",
			1132 => "11111110101000010001001000000001",
			1133 => "0000000000000000001101010000010000",
			1134 => "0000000110000000001000010000001000",
			1135 => "0000001111000000001011110000000100",
			1136 => "00000000110101010001001000000001",
			1137 => "11111110011101010001001000000001",
			1138 => "0000000111000000001000011000000100",
			1139 => "11111111010100100001001000000001",
			1140 => "00000010000000010001001000000001",
			1141 => "0000001110000000001110100100001000",
			1142 => "0000001110000000001000011100000100",
			1143 => "11111101111111100001001000000001",
			1144 => "00000000000000000001001000000001",
			1145 => "0000000101000000000011001000000100",
			1146 => "11111110111010100001001000000001",
			1147 => "00000001100011100001001000000001",
			1148 => "0000001011000000000110110100000100",
			1149 => "00000000100101010001001000000001",
			1150 => "11111110100001110001001000000001",
			1151 => "11111110001001010001001000000001",
			1152 => "0000001001000000000111101100110000",
			1153 => "0000001100000000001000000000001000",
			1154 => "0000001111000000001000000100000100",
			1155 => "11111110100100110001001011100101",
			1156 => "00000000000000000001001011100101",
			1157 => "0000001101000000001010000100100000",
			1158 => "0000000001000000000101011100010000",
			1159 => "0000001100000000000110100100001000",
			1160 => "0000000001000000001101011100000100",
			1161 => "00000000010111100001001011100101",
			1162 => "00000000000000000001001011100101",
			1163 => "0000001110000000000010010100000100",
			1164 => "11111111011000000001001011100101",
			1165 => "00000000000000000001001011100101",
			1166 => "0000000000000000000010101000000100",
			1167 => "00000000000000000001001011100101",
			1168 => "0000000100000000000011010100001000",
			1169 => "0000001010000000001010110000000100",
			1170 => "00000001000001000001001011100101",
			1171 => "00000000000000000001001011100101",
			1172 => "00000000000000000001001011100101",
			1173 => "0000001110000000000101000000000100",
			1174 => "11111111000111010001001011100101",
			1175 => "00000000000000000001001011100101",
			1176 => "0000000011000000001000100000011100",
			1177 => "0000000101000000001100100100010100",
			1178 => "0000000100000000001011101100001100",
			1179 => "0000001001000000000000001000000100",
			1180 => "00000000000000000001001011100101",
			1181 => "0000001110000000001110110100000100",
			1182 => "00000000000000000001001011100101",
			1183 => "00000000111110000001001011100101",
			1184 => "0000001100000000001010111000000100",
			1185 => "00000000000000000001001011100101",
			1186 => "11111111100100010001001011100101",
			1187 => "0000000000000000000111000100000100",
			1188 => "00000000000000000001001011100101",
			1189 => "00000001101010100001001011100101",
			1190 => "0000001000000000000001010100000100",
			1191 => "11111111000010000001001011100101",
			1192 => "0000001000000000000001110000010000",
			1193 => "0000001001000000000010101100001100",
			1194 => "0000000101000000000001000000000100",
			1195 => "00000000000000000001001011100101",
			1196 => "0000000101000000000111111100000100",
			1197 => "00000001010011010001001011100101",
			1198 => "00000000000000000001001011100101",
			1199 => "00000000000000000001001011100101",
			1200 => "0000001101000000001100010100000100",
			1201 => "11111110111001000001001011100101",
			1202 => "0000000100000000001110111000001000",
			1203 => "0000001100000000001000011000000100",
			1204 => "00000001010001010001001011100101",
			1205 => "00000000000000000001001011100101",
			1206 => "0000001110000000000011110000000100",
			1207 => "11111111101111010001001011100101",
			1208 => "00000000000000000001001011100101",
			1209 => "0000000001000000001101111101000000",
			1210 => "0000001100000000000100011000001000",
			1211 => "0000000011000000000010010100000100",
			1212 => "11111110011100110001001111011001",
			1213 => "00000000000000000001001111011001",
			1214 => "0000000100000000000101000000010100",
			1215 => "0000000110000000001001100100001100",
			1216 => "0000000010000000001010001000001000",
			1217 => "0000000100000000000010000000000100",
			1218 => "00000000000000000001001111011001",
			1219 => "00000000001010100001001111011001",
			1220 => "11111110111101110001001111011001",
			1221 => "0000001011000000000110110100000100",
			1222 => "00000000000000000001001111011001",
			1223 => "00000001010110000001001111011001",
			1224 => "0000001110000000001000011100010000",
			1225 => "0000001001000000001001111100001100",
			1226 => "0000001001000000001000010000000100",
			1227 => "11111111000100000001001111011001",
			1228 => "0000000000000000001000101100000100",
			1229 => "00000000000110010001001111011001",
			1230 => "00000000000000000001001111011001",
			1231 => "11111110011101100001001111011001",
			1232 => "0000001011000000000111100000001100",
			1233 => "0000000011000000001110100100000100",
			1234 => "00000000000000000001001111011001",
			1235 => "0000000000000000001100001000000100",
			1236 => "00000001001110010001001111011001",
			1237 => "00000000000000000001001111011001",
			1238 => "0000001101000000001111100100000100",
			1239 => "00000000000000000001001111011001",
			1240 => "11111111011010000001001111011001",
			1241 => "0000001100000000001000011000110000",
			1242 => "0000001101000000000111111100010100",
			1243 => "0000000110000000000100111100010000",
			1244 => "0000000100000000001111101000001000",
			1245 => "0000001001000000001010100000000100",
			1246 => "00000000000000000001001111011001",
			1247 => "00000001100100110001001111011001",
			1248 => "0000001100000000001011000000000100",
			1249 => "11111111100100010001001111011001",
			1250 => "00000000000000000001001111011001",
			1251 => "11111110101100010001001111011001",
			1252 => "0000000000000000000010101000001000",
			1253 => "0000001011000000000010001000000100",
			1254 => "00000000101110100001001111011001",
			1255 => "11111111000110010001001111011001",
			1256 => "0000001110000000001111101000001000",
			1257 => "0000000000000000001000101100000100",
			1258 => "00000010010011100001001111011001",
			1259 => "00000000000000000001001111011001",
			1260 => "0000000100000000001100001100000100",
			1261 => "11111110100110000001001111011001",
			1262 => "0000001101000000000011001000000100",
			1263 => "11111111110011000001001111011001",
			1264 => "00000001101111010001001111011001",
			1265 => "0000000001000000000100110100000100",
			1266 => "00000000110001100001001111011001",
			1267 => "0000001110000000000010111000000100",
			1268 => "11111110101101110001001111011001",
			1269 => "00000000000000000001001111011001",
			1270 => "0000000001000000001101111101000100",
			1271 => "0000001100000000000100011000001000",
			1272 => "0000000011000000000010010100000100",
			1273 => "11111110011101110001010011010101",
			1274 => "00000000000000000001010011010101",
			1275 => "0000000100000000000101000000011000",
			1276 => "0000000011000000001011111000001000",
			1277 => "0000001111000000001010001000000100",
			1278 => "00000000000000100001010011010101",
			1279 => "11111111000100010001010011010101",
			1280 => "0000000101000000000111111100001100",
			1281 => "0000000000000000000110001000000100",
			1282 => "00000000000000000001010011010101",
			1283 => "0000000001000000000001111000000100",
			1284 => "00000001011111110001010011010101",
			1285 => "00000000000000000001010011010101",
			1286 => "00000000000000000001010011010101",
			1287 => "0000001110000000001000011100010000",
			1288 => "0000001001000000001001111100001100",
			1289 => "0000001001000000001000010000000100",
			1290 => "11111111001010010001010011010101",
			1291 => "0000000101000000001100010100000100",
			1292 => "00000000100110110001010011010101",
			1293 => "00000000000000000001010011010101",
			1294 => "11111110100111110001010011010101",
			1295 => "0000001011000000000111100000001100",
			1296 => "0000000011000000001110100100000100",
			1297 => "00000000000000000001010011010101",
			1298 => "0000000000000000001100001000000100",
			1299 => "00000001001010000001010011010101",
			1300 => "00000000000000000001010011010101",
			1301 => "0000001101000000001111100100000100",
			1302 => "00000000000000000001010011010101",
			1303 => "11111111100001000001010011010101",
			1304 => "0000001100000000001000011000110000",
			1305 => "0000001101000000000100101000010100",
			1306 => "0000001010000000000111110100001000",
			1307 => "0000001001000000001010100000000100",
			1308 => "00000000000000000001010011010101",
			1309 => "00000001010010100001010011010101",
			1310 => "0000001001000000001010100100001000",
			1311 => "0000000001000000001101111100000100",
			1312 => "00000000000000000001010011010101",
			1313 => "11111110110000000001010011010101",
			1314 => "00000000000000000001010011010101",
			1315 => "0000001111000000000011000000001000",
			1316 => "0000001001000000001010100100000100",
			1317 => "00000000000000000001010011010101",
			1318 => "00000010010000000001010011010101",
			1319 => "0000000000000000000111000000001000",
			1320 => "0000000001000000001010011000000100",
			1321 => "11111110101000110001010011010101",
			1322 => "00000000000000000001010011010101",
			1323 => "0000000101000000001001010000000100",
			1324 => "11111111101010000001010011010101",
			1325 => "0000001000000000001001101000000100",
			1326 => "00000001101111110001010011010101",
			1327 => "00000000000000000001010011010101",
			1328 => "0000000001000000000100110100000100",
			1329 => "00000000100111110001010011010101",
			1330 => "0000001110000000000010111000000100",
			1331 => "11111110110100000001010011010101",
			1332 => "00000000000000000001010011010101",
			1333 => "0000001100000000001010111000001000",
			1334 => "0000000001000000001100011000000100",
			1335 => "11111110100100110001010110100001",
			1336 => "00000000000000000001010110100001",
			1337 => "0000000100000000000011001101000000",
			1338 => "0000001010000000001000010100100100",
			1339 => "0000000101000000001110101100001100",
			1340 => "0000000100000000000110101100001000",
			1341 => "0000000000000000000001010100000100",
			1342 => "00000000000000000001010110100001",
			1343 => "00000001001000010001010110100001",
			1344 => "00000000000000000001010110100001",
			1345 => "0000000000000000001111001000001000",
			1346 => "0000001011000000000100000100000100",
			1347 => "00000000000000000001010110100001",
			1348 => "11111110111100110001010110100001",
			1349 => "0000000010000000001100111000001000",
			1350 => "0000001101000000000101110000000100",
			1351 => "11111111110100110001010110100001",
			1352 => "00000001001000000001010110100001",
			1353 => "0000000000000000000010101000000100",
			1354 => "11111111001010110001010110100001",
			1355 => "00000000000000000001010110100001",
			1356 => "0000001101000000000010000100010100",
			1357 => "0000000111000000001000011000001000",
			1358 => "0000000111000000000110100100000100",
			1359 => "00000000000000000001010110100001",
			1360 => "11111111111011000001010110100001",
			1361 => "0000001010000000000001010000001000",
			1362 => "0000001101000000001001011100000100",
			1363 => "00000000000000000001010110100001",
			1364 => "00000001011111010001010110100001",
			1365 => "00000000000000000001010110100001",
			1366 => "0000001000000000001100000100000100",
			1367 => "11111111110001010001010110100001",
			1368 => "00000000000000000001010110100001",
			1369 => "0000001110000000001000110100001000",
			1370 => "0000000100000000000011001100000100",
			1371 => "00000000000000000001010110100001",
			1372 => "11111110110010100001010110100001",
			1373 => "0000000101000000001100010000010000",
			1374 => "0000001001000000001010100100001100",
			1375 => "0000000101000000001110010000000100",
			1376 => "00000000000000000001010110100001",
			1377 => "0000000010000000000011110100000100",
			1378 => "00000001001011110001010110100001",
			1379 => "00000000000000000001010110100001",
			1380 => "00000000000000000001010110100001",
			1381 => "0000000110000000001001111100000100",
			1382 => "11111110111100000001010110100001",
			1383 => "00000000000000000001010110100001",
			1384 => "0000000001000000000101011100011100",
			1385 => "0000000000000000000111000000011000",
			1386 => "0000000000000000000001010100000100",
			1387 => "11111110011001010001011001100101",
			1388 => "0000000000000000000001010100000100",
			1389 => "00000000001101010001011001100101",
			1390 => "0000000000000000000111000000001100",
			1391 => "0000000000000000000110001000000100",
			1392 => "11111110011110000001011001100101",
			1393 => "0000000000000000001111001000000100",
			1394 => "00000011111001010001011001100101",
			1395 => "11111110100000010001011001100101",
			1396 => "00000000000000000001011001100101",
			1397 => "11111110011000010001011001100101",
			1398 => "0000000001000000001100011001000000",
			1399 => "0000000101000000001001010000100000",
			1400 => "0000000100000000001011110000011100",
			1401 => "0000000001000000001101111100010000",
			1402 => "0000001000000000000110011100001000",
			1403 => "0000000010000000001100000000000100",
			1404 => "11111111011000000001011001100101",
			1405 => "11111110011010100001011001100101",
			1406 => "0000000101000000001100100100000100",
			1407 => "11111110111010000001011001100101",
			1408 => "00001010101111010001011001100101",
			1409 => "0000001000000000000110011100000100",
			1410 => "00001000111110110001011001100101",
			1411 => "0000000001000000000100110100000100",
			1412 => "11111110111101110001011001100101",
			1413 => "00000010111001000001011001100101",
			1414 => "11111110010100010001011001100101",
			1415 => "0000000110000000000100111100001100",
			1416 => "0000001011000000000101110100000100",
			1417 => "00000100011110100001011001100101",
			1418 => "0000000000000000000111000000000100",
			1419 => "11111110011001110001011001100101",
			1420 => "11111100101100100001011001100101",
			1421 => "0000000010000000001110000000001000",
			1422 => "0000000100000000001000011100000100",
			1423 => "00000000101111000001011001100101",
			1424 => "00000110111110010001011001100101",
			1425 => "0000001011000000001100100100001000",
			1426 => "0000001110000000000010010100000100",
			1427 => "11111110111011100001011001100101",
			1428 => "00000010001110010001011001100101",
			1429 => "11111111011110110001011001100101",
			1430 => "0000000011000000000001011100000100",
			1431 => "00000011101001010001011001100101",
			1432 => "11111110011000100001011001100101",
			1433 => "0000001100000000001101010100000100",
			1434 => "11111110011101010001011100010001",
			1435 => "0000001001000000001010100101000000",
			1436 => "0000001011000000000111010000010000",
			1437 => "0000000000000000000110001000001100",
			1438 => "0000000110000000000100110100000100",
			1439 => "00000000000000000001011100010001",
			1440 => "0000000111000000000011100000000100",
			1441 => "00000000000000000001011100010001",
			1442 => "00000001101000000001011100010001",
			1443 => "11111111111011110001011100010001",
			1444 => "0000001011000000000110110100011000",
			1445 => "0000001011000000000100000100001100",
			1446 => "0000000010000000000110111100001000",
			1447 => "0000000010000000001100010000000100",
			1448 => "00000000000000000001011100010001",
			1449 => "00000000010001010001011100010001",
			1450 => "00000000000000000001011100010001",
			1451 => "0000000101000000001100100100000100",
			1452 => "11111110101110100001011100010001",
			1453 => "0000000101000000000111100000000100",
			1454 => "00000000000000000001011100010001",
			1455 => "11111111011000110001011100010001",
			1456 => "0000000011000000001100111000001100",
			1457 => "0000000110000000001001100100000100",
			1458 => "11111111011010110001011100010001",
			1459 => "0000000000000000000010101000000100",
			1460 => "00000001100011010001011100010001",
			1461 => "00000000000000000001011100010001",
			1462 => "0000000111000000001111011100000100",
			1463 => "11111110011010110001011100010001",
			1464 => "0000001101000000000111010100000100",
			1465 => "00000000101000100001011100010001",
			1466 => "11111111011101010001011100010001",
			1467 => "0000001100000000001000000000010000",
			1468 => "0000001100000000001011000000001000",
			1469 => "0000001011000000000101100100000100",
			1470 => "00000000000000000001011100010001",
			1471 => "11111111010101010001011100010001",
			1472 => "0000000000000000001101010000000100",
			1473 => "00000001010011010001011100010001",
			1474 => "00000000000000000001011100010001",
			1475 => "11111110011011010001011100010001",
			1476 => "0000001100000000001101010100000100",
			1477 => "11111110100000110001011111011101",
			1478 => "0000001001000000001010100000101100",
			1479 => "0000000111000000001111011100001100",
			1480 => "0000000010000000001110010000001000",
			1481 => "0000000110000000000100110100000100",
			1482 => "00000000000000000001011111011101",
			1483 => "00000000110110100001011111011101",
			1484 => "11111110100011010001011111011101",
			1485 => "0000001101000000000111010100011000",
			1486 => "0000001110000000000110111000010000",
			1487 => "0000000111000000001011011100001000",
			1488 => "0000000000000000001000110000000100",
			1489 => "00000000111100000001011111011101",
			1490 => "11111111011100100001011111011101",
			1491 => "0000000110000000000101010000000100",
			1492 => "11111110111001000001011111011101",
			1493 => "00000000000000000001011111011101",
			1494 => "0000000000000000000011010000000100",
			1495 => "00000001001100100001011111011101",
			1496 => "00000000000000000001011111011101",
			1497 => "0000000001000000000111101000000100",
			1498 => "11111110101101100001011111011101",
			1499 => "00000000000000000001011111011101",
			1500 => "0000001100000000001000000000010100",
			1501 => "0000001001000000001010100100001000",
			1502 => "0000000110000000001111000000000100",
			1503 => "00000000110001100001011111011101",
			1504 => "11111110111101100001011111011101",
			1505 => "0000000000000000001000101100001000",
			1506 => "0000001011000000001011011100000100",
			1507 => "00000000000000000001011111011101",
			1508 => "00000001110001000001011111011101",
			1509 => "11111111111000000001011111011101",
			1510 => "0000001000000000000001110000001100",
			1511 => "0000001001000000001010100100001000",
			1512 => "0000001001000000001010100100000100",
			1513 => "11111111000100110001011111011101",
			1514 => "00000000101001110001011111011101",
			1515 => "11111110100101000001011111011101",
			1516 => "0000001101000000001110110100001100",
			1517 => "0000001000000000001100000100001000",
			1518 => "0000000001000000000100110100000100",
			1519 => "00000000100110110001011111011101",
			1520 => "00000000000000000001011111011101",
			1521 => "11111111001111100001011111011101",
			1522 => "0000001110000000001110000000000100",
			1523 => "00000000000000000001011111011101",
			1524 => "0000000001000000001100011000000100",
			1525 => "00000001101000010001011111011101",
			1526 => "00000000000000000001011111011101",
			1527 => "0000000111000000000011100000000100",
			1528 => "11111110011100000001100010010001",
			1529 => "0000001011000000001010001100010000",
			1530 => "0000001010000000000111110100001100",
			1531 => "0000000100000000001111100100001000",
			1532 => "0000001111000000001001011100000100",
			1533 => "00000000000000000001100010010001",
			1534 => "00000010001100010001100010010001",
			1535 => "00000000000000000001100010010001",
			1536 => "00000000000000000001100010010001",
			1537 => "0000000001000000001100011000110000",
			1538 => "0000001110000000000010010100011100",
			1539 => "0000000010000000001000100000010000",
			1540 => "0000000100000000000001011100001000",
			1541 => "0000001011000000000100000100000100",
			1542 => "00000000000000000001100010010001",
			1543 => "11111110101000110001100010010001",
			1544 => "0000000101000000001100100100000100",
			1545 => "11111111010010000001100010010001",
			1546 => "00000010000000000001100010010001",
			1547 => "0000001100000000001001001000000100",
			1548 => "11111110001000110001100010010001",
			1549 => "0000000111000000001111011100000100",
			1550 => "00000000010111010001100010010001",
			1551 => "11111110111000110001100010010001",
			1552 => "0000001011000000000001000000001100",
			1553 => "0000000110000000001000010000000100",
			1554 => "11111110111000100001100010010001",
			1555 => "0000001011000000001011110100000100",
			1556 => "11111111000000010001100010010001",
			1557 => "00000001001010010001100010010001",
			1558 => "0000000101000000001111010100000100",
			1559 => "00000000000000000001100010010001",
			1560 => "11111110100101000001100010010001",
			1561 => "0000000111000000000000011100010100",
			1562 => "0000001011000000000010001000001000",
			1563 => "0000000110000000001000010000000100",
			1564 => "00000000111000010001100010010001",
			1565 => "11111111010100000001100010010001",
			1566 => "0000001000000000001001101000001000",
			1567 => "0000001001000000000010101100000100",
			1568 => "00000010001010110001100010010001",
			1569 => "00000000000000000001100010010001",
			1570 => "00000000000000000001100010010001",
			1571 => "11111110101000010001100010010001",
			1572 => "0000001100000000001010111000001000",
			1573 => "0000001001000000000010101100000100",
			1574 => "11111110011010110001100100111101",
			1575 => "00000000000000000001100100111101",
			1576 => "0000001101000000001111100101001100",
			1577 => "0000001110000000000101000000111100",
			1578 => "0000000010000000001110000000100000",
			1579 => "0000000000000000000111000000010000",
			1580 => "0000001110000000001101101100001000",
			1581 => "0000000100000000001111101000000100",
			1582 => "00000000000111010001100100111101",
			1583 => "00000001101101010001100100111101",
			1584 => "0000000001000000001101111100000100",
			1585 => "00000000010101100001100100111101",
			1586 => "11111101110001010001100100111101",
			1587 => "0000001001000000001010100100001000",
			1588 => "0000000111000000000111010000000100",
			1589 => "11111110100110100001100100111101",
			1590 => "00000000111010100001100100111101",
			1591 => "0000001100000000000001101000000100",
			1592 => "00000010011100100001100100111101",
			1593 => "11111111111110010001100100111101",
			1594 => "0000001110000000001011110000010000",
			1595 => "0000000010000000001000110100001000",
			1596 => "0000000001000000000111101000000100",
			1597 => "00000000100010000001100100111101",
			1598 => "11111111010001110001100100111101",
			1599 => "0000001010000000001001000100000100",
			1600 => "00000000000000000001100100111101",
			1601 => "11111110000010100001100100111101",
			1602 => "0000001000000000001100000100000100",
			1603 => "11111110101000010001100100111101",
			1604 => "0000001000000000001001101000000100",
			1605 => "00000001000111000001100100111101",
			1606 => "11111110110000000001100100111101",
			1607 => "0000000001000000001100011000001100",
			1608 => "0000000000000000001011000100001000",
			1609 => "0000000111000000000111010000000100",
			1610 => "00000000000000000001100100111101",
			1611 => "00000001101110000001100100111101",
			1612 => "00000000000000000001100100111101",
			1613 => "11111111010001000001100100111101",
			1614 => "11111110010010110001100100111101",
			1615 => "0000000001000000001101011100000100",
			1616 => "11111110011010000001100111010011",
			1617 => "0000001001000000000010101101000000",
			1618 => "0000000110000000001011001100000100",
			1619 => "11111110100010000001100111010011",
			1620 => "0000000100000000001011110000011100",
			1621 => "0000000101000000001100100100010000",
			1622 => "0000000100000000001111100100001000",
			1623 => "0000001001000000000111101100000100",
			1624 => "00000000000000000001100111010011",
			1625 => "00000010100010000001100111010011",
			1626 => "0000001001000000001010100100000100",
			1627 => "11111110100110110001100111010011",
			1628 => "00000000001100110001100111010011",
			1629 => "0000000011000000001101101100001000",
			1630 => "0000000000000000000110001000000100",
			1631 => "11111111100011110001100111010011",
			1632 => "00000011011000100001100111010011",
			1633 => "11111111000011110001100111010011",
			1634 => "0000000000000000000111000000010000",
			1635 => "0000000011000000000001011100001000",
			1636 => "0000000110000000000100111100000100",
			1637 => "11111110111010010001100111010011",
			1638 => "00000001011111000001100111010011",
			1639 => "0000000000000000000111000000000100",
			1640 => "11111101111000000001100111010011",
			1641 => "11111111110110110001100111010011",
			1642 => "0000000000000000001000101100001000",
			1643 => "0000001010000000001000010100000100",
			1644 => "11111110111110010001100111010011",
			1645 => "00000010101110110001100111010011",
			1646 => "0000000101000000000111111100000100",
			1647 => "11111110010010010001100111010011",
			1648 => "00000000110101000001100111010011",
			1649 => "0000001101000000000100101000000100",
			1650 => "00000000100101010001100111010011",
			1651 => "11111110100000010001100111010011",
			1652 => "00000000000000000001100111010101",
			1653 => "00000000000000000001100111011001",
			1654 => "00000000000000000001100111011101",
			1655 => "00000000000000000001100111100001",
			1656 => "00000000000000000001100111100101",
			1657 => "00000000000000000001100111101001",
			1658 => "00000000000000000001100111101101",
			1659 => "00000000000000000001100111110001",
			1660 => "00000000000000000001100111110101",
			1661 => "00000000000000000001100111111001",
			1662 => "00000000000000000001100111111101",
			1663 => "00000000000000000001101000000001",
			1664 => "00000000000000000001101000000101",
			1665 => "00000000000000000001101000001001",
			1666 => "00000000000000000001101000001101",
			1667 => "00000000000000000001101000010001",
			1668 => "00000000000000000001101000010101",
			1669 => "00000000000000000001101000011001",
			1670 => "00000000000000000001101000011101",
			1671 => "00000000000000000001101000100001",
			1672 => "0000000110000000000100111100000100",
			1673 => "00000000000000000001101000110101",
			1674 => "0000000110000000001001111100000100",
			1675 => "00000000000100110001101000110101",
			1676 => "00000000000000000001101000110101",
			1677 => "0000001110000000001100001100001000",
			1678 => "0000000011000000001011101100000100",
			1679 => "00000000000000000001101001001001",
			1680 => "11111111111100010001101001001001",
			1681 => "00000000000000000001101001001001",
			1682 => "0000000110000000000100111100000100",
			1683 => "00000000000000000001101001011101",
			1684 => "0000000110000000001001111100000100",
			1685 => "00000000000101110001101001011101",
			1686 => "00000000000000000001101001011101",
			1687 => "0000001000000000001011010100001000",
			1688 => "0000001000000000001010110000000100",
			1689 => "00000000000000000001101001110001",
			1690 => "00000000000001010001101001110001",
			1691 => "00000000000000000001101001110001",
			1692 => "0000000111000000001111011100001000",
			1693 => "0000000111000000000001101000000100",
			1694 => "00000000000000000001101010001101",
			1695 => "11111111111001000001101010001101",
			1696 => "0000000111000000000100010000000100",
			1697 => "00000000001110110001101010001101",
			1698 => "00000000000000000001101010001101",
			1699 => "0000000000000000000010101000001100",
			1700 => "0000000000000000000010101000000100",
			1701 => "00000000000000000001101010101001",
			1702 => "0000001000000000000101000100000100",
			1703 => "00000000000000000001101010101001",
			1704 => "00000000001011110001101010101001",
			1705 => "11111111111101100001101010101001",
			1706 => "0000001101000000001111100100001100",
			1707 => "0000001011000000001011110100000100",
			1708 => "00000000000000000001101011000101",
			1709 => "0000001101000000000011001000000100",
			1710 => "00000000000000000001101011000101",
			1711 => "00000000000110010001101011000101",
			1712 => "00000000000000000001101011000101",
			1713 => "0000000001000000001100011000001100",
			1714 => "0000000111000000001000011000000100",
			1715 => "00000000000000000001101011100001",
			1716 => "0000000000000000000011111100000100",
			1717 => "11111111111000010001101011100001",
			1718 => "00000000000000000001101011100001",
			1719 => "00000000000000000001101011100001",
			1720 => "0000001001000000001010100000000100",
			1721 => "00000000000000000001101011111101",
			1722 => "0000000101000000000111011000001000",
			1723 => "0000001001000000000011101000000100",
			1724 => "00000000001111010001101011111101",
			1725 => "00000000000000000001101011111101",
			1726 => "00000000000000000001101011111101",
			1727 => "0000000000000000001101010000010000",
			1728 => "0000001001000000001010100000000100",
			1729 => "00000000000000000001101100100001",
			1730 => "0000001100000000001001110100001000",
			1731 => "0000001010000000001001000100000100",
			1732 => "00000000001110110001101100100001",
			1733 => "00000000000000000001101100100001",
			1734 => "00000000000000000001101100100001",
			1735 => "11111111111010110001101100100001",
			1736 => "0000000011000000000011110000010000",
			1737 => "0000000100000000001011110000000100",
			1738 => "00000000000000000001101101000101",
			1739 => "0000000001000000001100011000001000",
			1740 => "0000000001000000000111101000000100",
			1741 => "00000000000000000001101101000101",
			1742 => "11111111101011010001101101000101",
			1743 => "00000000000000000001101101000101",
			1744 => "00000000000000000001101101000101",
			1745 => "0000000100000000001000011100010000",
			1746 => "0000001001000000000000001000000100",
			1747 => "00000000000000000001101101110001",
			1748 => "0000000011000000000010010100001000",
			1749 => "0000001010000000000011101000000100",
			1750 => "00000000000000000001101101110001",
			1751 => "00000000001001000001101101110001",
			1752 => "00000000000000000001101101110001",
			1753 => "0000001001000000000100101100000100",
			1754 => "00000000000000000001101101110001",
			1755 => "11111111110111010001101101110001",
			1756 => "0000000000000000000010101000010000",
			1757 => "0000001111000000000011000000001100",
			1758 => "0000001000000000001010110000000100",
			1759 => "00000000000000000001101110011101",
			1760 => "0000001111000000001100010000000100",
			1761 => "00000000000000000001101110011101",
			1762 => "00000000001011000001101110011101",
			1763 => "00000000000000000001101110011101",
			1764 => "0000000010000000000011110100000100",
			1765 => "11111111110110110001101110011101",
			1766 => "00000000000000000001101110011101",
			1767 => "0000000000000000001010101100001100",
			1768 => "0000001001000000001010100100000100",
			1769 => "00000000000000000001101111011001",
			1770 => "0000000010000000000001011100000100",
			1771 => "00000000100011100001101111011001",
			1772 => "00000000000000000001101111011001",
			1773 => "0000001110000000001110000000001000",
			1774 => "0000000001000000001100011000000100",
			1775 => "11111111011111100001101111011001",
			1776 => "00000000000000000001101111011001",
			1777 => "0000001101000000001111100100001000",
			1778 => "0000000111000000000111010000000100",
			1779 => "00000000000000000001101111011001",
			1780 => "00000000010001010001101111011001",
			1781 => "00000000000000000001101111011001",
			1782 => "0000000111000000000001101000010100",
			1783 => "0000000000000000000010101000010000",
			1784 => "0000000011000000001100111000001100",
			1785 => "0000000111000000001000000000000100",
			1786 => "00000000000000000001110000001101",
			1787 => "0000000000000000000001010100000100",
			1788 => "00000000000000000001110000001101",
			1789 => "00000000010000110001110000001101",
			1790 => "00000000000000000001110000001101",
			1791 => "00000000000000000001110000001101",
			1792 => "0000000111000000000111010000000100",
			1793 => "11111111110001110001110000001101",
			1794 => "00000000000000000001110000001101",
			1795 => "0000001001000000001010100000000100",
			1796 => "00000000000000000001110000111001",
			1797 => "0000001100000000001000011000010000",
			1798 => "0000000110000000001001111100001100",
			1799 => "0000001001000000000011101000001000",
			1800 => "0000001001000000001010100000000100",
			1801 => "00000000000000000001110000111001",
			1802 => "00000000010000100001110000111001",
			1803 => "00000000000000000001110000111001",
			1804 => "00000000000000000001110000111001",
			1805 => "00000000000000000001110000111001",
			1806 => "0000001000000000000001010100010100",
			1807 => "0000000101000000001100100100000100",
			1808 => "00000000000000000001110001111101",
			1809 => "0000000000000000001111001000000100",
			1810 => "00000000000000000001110001111101",
			1811 => "0000001011000000000101110100001000",
			1812 => "0000000010000000001000101000000100",
			1813 => "00000000100010110001110001111101",
			1814 => "00000000000000000001110001111101",
			1815 => "00000000000000000001110001111101",
			1816 => "0000001110000000001110000000001100",
			1817 => "0000000001000000001100011000001000",
			1818 => "0000000100000000001000110100000100",
			1819 => "00000000000000000001110001111101",
			1820 => "11111111100011010001110001111101",
			1821 => "00000000000000000001110001111101",
			1822 => "00000000000000000001110001111101",
			1823 => "0000001000000000000001010100011000",
			1824 => "0000000101000000001100100100001000",
			1825 => "0000000000000000000001110000000100",
			1826 => "00000000000000000001110011010001",
			1827 => "11111111111110100001110011010001",
			1828 => "0000000000000000001111001000000100",
			1829 => "00000000000000000001110011010001",
			1830 => "0000000011000000000010010100001000",
			1831 => "0000000111000000000000011100000100",
			1832 => "00000000011100100001110011010001",
			1833 => "00000000000000000001110011010001",
			1834 => "00000000000000000001110011010001",
			1835 => "0000000101000000000111111100001000",
			1836 => "0000000100000000000110111000000100",
			1837 => "00000000000000000001110011010001",
			1838 => "11111111100110110001110011010001",
			1839 => "0000000100000000001110111000001000",
			1840 => "0000000100000000000110001100000100",
			1841 => "00000000000000000001110011010001",
			1842 => "00000000010011110001110011010001",
			1843 => "00000000000000000001110011010001",
			1844 => "0000000100000000001011110000011000",
			1845 => "0000001110000000001011101100010100",
			1846 => "0000000111000000001000000000000100",
			1847 => "00000000000000000001110100001101",
			1848 => "0000001000000000001000100100000100",
			1849 => "00000000000000000001110100001101",
			1850 => "0000001101000000001100010100001000",
			1851 => "0000001010000000001000010100000100",
			1852 => "00000000011000010001110100001101",
			1853 => "00000000000000000001110100001101",
			1854 => "00000000000000000001110100001101",
			1855 => "00000000000000000001110100001101",
			1856 => "0000001110000000000010010100000100",
			1857 => "11111111110010010001110100001101",
			1858 => "00000000000000000001110100001101",
			1859 => "0000001000000000001100000100011000",
			1860 => "0000000110000000001011001100000100",
			1861 => "00000000000000000001110101001001",
			1862 => "0000001101000000001110110100010000",
			1863 => "0000000010000000001000011100001100",
			1864 => "0000000101000000001100100100000100",
			1865 => "00000000000000000001110101001001",
			1866 => "0000001000000000001100011100000100",
			1867 => "00000000000000000001110101001001",
			1868 => "00000000010010100001110101001001",
			1869 => "00000000000000000001110101001001",
			1870 => "00000000000000000001110101001001",
			1871 => "0000000010000000000011110100000100",
			1872 => "11111111111110000001110101001001",
			1873 => "00000000000000000001110101001001",
			1874 => "0000001101000000001111100100011000",
			1875 => "0000000001000000000101011100000100",
			1876 => "00000000000000000001110101111101",
			1877 => "0000000111000000001111011100000100",
			1878 => "00000000000000000001110101111101",
			1879 => "0000000001000000000100110100001100",
			1880 => "0000001101000000000011001000000100",
			1881 => "00000000000000000001110101111101",
			1882 => "0000000110000000001000010000000100",
			1883 => "00000000000000000001110101111101",
			1884 => "00000000100100000001110101111101",
			1885 => "00000000000000000001110101111101",
			1886 => "00000000000000000001110101111101",
			1887 => "0000000101000000001001010000000100",
			1888 => "00000000000000000001110110110001",
			1889 => "0000001101000000001011111000010100",
			1890 => "0000001001000000000010101100010000",
			1891 => "0000001101000000001110010000000100",
			1892 => "00000000000000000001110110110001",
			1893 => "0000000110000000001001100100000100",
			1894 => "00000000000000000001110110110001",
			1895 => "0000001010000000000110011100000100",
			1896 => "00000000010110110001110110110001",
			1897 => "00000000000000000001110110110001",
			1898 => "00000000000000000001110110110001",
			1899 => "00000000000000000001110110110001",
			1900 => "0000000000000000001010101100011000",
			1901 => "0000001011000000000101110100010100",
			1902 => "0000001100000000001001110100010000",
			1903 => "0000000110000000000100110100000100",
			1904 => "00000000000000000001110111111101",
			1905 => "0000001100000000001010111000000100",
			1906 => "00000000000000000001110111111101",
			1907 => "0000000010000000001000101000000100",
			1908 => "00000000011001110001110111111101",
			1909 => "00000000000000000001110111111101",
			1910 => "00000000000000000001110111111101",
			1911 => "00000000000000000001110111111101",
			1912 => "0000000110000000001000010000000100",
			1913 => "11111111110100000001110111111101",
			1914 => "0000001010000000001010110000001000",
			1915 => "0000001010000000001001000100000100",
			1916 => "00000000000000000001110111111101",
			1917 => "00000000001011010001110111111101",
			1918 => "00000000000000000001110111111101",
			1919 => "0000000111000000001000011000100000",
			1920 => "0000001100000000000100011000001100",
			1921 => "0000000100000000001000100000000100",
			1922 => "00000000000000000001111001011001",
			1923 => "0000000001000000001100011000000100",
			1924 => "11111111101110110001111001011001",
			1925 => "00000000000000000001111001011001",
			1926 => "0000001100000000001000000000010000",
			1927 => "0000000000000000001000101100001100",
			1928 => "0000000111000000000110100100000100",
			1929 => "00000000000000000001111001011001",
			1930 => "0000000110000000000100110100000100",
			1931 => "00000000000000000001111001011001",
			1932 => "00000000101010000001111001011001",
			1933 => "00000000000000000001111001011001",
			1934 => "00000000000000000001111001011001",
			1935 => "0000000010000000000011110100001100",
			1936 => "0000000001000000000111101000000100",
			1937 => "00000000000000000001111001011001",
			1938 => "0000000110000000001001111100000100",
			1939 => "11111111011001010001111001011001",
			1940 => "00000000000000000001111001011001",
			1941 => "00000000000000000001111001011001",
			1942 => "0000000100000000001110111000100000",
			1943 => "0000001011000000001011011100001000",
			1944 => "0000000100000000001011101100000100",
			1945 => "00000000000000000001111010100101",
			1946 => "11111111110010100001111010100101",
			1947 => "0000000111000000000100010000010100",
			1948 => "0000000110000000001001100100000100",
			1949 => "00000000000000000001111010100101",
			1950 => "0000001001000000000011101000001100",
			1951 => "0000001100000000000100011000000100",
			1952 => "00000000000000000001111010100101",
			1953 => "0000001000000000001011010100000100",
			1954 => "00000000100011110001111010100101",
			1955 => "00000000000000000001111010100101",
			1956 => "00000000000000000001111010100101",
			1957 => "00000000000000000001111010100101",
			1958 => "0000001010000000001100011100000100",
			1959 => "11111111110011000001111010100101",
			1960 => "00000000000000000001111010100101",
			1961 => "0000001100000000001011000000001000",
			1962 => "0000001110000000001000101000000100",
			1963 => "11111111010011010001111011101001",
			1964 => "00000000000000000001111011101001",
			1965 => "0000001101000000001111100100011000",
			1966 => "0000001011000000000010001000000100",
			1967 => "00000000000000000001111011101001",
			1968 => "0000000100000000001011110000000100",
			1969 => "00000000000000000001111011101001",
			1970 => "0000001011000000000010110100001100",
			1971 => "0000000100000000001001001100001000",
			1972 => "0000001101000000001010001000000100",
			1973 => "00000000000000000001111011101001",
			1974 => "00000000011111010001111011101001",
			1975 => "00000000000000000001111011101001",
			1976 => "00000000000000000001111011101001",
			1977 => "11111111111000000001111011101001",
			1978 => "0000000000000000000010101000010100",
			1979 => "0000001001000000000000001000000100",
			1980 => "00000000000000000001111101001101",
			1981 => "0000000111000000001000011000001100",
			1982 => "0000000010000000001000101000001000",
			1983 => "0000001110000000000110010000000100",
			1984 => "00000000000000000001111101001101",
			1985 => "00000000110111110001111101001101",
			1986 => "00000000000000000001111101001101",
			1987 => "00000000000000000001111101001101",
			1988 => "0000000111000000001111011100000100",
			1989 => "11111111000111100001111101001101",
			1990 => "0000000111000000000101100100001100",
			1991 => "0000001000000000001011010100001000",
			1992 => "0000001001000000000010101100000100",
			1993 => "00000000100110100001111101001101",
			1994 => "00000000000000000001111101001101",
			1995 => "00000000000000000001111101001101",
			1996 => "0000000110000000000101010000001000",
			1997 => "0000000100000000000110001100000100",
			1998 => "00000000000000000001111101001101",
			1999 => "11111111101011000001111101001101",
			2000 => "0000000110000000001001111100000100",
			2001 => "00000000000100100001111101001101",
			2002 => "00000000000000000001111101001101",
			2003 => "0000001000000000000110011100010100",
			2004 => "0000001010000000000011101000000100",
			2005 => "00000000000000000001111111000001",
			2006 => "0000001010000000000111110100001100",
			2007 => "0000000110000000001111000000001000",
			2008 => "0000000110000000001011001100000100",
			2009 => "00000000000000000001111111000001",
			2010 => "00000000000111010001111111000001",
			2011 => "00000000000000000001111111000001",
			2012 => "00000000000000000001111111000001",
			2013 => "0000000110000000001000010000001100",
			2014 => "0000001001000000001010100100001000",
			2015 => "0000000001000000000001000100000100",
			2016 => "00000000000000000001111111000001",
			2017 => "11111111001000110001111111000001",
			2018 => "00000000000000000001111111000001",
			2019 => "0000000100000000001001001100010000",
			2020 => "0000000111000000001000011000000100",
			2021 => "00000000000000000001111111000001",
			2022 => "0000001000000000001001101000001000",
			2023 => "0000001010000000001000010100000100",
			2024 => "00000000000000000001111111000001",
			2025 => "00000000011001100001111111000001",
			2026 => "00000000000000000001111111000001",
			2027 => "0000001010000000001010110000001000",
			2028 => "0000000100000000001110111000000100",
			2029 => "00000000000000000001111111000001",
			2030 => "11111111101101100001111111000001",
			2031 => "00000000000000000001111111000001",
			2032 => "0000000111000000001000011000100000",
			2033 => "0000001000000000000001110000011000",
			2034 => "0000001100000000001000000000010100",
			2035 => "0000001100000000000100011000000100",
			2036 => "00000000000000000010000000110101",
			2037 => "0000000110000000001000010000001100",
			2038 => "0000000111000000000110100100000100",
			2039 => "00000000000000000010000000110101",
			2040 => "0000000110000000000100110100000100",
			2041 => "00000000000000000010000000110101",
			2042 => "00000000101000100010000000110101",
			2043 => "00000000000000000010000000110101",
			2044 => "00000000000000000010000000110101",
			2045 => "0000001011000000000101110100000100",
			2046 => "11111111111101010010000000110101",
			2047 => "00000000000000000010000000110101",
			2048 => "0000001110000000001111101000001100",
			2049 => "0000000001000000001100011000001000",
			2050 => "0000000111000000000111010000000100",
			2051 => "11111111001001100010000000110101",
			2052 => "00000000000000000010000000110101",
			2053 => "00000000000000000010000000110101",
			2054 => "0000001011000000000001000000001100",
			2055 => "0000000111000000001111011100000100",
			2056 => "00000000000000000010000000110101",
			2057 => "0000000101000000001001010000000100",
			2058 => "00000000000000000010000000110101",
			2059 => "00000000010001000010000000110101",
			2060 => "11111111101101010010000000110101",
			2061 => "0000001001000000000111101100001100",
			2062 => "0000001100000000001000000000001000",
			2063 => "0000001110000000001000101000000100",
			2064 => "11111111001001010010000010100001",
			2065 => "00000000000000000010000010100001",
			2066 => "00000000000000000010000010100001",
			2067 => "0000001100000000000100011000010000",
			2068 => "0000001000000000000001010100001100",
			2069 => "0000001001000000000000001000000100",
			2070 => "00000000000000000010000010100001",
			2071 => "0000001110000000000110010000000100",
			2072 => "00000000000000000010000010100001",
			2073 => "00000000110100000010000010100001",
			2074 => "00000000000000000010000010100001",
			2075 => "0000000110000000001000010000001000",
			2076 => "0000000011000000001000100000000100",
			2077 => "00000000000000000010000010100001",
			2078 => "11111111011110110010000010100001",
			2079 => "0000001011000000000001000000010000",
			2080 => "0000000101000000000010011100000100",
			2081 => "00000000000000000010000010100001",
			2082 => "0000001110000000000011000000000100",
			2083 => "00000000000000000010000010100001",
			2084 => "0000001010000000000110011100000100",
			2085 => "00000000110110010010000010100001",
			2086 => "00000000000000000010000010100001",
			2087 => "11111111111010110010000010100001",
			2088 => "0000001000000000000001110000011100",
			2089 => "0000001101000000001100010100010100",
			2090 => "0000001100000000000100011000000100",
			2091 => "00000000000000000010000100010101",
			2092 => "0000001101000000000101110000000100",
			2093 => "00000000000000000010000100010101",
			2094 => "0000000000000000000111000100000100",
			2095 => "00000000000000000010000100010101",
			2096 => "0000000110000000001000010000000100",
			2097 => "00000000111011010010000100010101",
			2098 => "00000000000000000010000100010101",
			2099 => "0000000110000000000100111100000100",
			2100 => "11111111101010110010000100010101",
			2101 => "00000000000000000010000100010101",
			2102 => "0000000111000000001111011100000100",
			2103 => "11111111001010010010000100010101",
			2104 => "0000000001000000000100110100010100",
			2105 => "0000000001000000001110010100001000",
			2106 => "0000000101000000001110110100000100",
			2107 => "00000000000000000010000100010101",
			2108 => "11111111111001000010000100010101",
			2109 => "0000001110000000000011000000000100",
			2110 => "00000000000000000010000100010101",
			2111 => "0000000101000000000101110000000100",
			2112 => "00000000000000000010000100010101",
			2113 => "00000000110000010010000100010101",
			2114 => "0000001111000000001000110100000100",
			2115 => "00000000000000000010000100010101",
			2116 => "11111111110011110010000100010101",
			2117 => "0000001000000000000110011100010100",
			2118 => "0000001010000000000011101000000100",
			2119 => "00000000000000000010000110010001",
			2120 => "0000001010000000000111110100001100",
			2121 => "0000000110000000001111000000001000",
			2122 => "0000000110000000001011001100000100",
			2123 => "00000000000000000010000110010001",
			2124 => "00000000000111110010000110010001",
			2125 => "00000000000000000010000110010001",
			2126 => "00000000000000000010000110010001",
			2127 => "0000000110000000001000010000001100",
			2128 => "0000001001000000001010100100001000",
			2129 => "0000001001000000000101010000000100",
			2130 => "00000000000000000010000110010001",
			2131 => "11111111000101110010000110010001",
			2132 => "00000000000000000010000110010001",
			2133 => "0000000000000000001101010000010100",
			2134 => "0000000111000000001000011000000100",
			2135 => "00000000000000000010000110010001",
			2136 => "0000000000000000000111000000000100",
			2137 => "00000000000000000010000110010001",
			2138 => "0000000101000000001001010000000100",
			2139 => "00000000000000000010000110010001",
			2140 => "0000001000000000000001110000000100",
			2141 => "00000000000000000010000110010001",
			2142 => "00000000100001010010000110010001",
			2143 => "0000000000000000000011111100001000",
			2144 => "0000001010000000001100011100000100",
			2145 => "11111111101100000010000110010001",
			2146 => "00000000000000000010000110010001",
			2147 => "00000000000000000010000110010001",
			2148 => "0000001000000000000001110000101000",
			2149 => "0000000111000000000001101000010100",
			2150 => "0000001001000000000000001000000100",
			2151 => "00000000000000000010001000011101",
			2152 => "0000000000000000001010101100001100",
			2153 => "0000000011000000001100111000001000",
			2154 => "0000001110000000000110010000000100",
			2155 => "00000000000000000010001000011101",
			2156 => "00000000110101000010001000011101",
			2157 => "00000000000000000010001000011101",
			2158 => "00000000000000000010001000011101",
			2159 => "0000000000000000000111000000001100",
			2160 => "0000000111000000000111010000001000",
			2161 => "0000001011000000000000011100000100",
			2162 => "00000000000000000010001000011101",
			2163 => "11111111010101110010001000011101",
			2164 => "00000000000000000010001000011101",
			2165 => "0000001110000000000110111000000100",
			2166 => "00000000100111000010001000011101",
			2167 => "00000000000000000010001000011101",
			2168 => "0000000111000000001111011100000100",
			2169 => "11111111000110110010001000011101",
			2170 => "0000000001000000000100110100010100",
			2171 => "0000000001000000001110010100001000",
			2172 => "0000000101000000001110110100000100",
			2173 => "00000000000000000010001000011101",
			2174 => "11111111110101110010001000011101",
			2175 => "0000001110000000000011000000000100",
			2176 => "00000000000000000010001000011101",
			2177 => "0000000101000000000101110000000100",
			2178 => "00000000000000000010001000011101",
			2179 => "00000000110011000010001000011101",
			2180 => "0000001111000000001000110100000100",
			2181 => "00000000000000000010001000011101",
			2182 => "11111111110001100010001000011101",
			2183 => "0000000001000000000001111000010000",
			2184 => "0000001110000000000001011100001100",
			2185 => "0000000100000000001100010000000100",
			2186 => "00000000000000000010001010100001",
			2187 => "0000001100000000001111011100000100",
			2188 => "11111111001001000010001010100001",
			2189 => "00000000000000000010001010100001",
			2190 => "00000000000000000010001010100001",
			2191 => "0000001110000000001011101100010000",
			2192 => "0000000111000000000110100100000100",
			2193 => "00000000000000000010001010100001",
			2194 => "0000000000000000000111000100000100",
			2195 => "00000000000000000010001010100001",
			2196 => "0000000000000000000010101000000100",
			2197 => "00000000110000100010001010100001",
			2198 => "00000000000000000010001010100001",
			2199 => "0000000000000000000111000000001000",
			2200 => "0000001000000000000001010100000100",
			2201 => "00000000000000000010001010100001",
			2202 => "11111111100100110010001010100001",
			2203 => "0000000111000000000101100100010000",
			2204 => "0000000100000000001110111000001100",
			2205 => "0000001101000000001010001000000100",
			2206 => "00000000000000000010001010100001",
			2207 => "0000000111000000001000011000000100",
			2208 => "00000000000000000010001010100001",
			2209 => "00000000101001010010001010100001",
			2210 => "00000000000000000010001010100001",
			2211 => "0000000100000000001110111000001000",
			2212 => "0000000111000000001011011100000100",
			2213 => "00000000000000000010001010100001",
			2214 => "11111111011101000010001010100001",
			2215 => "00000000000000000010001010100001",
			2216 => "0000000100000000001011110000010000",
			2217 => "0000001110000000001011101100001100",
			2218 => "0000001011000000000110110100001000",
			2219 => "0000001001000000001010100000000100",
			2220 => "00000000000000000010001100001101",
			2221 => "00000000111110100010001100001101",
			2222 => "00000000000000000010001100001101",
			2223 => "00000000000000000010001100001101",
			2224 => "0000000101000000001001010000000100",
			2225 => "11111110111100100010001100001101",
			2226 => "0000001011000000000001000000100000",
			2227 => "0000000000000000000111000000001100",
			2228 => "0000001110000000001000101000000100",
			2229 => "00000000000000000010001100001101",
			2230 => "0000000000000000000111000000000100",
			2231 => "11111111101100110010001100001101",
			2232 => "00000000000000000010001100001101",
			2233 => "0000001110000000001000101000000100",
			2234 => "00000000000000000010001100001101",
			2235 => "0000000000000000000010011000001000",
			2236 => "0000001001000000000010101100000100",
			2237 => "00000000111100000010001100001101",
			2238 => "00000000000000000010001100001101",
			2239 => "0000001110000000000011110000000100",
			2240 => "11111111101101100010001100001101",
			2241 => "00000000011011000010001100001101",
			2242 => "11111111011100100010001100001101",
			2243 => "0000000111000000000001101000010100",
			2244 => "0000000100000000001000100000001100",
			2245 => "0000001010000000001010100000000100",
			2246 => "00000000000000000010001110111001",
			2247 => "0000001100000000001101010100000100",
			2248 => "00000000000000000010001110111001",
			2249 => "00000000001111110010001110111001",
			2250 => "0000001001000000000010101100000100",
			2251 => "11111110101101010010001110111001",
			2252 => "00000000000000000010001110111001",
			2253 => "0000001100000000001001110100011000",
			2254 => "0000001011000000000110110100001000",
			2255 => "0000000011000000001011111000000100",
			2256 => "00000000000000000010001110111001",
			2257 => "11111111101100110010001110111001",
			2258 => "0000001000000000001100000100001000",
			2259 => "0000000100000000001111101000000100",
			2260 => "00000000000000000010001110111001",
			2261 => "00000001010001000010001110111001",
			2262 => "0000001100000000001001110100000100",
			2263 => "11111111111011110010001110111001",
			2264 => "00000000000000000010001110111001",
			2265 => "0000001110000000001000011100011000",
			2266 => "0000001001000000000100101100001100",
			2267 => "0000000100000000001101001000001000",
			2268 => "0000000100000000001000110100000100",
			2269 => "00000000000000000010001110111001",
			2270 => "00000000001100010010001110111001",
			2271 => "11111111101100100010001110111001",
			2272 => "0000000101000000000010011100000100",
			2273 => "00000000000000000010001110111001",
			2274 => "0000001110000000001110000000000100",
			2275 => "11111111000100010010001110111001",
			2276 => "00000000000000000010001110111001",
			2277 => "0000001011000000000111100000010000",
			2278 => "0000001000000000000110001000001100",
			2279 => "0000001001000000000010101100001000",
			2280 => "0000000100000000000010111000000100",
			2281 => "00000000000000000010001110111001",
			2282 => "00000001001110110010001110111001",
			2283 => "00000000000000000010001110111001",
			2284 => "00000000000000000010001110111001",
			2285 => "11111111111010000010001110111001",
			2286 => "0000001001000000001010100000011000",
			2287 => "0000001110000000001011110000001000",
			2288 => "0000000000000000001000101100000100",
			2289 => "00000000000000000010010000111101",
			2290 => "11111111000000000010010000111101",
			2291 => "0000000100000000000011110100001100",
			2292 => "0000000000000000001000110000000100",
			2293 => "00000000000000000010010000111101",
			2294 => "0000000101000000001110010000000100",
			2295 => "00000000000000000010010000111101",
			2296 => "00000000010111110010010000111101",
			2297 => "00000000000000000010010000111101",
			2298 => "0000001100000000001011011100101000",
			2299 => "0000001011000000001011011100001000",
			2300 => "0000000100000000000011000000000100",
			2301 => "00000000000000000010010000111101",
			2302 => "11111111101110010010010000111101",
			2303 => "0000000000000000000111000100000100",
			2304 => "00000000000000000010010000111101",
			2305 => "0000001110000000001111101000001100",
			2306 => "0000000111000000001111011100001000",
			2307 => "0000001100000000000100011000000100",
			2308 => "00000000000000000010010000111101",
			2309 => "00000001000101100010010000111101",
			2310 => "00000000000000000010010000111101",
			2311 => "0000001110000000000110001100001000",
			2312 => "0000001001000000001010100100000100",
			2313 => "00000000000000000010010000111101",
			2314 => "11111111100001010010010000111101",
			2315 => "0000001001000000000010101100000100",
			2316 => "00000000111011000010010000111101",
			2317 => "00000000000000000010010000111101",
			2318 => "11111111101110010010010000111101",
			2319 => "0000001001000000001010100000101100",
			2320 => "0000000111000000001111011100001000",
			2321 => "0000000100000000000110101100000100",
			2322 => "00000000000000000010010011110001",
			2323 => "11111110101111000010010011110001",
			2324 => "0000001011000000000010110100010100",
			2325 => "0000000100000000000011001100010000",
			2326 => "0000001111000000000000010000000100",
			2327 => "00000000000000000010010011110001",
			2328 => "0000001000000000001100011100000100",
			2329 => "00000000000000000010010011110001",
			2330 => "0000000101000000001100010100000100",
			2331 => "00000000101101010010010011110001",
			2332 => "00000000000000000010010011110001",
			2333 => "00000000000000000010010011110001",
			2334 => "0000001100000000001111011100000100",
			2335 => "00000000000000000010010011110001",
			2336 => "0000001000000000001011010100001000",
			2337 => "0000000111000000000010001000000100",
			2338 => "00000000000000000010010011110001",
			2339 => "11111111100101110010010011110001",
			2340 => "00000000000000000010010011110001",
			2341 => "0000001100000000001001110100011100",
			2342 => "0000000000000000001000101100011000",
			2343 => "0000000101000000001100100100001000",
			2344 => "0000001100000000001010111000000100",
			2345 => "00000000010000000010010011110001",
			2346 => "00000000000000000010010011110001",
			2347 => "0000001100000000000100011000000100",
			2348 => "00000000000000000010010011110001",
			2349 => "0000000001000000001101111100000100",
			2350 => "00000000000000000010010011110001",
			2351 => "0000001001000000001010100000000100",
			2352 => "00000000000000000010010011110001",
			2353 => "00000001010010100010010011110001",
			2354 => "00000000000000000010010011110001",
			2355 => "0000000001000000000100110100001100",
			2356 => "0000000110000000001000010000000100",
			2357 => "00000000000000000010010011110001",
			2358 => "0000000101000000000111111100000100",
			2359 => "00000000000000000010010011110001",
			2360 => "00000000100110110010010011110001",
			2361 => "0000001011000000000101110100000100",
			2362 => "00000000000000000010010011110001",
			2363 => "11111111001000110010010011110001",
			2364 => "0000001110000000001110110100010000",
			2365 => "0000000111000000000110100100000100",
			2366 => "11111110011011100010010101110101",
			2367 => "0000000111000000000110100100001000",
			2368 => "0000001101000000000001000000000100",
			2369 => "00000000111000100010010101110101",
			2370 => "00000000000000000010010101110101",
			2371 => "11111111001000010010010101110101",
			2372 => "0000001101000000001111100100110000",
			2373 => "0000001110000000000110001100011100",
			2374 => "0000001000000000001001101000010100",
			2375 => "0000001010000000000011101000000100",
			2376 => "11111110110111100010010101110101",
			2377 => "0000000010000000001000100000001000",
			2378 => "0000000110000000001001100100000100",
			2379 => "00000001110010100010010101110101",
			2380 => "00000000000000000010010101110101",
			2381 => "0000000000000000000111000000000100",
			2382 => "11111111010001100010010101110101",
			2383 => "00000000101010010010010101110101",
			2384 => "0000001110000000001100001100000100",
			2385 => "11111110101010110010010101110101",
			2386 => "00000000000000000010010101110101",
			2387 => "0000001000000000000111000100010000",
			2388 => "0000000100000000001001001100000100",
			2389 => "00000000000000000010010101110101",
			2390 => "0000000001000000001010011000001000",
			2391 => "0000001101000000001100000000000100",
			2392 => "00000011110111110010010101110101",
			2393 => "00000001101000010010010101110101",
			2394 => "00000000000000000010010101110101",
			2395 => "00000000000000000010010101110101",
			2396 => "11111110100110110010010101110101",
			2397 => "0000000000000000000010101000011000",
			2398 => "0000000001000000000001111000000100",
			2399 => "00000000000000000010011000001001",
			2400 => "0000000111000000001000011000010000",
			2401 => "0000000010000000001000101000001100",
			2402 => "0000001010000000000011101000000100",
			2403 => "00000000000000000010011000001001",
			2404 => "0000001110000000000110010000000100",
			2405 => "00000000000000000010011000001001",
			2406 => "00000000111001110010011000001001",
			2407 => "00000000000000000010011000001001",
			2408 => "00000000000000000010011000001001",
			2409 => "0000000111000000001111011100000100",
			2410 => "11111111000100100010011000001001",
			2411 => "0000000111000000000101100100010000",
			2412 => "0000001000000000001011010100001100",
			2413 => "0000001000000000000001010100000100",
			2414 => "00000000000000000010011000001001",
			2415 => "0000000001000000001100011000000100",
			2416 => "00000000101100010010011000001001",
			2417 => "00000000000000000010011000001001",
			2418 => "00000000000000000010011000001001",
			2419 => "0000001110000000001000011100010000",
			2420 => "0000000100000000000110001100000100",
			2421 => "00000000000000000010011000001001",
			2422 => "0000000110000000000101010000001000",
			2423 => "0000001100000000000001011000000100",
			2424 => "11111111100111010010011000001001",
			2425 => "00000000000000000010011000001001",
			2426 => "00000000000000000010011000001001",
			2427 => "0000001101000000001011111000001100",
			2428 => "0000000110000000001001111100001000",
			2429 => "0000000110000000001000010000000100",
			2430 => "00000000000000000010011000001001",
			2431 => "00000000100001000010011000001001",
			2432 => "00000000000000000010011000001001",
			2433 => "00000000000000000010011000001001",
			2434 => "0000000100000000001011110000011100",
			2435 => "0000001110000000001011101100011000",
			2436 => "0000000110000000000100110100000100",
			2437 => "00000000000000000010011010001101",
			2438 => "0000001011000000000110110100010000",
			2439 => "0000001001000000001010100000001100",
			2440 => "0000000010000000000110111100001000",
			2441 => "0000000000000000000110001000000100",
			2442 => "00000000010101100010011010001101",
			2443 => "00000000000000000010011010001101",
			2444 => "00000000000000000010011010001101",
			2445 => "00000001000001000010011010001101",
			2446 => "00000000000000000010011010001101",
			2447 => "00000000000000000010011010001101",
			2448 => "0000000110000000000100111100000100",
			2449 => "11111110111101110010011010001101",
			2450 => "0000001011000000000001000000100000",
			2451 => "0000000101000000000111111100010000",
			2452 => "0000000100000000000110001100001100",
			2453 => "0000001001000000000010101100001000",
			2454 => "0000001101000000001110010000000100",
			2455 => "00000000000000000010011010001101",
			2456 => "00000000011111010010011010001101",
			2457 => "00000000000000000010011010001101",
			2458 => "11111111101100000010011010001101",
			2459 => "0000000110000000001001111100001100",
			2460 => "0000001001000000000010101100001000",
			2461 => "0000000001000000000101011100000100",
			2462 => "00000000000000000010011010001101",
			2463 => "00000000101110010010011010001101",
			2464 => "00000000000000000010011010001101",
			2465 => "00000000000000000010011010001101",
			2466 => "11111111100001110010011010001101",
			2467 => "0000001100000000001000000000100000",
			2468 => "0000000001000000000001111000001000",
			2469 => "0000001110000000001111101000000100",
			2470 => "11111111000101000010011100100001",
			2471 => "00000000000000000010011100100001",
			2472 => "0000001011000000000110110100001000",
			2473 => "0000001011000000000100000100000100",
			2474 => "00000000000000000010011100100001",
			2475 => "11111111110100110010011100100001",
			2476 => "0000001011000000000100010000001100",
			2477 => "0000000001000000001100011000001000",
			2478 => "0000000101000000000111100000000100",
			2479 => "00000000000000000010011100100001",
			2480 => "00000000010100110010011100100001",
			2481 => "00000000000000000010011100100001",
			2482 => "00000000000000000010011100100001",
			2483 => "0000000101000000000110111100101000",
			2484 => "0000000001000000001010011000100100",
			2485 => "0000000000000000001111001000000100",
			2486 => "00000000000000000010011100100001",
			2487 => "0000000111000000000101100100010000",
			2488 => "0000000110000000001000010000001000",
			2489 => "0000000100000000000011001100000100",
			2490 => "00000000110110010010011100100001",
			2491 => "00000000000000000010011100100001",
			2492 => "0000001011000000001010010100000100",
			2493 => "00000000000000000010011100100001",
			2494 => "00000000000000110010011100100001",
			2495 => "0000001110000000001000011100001000",
			2496 => "0000000110000000001000010000000100",
			2497 => "11111111101001100010011100100001",
			2498 => "00000000000000000010011100100001",
			2499 => "0000000110000000001001111100000100",
			2500 => "00000000100111010010011100100001",
			2501 => "00000000000000000010011100100001",
			2502 => "00000000000000000010011100100001",
			2503 => "11111111011101010010011100100001",
			2504 => "0000001001000000001010100000101100",
			2505 => "0000001100000000001011000000001000",
			2506 => "0000000100000000000110101100000100",
			2507 => "00000000000000000010011111001101",
			2508 => "11111111001101000010011111001101",
			2509 => "0000000010000000000010010100001100",
			2510 => "0000001000000000001000100100000100",
			2511 => "00000000000000000010011111001101",
			2512 => "0000000100000000001000011100000100",
			2513 => "00000000000111010010011111001101",
			2514 => "00000000000000000010011111001101",
			2515 => "0000001110000000001011110000001000",
			2516 => "0000001111000000001000110100000100",
			2517 => "00000000000000000010011111001101",
			2518 => "11111111011111000010011111001101",
			2519 => "0000000011000000000100001100001100",
			2520 => "0000001110000000001000000100000100",
			2521 => "00000000000000000010011111001101",
			2522 => "0000001111000000001111100000000100",
			2523 => "00000000010001000010011111001101",
			2524 => "00000000000000000010011111001101",
			2525 => "00000000000000000010011111001101",
			2526 => "0000001100000000001011011100101000",
			2527 => "0000001011000000001011011100001000",
			2528 => "0000000100000000000011000000000100",
			2529 => "00000000000000000010011111001101",
			2530 => "11111111110001100010011111001101",
			2531 => "0000000100000000000110111000000100",
			2532 => "00000000000000000010011111001101",
			2533 => "0000001110000000001111101000001100",
			2534 => "0000000111000000001111011100001000",
			2535 => "0000001100000000000100011000000100",
			2536 => "00000000000000000010011111001101",
			2537 => "00000001000110100010011111001101",
			2538 => "00000000000000000010011111001101",
			2539 => "0000001110000000000110001100001000",
			2540 => "0000000001000000001100011000000100",
			2541 => "00000000000000000010011111001101",
			2542 => "11111111011001010010011111001101",
			2543 => "0000000001000000001100011000000100",
			2544 => "00000000110101010010011111001101",
			2545 => "00000000000000000010011111001101",
			2546 => "11111111110001010010011111001101",
			2547 => "0000001100000000001101010100000100",
			2548 => "11111110101111010010100001010001",
			2549 => "0000001100000000000001011000110100",
			2550 => "0000000011000000000011110000101000",
			2551 => "0000000111000000000001101000010000",
			2552 => "0000000000000000000010101000001100",
			2553 => "0000001001000000000000001000000100",
			2554 => "00000000000000000010100001010001",
			2555 => "0000000011000000001100111000000100",
			2556 => "00000001001001110010100001010001",
			2557 => "00000000000000000010100001010001",
			2558 => "11111111100111110010100001010001",
			2559 => "0000000100000000001010110100010000",
			2560 => "0000000111000000000111010000001000",
			2561 => "0000001001000000001010100100000100",
			2562 => "11111110110010110010100001010001",
			2563 => "00000000001000110010100001010001",
			2564 => "0000001001000000001010100100000100",
			2565 => "00000000110000110010100001010001",
			2566 => "11111111110101010010100001010001",
			2567 => "0000001110000000001000011100000100",
			2568 => "11111110111110110010100001010001",
			2569 => "00000000000000000010100001010001",
			2570 => "0000001001000000000010101100001000",
			2571 => "0000000000000000001011000100000100",
			2572 => "00000001001101010010100001010001",
			2573 => "00000000000000000010100001010001",
			2574 => "00000000000000000010100001010001",
			2575 => "0000000111000000000100010000000100",
			2576 => "00000000000000000010100001010001",
			2577 => "0000001010000000001010110000000100",
			2578 => "11111110111110000010100001010001",
			2579 => "00000000000000000010100001010001",
			2580 => "0000001001000000001010100000111100",
			2581 => "0000000111000000001111011100011000",
			2582 => "0000000100000000001111100100010100",
			2583 => "0000001011000000000100000100010000",
			2584 => "0000000101000000000001001000000100",
			2585 => "00000000000000000010100100101101",
			2586 => "0000000000000000000001010100000100",
			2587 => "00000000000000000010100100101101",
			2588 => "0000000111000000001000000000000100",
			2589 => "00000000000000000010100100101101",
			2590 => "00000001000111100010100100101101",
			2591 => "11111111111011110010100100101101",
			2592 => "11111110011110000010100100101101",
			2593 => "0000001101000000000111010100011100",
			2594 => "0000000110000000001000010000001100",
			2595 => "0000000111000000000101100100001000",
			2596 => "0000000110000000001001100100000100",
			2597 => "00000000000000000010100100101101",
			2598 => "00000000101001100010100100101101",
			2599 => "11111111001001010010100100101101",
			2600 => "0000000100000000000011101100001000",
			2601 => "0000000101000000000111111100000100",
			2602 => "00000000000000000010100100101101",
			2603 => "00000001001100100010100100101101",
			2604 => "0000001011000000001101000100000100",
			2605 => "11111111110111100010100100101101",
			2606 => "00000000000000000010100100101101",
			2607 => "0000000110000000001001111100000100",
			2608 => "11111110111010000010100100101101",
			2609 => "00000000000000000010100100101101",
			2610 => "0000000011000000001101101100010000",
			2611 => "0000000000000000001010101100001100",
			2612 => "0000001011000000001011011100001000",
			2613 => "0000001011000000000000011100000100",
			2614 => "00000000101010100010100100101101",
			2615 => "00000000000000000010100100101101",
			2616 => "00000001101101010010100100101101",
			2617 => "00000000000000000010100100101101",
			2618 => "0000000000000000000010101000000100",
			2619 => "11111111001010110010100100101101",
			2620 => "0000000000000000001101010000010100",
			2621 => "0000001001000000000010101100001100",
			2622 => "0000001101000000001010001000000100",
			2623 => "00000000000000000010100100101101",
			2624 => "0000000111000000000101100100000100",
			2625 => "00000001011010110010100100101101",
			2626 => "00000000000000000010100100101101",
			2627 => "0000001100000000001000000000000100",
			2628 => "00000000000011100010100100101101",
			2629 => "11111111010000110010100100101101",
			2630 => "0000000011000000000011110000001000",
			2631 => "0000000000000000001101010000000100",
			2632 => "00000000000000000010100100101101",
			2633 => "11111111001001100010100100101101",
			2634 => "00000000000000000010100100101101",
			2635 => "0000001001000000001010100000111100",
			2636 => "0000000111000000001111011100011000",
			2637 => "0000000100000000001111100100010100",
			2638 => "0000001011000000000100000100010000",
			2639 => "0000000101000000000001001000000100",
			2640 => "00000000000000000010101000001001",
			2641 => "0000000000000000000001010100000100",
			2642 => "00000000000000000010101000001001",
			2643 => "0000000111000000001000000000000100",
			2644 => "00000000000000000010101000001001",
			2645 => "00000001010001010010101000001001",
			2646 => "11111111110011000010101000001001",
			2647 => "11111110011100010010101000001001",
			2648 => "0000001101000000000111010100011100",
			2649 => "0000000110000000001000010000001100",
			2650 => "0000000111000000000101100100001000",
			2651 => "0000000110000000001001100100000100",
			2652 => "00000000000000000010101000001001",
			2653 => "00000000101100100010101000001001",
			2654 => "11111111000011000010101000001001",
			2655 => "0000000100000000000011101100001000",
			2656 => "0000000101000000000111111100000100",
			2657 => "00000000000000000010101000001001",
			2658 => "00000001001111110010101000001001",
			2659 => "0000001011000000001101000100000100",
			2660 => "11111111110000110010101000001001",
			2661 => "00000000000000000010101000001001",
			2662 => "0000000110000000001001111100000100",
			2663 => "11111110110011000010101000001001",
			2664 => "00000000000000000010101000001001",
			2665 => "0000000100000000001011110000010000",
			2666 => "0000000010000000001101101100001100",
			2667 => "0000000101000000001100100100001000",
			2668 => "0000000101000000001101000100000100",
			2669 => "00000000101100010010101000001001",
			2670 => "00000000000000000010101000001001",
			2671 => "00000001110100110010101000001001",
			2672 => "00000000000000000010101000001001",
			2673 => "0000001011000000000010001000000100",
			2674 => "11111111000101000010101000001001",
			2675 => "0000000000000000001101010000011000",
			2676 => "0000000000000000000010101000001000",
			2677 => "0000000100000000001011110000000100",
			2678 => "00000000000000000010101000001001",
			2679 => "11111111001111100010101000001001",
			2680 => "0000001101000000000010000100001000",
			2681 => "0000000000000000001101010000000100",
			2682 => "00000001001101110010101000001001",
			2683 => "00000000000000000010101000001001",
			2684 => "0000001100000000000001101000000100",
			2685 => "00000000000000000010101000001001",
			2686 => "11111111101110100010101000001001",
			2687 => "0000000010000000000011001100000100",
			2688 => "11111111001100110010101000001001",
			2689 => "00000000000000000010101000001001",
			2690 => "0000000001000000000101011100010100",
			2691 => "0000000000000000000111000000010000",
			2692 => "0000000011000000001000100000001100",
			2693 => "0000001100000000001011000000000100",
			2694 => "11111110011010110010101010110101",
			2695 => "0000001110000000000111111100000100",
			2696 => "00000011110011010010101010110101",
			2697 => "11111110011110110010101010110101",
			2698 => "00000100100110000010101010110101",
			2699 => "11111110011000010010101010110101",
			2700 => "0000001001000000000010101100111100",
			2701 => "0000000101000000001001010000100000",
			2702 => "0000000100000000001011110000011100",
			2703 => "0000001001000000001010100000001100",
			2704 => "0000000010000000001100000000001000",
			2705 => "0000000010000000001100010000000100",
			2706 => "11111110101101010010101010110101",
			2707 => "00000010001011000010101010110101",
			2708 => "11111110011101100010101010110101",
			2709 => "0000000010000000001111100100001000",
			2710 => "0000000110000000001001100100000100",
			2711 => "00000100001011000010101010110101",
			2712 => "00000010000000010010101010110101",
			2713 => "0000001011000000000010001000000100",
			2714 => "11111110001011010010101010110101",
			2715 => "00000011111100110010101010110101",
			2716 => "11111110010001100010101010110101",
			2717 => "0000001000000000000101000100001000",
			2718 => "0000001001000000000101010000000100",
			2719 => "00000000110011010010101010110101",
			2720 => "11111110011100100010101010110101",
			2721 => "0000000010000000000110111000001000",
			2722 => "0000000011000000001111101000000100",
			2723 => "00000110000001010010101010110101",
			2724 => "00000001001001100010101010110101",
			2725 => "0000001110000000001000101000000100",
			2726 => "11111110001111010010101010110101",
			2727 => "0000001011000000001110101000000100",
			2728 => "00000001101010110010101010110101",
			2729 => "11111111011100000010101010110101",
			2730 => "0000000001000000001100011000000100",
			2731 => "00000000011100000010101010110101",
			2732 => "11111110011010010010101010110101",
			2733 => "0000001011000000001010001100000100",
			2734 => "11111110011011110010101100100001",
			2735 => "0000001101000000001111100100110000",
			2736 => "0000001110000000000110001100100000",
			2737 => "0000000000000000000010011000011100",
			2738 => "0000001010000000000011101000001100",
			2739 => "0000001011000000000100000100001000",
			2740 => "0000000111000000000110100100000100",
			2741 => "00000000000000000010101100100001",
			2742 => "00000000111101000010101100100001",
			2743 => "11111110101011000010101100100001",
			2744 => "0000000110000000001001100100001000",
			2745 => "0000000010000000001000100000000100",
			2746 => "00000001110011010010101100100001",
			2747 => "11111111011010010010101100100001",
			2748 => "0000001100000000000100011000000100",
			2749 => "11111110110111110010101100100001",
			2750 => "00000000010101110010101100100001",
			2751 => "11111110101011110010101100100001",
			2752 => "0000001000000000000111000100001100",
			2753 => "0000000100000000001001001100000100",
			2754 => "00000000000000000010101100100001",
			2755 => "0000000001000000001010011000000100",
			2756 => "00000010000010110010101100100001",
			2757 => "00000000000000000010101100100001",
			2758 => "00000000000000000010101100100001",
			2759 => "11111110101010100010101100100001",
			2760 => "0000000000000000000001110100101100",
			2761 => "0000001110000000001011111000101000",
			2762 => "0000001010000000000011101000011000",
			2763 => "0000001011000000000111010000010000",
			2764 => "0000001011000000001010011100000100",
			2765 => "00000000000000000010101111110101",
			2766 => "0000000100000000001000001100001000",
			2767 => "0000000100000000000010000100000100",
			2768 => "00000000000000000010101111110101",
			2769 => "00000000100101110010101111110101",
			2770 => "00000000000000000010101111110101",
			2771 => "0000001011000000000100000100000100",
			2772 => "00000000000000000010101111110101",
			2773 => "11111111101100100010101111110101",
			2774 => "0000001110000000001110110100000100",
			2775 => "00000000000000000010101111110101",
			2776 => "0000001101000000001100100100000100",
			2777 => "00000000000000000010101111110101",
			2778 => "0000000100000000000010010100000100",
			2779 => "00000001001111000010101111110101",
			2780 => "00000000000000000010101111110101",
			2781 => "11111111011101010010101111110101",
			2782 => "0000001110000000001000101000010000",
			2783 => "0000001001000000000010101100001000",
			2784 => "0000000001000000001010011000000100",
			2785 => "11111110101010010010101111110101",
			2786 => "00000000000000000010101111110101",
			2787 => "0000000001000000001010011000000100",
			2788 => "00000000001010110010101111110101",
			2789 => "00000000000000000010101111110101",
			2790 => "0000000000000000000111000000001000",
			2791 => "0000000010000000001110000000000100",
			2792 => "11111110111001010010101111110101",
			2793 => "00000000000000000010101111110101",
			2794 => "0000000010000000001110000000001100",
			2795 => "0000001101000000001010001000000100",
			2796 => "00000000000000000010101111110101",
			2797 => "0000001101000000001001100000000100",
			2798 => "00000001000100010010101111110101",
			2799 => "00000000000000000010101111110101",
			2800 => "0000001011000000000010110100010000",
			2801 => "0000001100000000001000011000001000",
			2802 => "0000001101000000000010000100000100",
			2803 => "11111111110010100010101111110101",
			2804 => "00000000000000000010101111110101",
			2805 => "0000000110000000001000010000000100",
			2806 => "00000000000000000010101111110101",
			2807 => "00000000011001000010101111110101",
			2808 => "0000001100000000001111011100000100",
			2809 => "00000000000000000010101111110101",
			2810 => "0000001111000000001001001100000100",
			2811 => "11111111001010100010101111110101",
			2812 => "00000000000000000010101111110101",
			2813 => "0000000001000000000101011100010100",
			2814 => "0000000000000000000111000100010000",
			2815 => "0000000011000000001000100000001100",
			2816 => "0000000001000000001101101000001000",
			2817 => "0000000111000000000100001000000100",
			2818 => "11111110100010000010110010011001",
			2819 => "00000011110110000010110010011001",
			2820 => "11111110011011000010110010011001",
			2821 => "00000100010001010010110010011001",
			2822 => "11111110011000110010110010011001",
			2823 => "0000000001000000001010011000111100",
			2824 => "0000000101000000001001010000011100",
			2825 => "0000000100000000001011110000011000",
			2826 => "0000000001000000001101111100001100",
			2827 => "0000000010000000001100000000001000",
			2828 => "0000000010000000001100010000000100",
			2829 => "11111110110000100010110010011001",
			2830 => "00000010000000100010110010011001",
			2831 => "11111110011110110010110010011001",
			2832 => "0000000011000000001100111000001000",
			2833 => "0000000000000000001010101100000100",
			2834 => "00000010101000110010110010011001",
			2835 => "11111110111100110010110010011001",
			2836 => "11111110000100100010110010011001",
			2837 => "11111110010010100010110010011001",
			2838 => "0000001000000000000101000100001000",
			2839 => "0000000001000000000001000100000100",
			2840 => "00000000011011110010110010011001",
			2841 => "11111110011100010010110010011001",
			2842 => "0000001101000000000111010100001100",
			2843 => "0000000010000000001111101000000100",
			2844 => "00000101000000100010110010011001",
			2845 => "0000001010000000001000010100000100",
			2846 => "11111110111100100010110010011001",
			2847 => "00000001100011100010110010011001",
			2848 => "0000000110000000001001111100000100",
			2849 => "11111011101011000010110010011001",
			2850 => "0000001000000000001011010100000100",
			2851 => "00000000110010110010110010011001",
			2852 => "00000010110111100010110010011001",
			2853 => "11111110011010110010110010011001",
			2854 => "0000001001000000001000010000011100",
			2855 => "0000000000000000000111000000011000",
			2856 => "0000000000000000000001010100000100",
			2857 => "11111110011001000010110101010101",
			2858 => "0000000000000000000001010100000100",
			2859 => "00000000010010000010110101010101",
			2860 => "0000000000000000000111000000001100",
			2861 => "0000000000000000000110001000000100",
			2862 => "11111110011101100010110101010101",
			2863 => "0000000000000000001111001000000100",
			2864 => "00000101100010100010110101010101",
			2865 => "11111110011111100010110101010101",
			2866 => "00000000000000000010110101010101",
			2867 => "11111110011000000010110101010101",
			2868 => "0000001001000000000010101100111100",
			2869 => "0000001101000000001110010000011100",
			2870 => "0000001001000000001010100100010100",
			2871 => "0000000010000000001100000000001000",
			2872 => "0000001010000000000011101000000100",
			2873 => "11111110011111000010110101010101",
			2874 => "00010111010110110010110101010101",
			2875 => "0000000100000000000010010100001000",
			2876 => "0000000000000000000111000100000100",
			2877 => "11111110011010100010110101010101",
			2878 => "00000101110001100010110101010101",
			2879 => "11111110010100110010110101010101",
			2880 => "0000001010000000001000010100000100",
			2881 => "00000100100000100010110101010101",
			2882 => "11111110011001110010110101010101",
			2883 => "0000000110000000000100111100001100",
			2884 => "0000000101000000000010011100000100",
			2885 => "00000011100101000010110101010101",
			2886 => "0000000000000000000111000000000100",
			2887 => "11111110011001000010110101010101",
			2888 => "11111100101100100010110101010101",
			2889 => "0000000010000000001110000000000100",
			2890 => "00001011000110110010110101010101",
			2891 => "0000001001000000001010100000001000",
			2892 => "0000001101000000000111010100000100",
			2893 => "00000010001001110010110101010101",
			2894 => "00000000001110010010110101010101",
			2895 => "0000000100000000001110111000000100",
			2896 => "00000110010001110010110101010101",
			2897 => "00000001001110000010110101010101",
			2898 => "0000000011000000000001011100000100",
			2899 => "00000100001110010010110101010101",
			2900 => "11111110011000010010110101010101",
			2901 => "0000001100000000001010111000001000",
			2902 => "0000000001000000001100011000000100",
			2903 => "11111110100110000010111000010001",
			2904 => "00000000000000000010111000010001",
			2905 => "0000000100000000000011001100111100",
			2906 => "0000001000000000000101000100100000",
			2907 => "0000000101000000001110101100001100",
			2908 => "0000000100000000000110101100001000",
			2909 => "0000000010000000001010001000000100",
			2910 => "00000000000000000010111000010001",
			2911 => "00000001000011010010111000010001",
			2912 => "00000000000000000010111000010001",
			2913 => "0000001101000000000011001000001100",
			2914 => "0000001001000000001010100100001000",
			2915 => "0000001011000000000100000100000100",
			2916 => "00000000000000000010111000010001",
			2917 => "11111110111100000010111000010001",
			2918 => "00000000000000000010111000010001",
			2919 => "0000001011000000001011110100000100",
			2920 => "00000000010010000010111000010001",
			2921 => "00000000000000000010111000010001",
			2922 => "0000001101000000000110010000010000",
			2923 => "0000001011000000001011011100000100",
			2924 => "11111111111110000010111000010001",
			2925 => "0000001000000000001100000100001000",
			2926 => "0000001100000000000100011000000100",
			2927 => "00000000000000000010111000010001",
			2928 => "00000001010101010010111000010001",
			2929 => "00000000000000000010111000010001",
			2930 => "0000000110000000001000010000000100",
			2931 => "11111111000100110010111000010001",
			2932 => "0000000001000000001100011000000100",
			2933 => "00000000110100100010111000010001",
			2934 => "00000000000000000010111000010001",
			2935 => "0000001110000000001000000100000100",
			2936 => "11111110110001100010111000010001",
			2937 => "0000000101000000001100010000010000",
			2938 => "0000001101000000001001100000000100",
			2939 => "11111111111100010010111000010001",
			2940 => "0000000001000000001100011000001000",
			2941 => "0000000001000000001011111100000100",
			2942 => "00000000000000000010111000010001",
			2943 => "00000001001011010010111000010001",
			2944 => "00000000000000000010111000010001",
			2945 => "0000000110000000001001111100000100",
			2946 => "11111110111111110010111000010001",
			2947 => "00000000000000000010111000010001",
			2948 => "0000001100000000001101010100000100",
			2949 => "11111110101101110010111010100101",
			2950 => "0000001100000000000001011000111100",
			2951 => "0000000111000000000001101000010100",
			2952 => "0000000000000000000010101000010000",
			2953 => "0000001001000000000000001000000100",
			2954 => "00000000000000000010111010100101",
			2955 => "0000001100000000001000000000001000",
			2956 => "0000000100000000001011110000000100",
			2957 => "00000001001110100010111010100101",
			2958 => "00000000000000000010111010100101",
			2959 => "00000000000000000010111010100101",
			2960 => "11111111100101000010111010100101",
			2961 => "0000001110000000001000110100011000",
			2962 => "0000000100000000000011001100010000",
			2963 => "0000000000000000000111000000001000",
			2964 => "0000000001000000001001011000000100",
			2965 => "00000000000000000010111010100101",
			2966 => "11111111011101010010111010100101",
			2967 => "0000001011000000001011110100000100",
			2968 => "11111111111110100010111010100101",
			2969 => "00000000110010000010111010100101",
			2970 => "0000001110000000001000000100000100",
			2971 => "11111110111100000010111010100101",
			2972 => "00000000000000000010111010100101",
			2973 => "0000001011000000000000110100000100",
			2974 => "00000000000000000010111010100101",
			2975 => "0000001001000000000010101100001000",
			2976 => "0000000000000000000100000000000100",
			2977 => "00000001010011010010111010100101",
			2978 => "00000000000000000010111010100101",
			2979 => "00000000000000000010111010100101",
			2980 => "0000000111000000000100010000000100",
			2981 => "00000000000000000010111010100101",
			2982 => "0000000110000000001001111100000100",
			2983 => "11111110110011100010111010100101",
			2984 => "00000000000000000010111010100101",
			2985 => "0000000001000000001101011100000100",
			2986 => "11111110011001110010111100100001",
			2987 => "0000001001000000000010101100110100",
			2988 => "0000000000000000001011010100000100",
			2989 => "11111110100000010010111100100001",
			2990 => "0000000100000000001011110000011000",
			2991 => "0000000101000000001100100100001100",
			2992 => "0000000100000000001111100100000100",
			2993 => "00000010101110110010111100100001",
			2994 => "0000000001000000000100110100000100",
			2995 => "11111110100110100010111100100001",
			2996 => "00000000000101100010111100100001",
			2997 => "0000001110000000001011101100001000",
			2998 => "0000000000000000000110001000000100",
			2999 => "00000000000000000010111100100001",
			3000 => "00000100011111000010111100100001",
			3001 => "11111111010000110010111100100001",
			3002 => "0000001110000000001100001100001100",
			3003 => "0000000100000000001001001100001000",
			3004 => "0000001011000000000010001000000100",
			3005 => "11111110011111000010111100100001",
			3006 => "00000000110111010010111100100001",
			3007 => "11111101110010000010111100100001",
			3008 => "0000001000000000001001101000000100",
			3009 => "11111111010001000010111100100001",
			3010 => "0000001001000000001010100000000100",
			3011 => "00000001010100110010111100100001",
			3012 => "00000011000100100010111100100001",
			3013 => "0000000100000000001011110000000100",
			3014 => "00000000101100000010111100100001",
			3015 => "11111110011110100010111100100001",
			3016 => "0000001100000000001101010100000100",
			3017 => "11111110100001100010111111101101",
			3018 => "0000001001000000001010100000101100",
			3019 => "0000001110000000001000011100011000",
			3020 => "0000001001000000000101010000010000",
			3021 => "0000000100000000000011110000001100",
			3022 => "0000000110000000000100110100000100",
			3023 => "00000000000000000010111111101101",
			3024 => "0000001100000000000100011000000100",
			3025 => "00000000000000000010111111101101",
			3026 => "00000000101111010010111111101101",
			3027 => "11111111101110010010111111101101",
			3028 => "0000001110000000001011110000000100",
			3029 => "11111110110110100010111111101101",
			3030 => "00000000000000000010111111101101",
			3031 => "0000000011000000001110111000001100",
			3032 => "0000000011000000001110100100000100",
			3033 => "00000000000000000010111111101101",
			3034 => "0000000000000000001011000100000100",
			3035 => "00000001000010010010111111101101",
			3036 => "00000000000000000010111111101101",
			3037 => "0000000101000000001100000000000100",
			3038 => "00000000000000000010111111101101",
			3039 => "11111111110010000010111111101101",
			3040 => "0000001100000000001000000000010100",
			3041 => "0000001001000000001010100100001000",
			3042 => "0000000110000000001111000000000100",
			3043 => "00000000101101110010111111101101",
			3044 => "11111111000001000010111111101101",
			3045 => "0000000000000000001000101100001000",
			3046 => "0000001011000000001011011100000100",
			3047 => "00000000000000000010111111101101",
			3048 => "00000001101100000010111111101101",
			3049 => "11111111111001000010111111101101",
			3050 => "0000001000000000000001110000001100",
			3051 => "0000001001000000001010100100001000",
			3052 => "0000001001000000001010100100000100",
			3053 => "11111111000110110010111111101101",
			3054 => "00000000100111000010111111101101",
			3055 => "11111110101000010010111111101101",
			3056 => "0000000101000000000011001000001100",
			3057 => "0000001000000000001100000100001000",
			3058 => "0000001001000000001010100100000100",
			3059 => "00000000101001100010111111101101",
			3060 => "00000000000000000010111111101101",
			3061 => "11111111010000010010111111101101",
			3062 => "0000001110000000001110000000000100",
			3063 => "00000000000000000010111111101101",
			3064 => "0000001001000000000010101100000100",
			3065 => "00000001011110110010111111101101",
			3066 => "00000000000000000010111111101101",
			3067 => "0000000101000000000001001000000100",
			3068 => "11111110011100010011000010000001",
			3069 => "0000000011000000001100111000100000",
			3070 => "0000001010000000000011101000001000",
			3071 => "0000000001000000001111001100000100",
			3072 => "00000001001110100011000010000001",
			3073 => "11111110110000100011000010000001",
			3074 => "0000000000000000000010101000010100",
			3075 => "0000000101000000001100100100001100",
			3076 => "0000000100000000001111100100000100",
			3077 => "00000001110110000011000010000001",
			3078 => "0000001001000000001010100100000100",
			3079 => "11111110101101110011000010000001",
			3080 => "00000000111110000011000010000001",
			3081 => "0000000100000000000001011100000100",
			3082 => "00000000000000000011000010000001",
			3083 => "00000001111000100011000010000001",
			3084 => "11111111001100010011000010000001",
			3085 => "0000000000000000000010101000000100",
			3086 => "11111110010010100011000010000001",
			3087 => "0000001011000000000010001000000100",
			3088 => "11111110100111000011000010000001",
			3089 => "0000001100000000001000011000010000",
			3090 => "0000000001000000001100011000001000",
			3091 => "0000000101000000001001010000000100",
			3092 => "11111110101100000011000010000001",
			3093 => "00000000101110010011000010000001",
			3094 => "0000001000000000001001101000000100",
			3095 => "00000001111100110011000010000001",
			3096 => "00000000000000000011000010000001",
			3097 => "0000001010000000001001000100001000",
			3098 => "0000000111000000000000011100000100",
			3099 => "00000000000000000011000010000001",
			3100 => "11111110101001000011000010000001",
			3101 => "0000001101000000001111100100000100",
			3102 => "00000000011100000011000010000001",
			3103 => "11111110100111110011000010000001",
			3104 => "0000000001000000001101111101001000",
			3105 => "0000001100000000000100011000001000",
			3106 => "0000000011000000000010010100000100",
			3107 => "11111110011101010011000110001101",
			3108 => "00000000000000000011000110001101",
			3109 => "0000000000000000000111000000011100",
			3110 => "0000000110000000001001100100001100",
			3111 => "0000000010000000001010001000001000",
			3112 => "0000001101000000000001000000000100",
			3113 => "00000000000100000011000110001101",
			3114 => "00000000000000000011000110001101",
			3115 => "11111111000001000011000110001101",
			3116 => "0000001011000000000110110100000100",
			3117 => "00000000000000000011000110001101",
			3118 => "0000000101000000000111111100001000",
			3119 => "0000000001000000000001111000000100",
			3120 => "00000001100011100011000110001101",
			3121 => "00000000000000000011000110001101",
			3122 => "00000000000000000011000110001101",
			3123 => "0000001110000000001000011100010000",
			3124 => "0000001001000000001001111100001100",
			3125 => "0000001001000000001000010000000100",
			3126 => "11111110111111100011000110001101",
			3127 => "0000001001000000000101010000000100",
			3128 => "00000000010101110011000110001101",
			3129 => "00000000000000000011000110001101",
			3130 => "11111110100010100011000110001101",
			3131 => "0000001011000000000111100000001100",
			3132 => "0000000011000000001110100100000100",
			3133 => "00000000000000000011000110001101",
			3134 => "0000000000000000001100001000000100",
			3135 => "00000001001100000011000110001101",
			3136 => "00000000000000000011000110001101",
			3137 => "0000001101000000001111100100000100",
			3138 => "00000000000000000011000110001101",
			3139 => "11111111011101100011000110001101",
			3140 => "0000001100000000001000011000110100",
			3141 => "0000001101000000000111111100010000",
			3142 => "0000000011000000001111100100001100",
			3143 => "0000001001000000001010100000000100",
			3144 => "11111111110100100011000110001101",
			3145 => "0000000000000000000001110100000100",
			3146 => "00000001010110000011000110001101",
			3147 => "00000000000000000011000110001101",
			3148 => "11111110101111100011000110001101",
			3149 => "0000000101000000001110000100001000",
			3150 => "0000001001000000001010100100000100",
			3151 => "00000000000000000011000110001101",
			3152 => "00000010110010100011000110001101",
			3153 => "0000000000000000000111000000001100",
			3154 => "0000000011000000000001011100001000",
			3155 => "0000001010000000001000100100000100",
			3156 => "00000000000000000011000110001101",
			3157 => "00000001010001000011000110001101",
			3158 => "11111110100011100011000110001101",
			3159 => "0000001000000000001001101000001000",
			3160 => "0000000101000000001001010000000100",
			3161 => "00000000000000000011000110001101",
			3162 => "00000001110100100011000110001101",
			3163 => "0000000010000000000011001100000100",
			3164 => "11111111111100010011000110001101",
			3165 => "00000000000000000011000110001101",
			3166 => "0000000001000000000100110100000100",
			3167 => "00000000101100010011000110001101",
			3168 => "0000001110000000000010111000000100",
			3169 => "11111110110000110011000110001101",
			3170 => "00000000000000000011000110001101",
			3171 => "0000001100000000001101010100000100",
			3172 => "11111110011101000011001001001001",
			3173 => "0000001001000000001010100101001000",
			3174 => "0000001011000000000111010000010100",
			3175 => "0000000000000000000110001000010000",
			3176 => "0000000110000000000100110100000100",
			3177 => "00000000000000000011001001001001",
			3178 => "0000000100000000001111100100001000",
			3179 => "0000000111000000000011100000000100",
			3180 => "00000000000000000011001001001001",
			3181 => "00000001110000100011001001001001",
			3182 => "00000000000000000011001001001001",
			3183 => "11111111110110100011001001001001",
			3184 => "0000001011000000000110110100011000",
			3185 => "0000001011000000000100000100001100",
			3186 => "0000000100000000001111100100001000",
			3187 => "0000001001000000000111101100000100",
			3188 => "00000000000000000011001001001001",
			3189 => "00000000011011000011001001001001",
			3190 => "00000000000000000011001001001001",
			3191 => "0000000101000000001100100100000100",
			3192 => "11111110101011110011001001001001",
			3193 => "0000000101000000000111100000000100",
			3194 => "00000000000000000011001001001001",
			3195 => "11111111010101100011001001001001",
			3196 => "0000000000000000001000101100001100",
			3197 => "0000000110000000001001100100000100",
			3198 => "11111111010000010011001001001001",
			3199 => "0000000001000000000001111000000100",
			3200 => "00000001100010110011001001001001",
			3201 => "00000000010010010011001001001001",
			3202 => "0000001110000000001011110000001000",
			3203 => "0000000000000000001000110000000100",
			3204 => "00000000000000000011001001001001",
			3205 => "11111110010110010011001001001001",
			3206 => "0000001101000000001111100100000100",
			3207 => "00000000111100110011001001001001",
			3208 => "11111110110010100011001001001001",
			3209 => "0000001100000000001000000000010000",
			3210 => "0000001100000000001011000000001000",
			3211 => "0000001011000000000101100100000100",
			3212 => "00000000000000000011001001001001",
			3213 => "11111111010010010011001001001001",
			3214 => "0000000000000000001101010000000100",
			3215 => "00000001010111100011001001001001",
			3216 => "00000000000000000011001001001001",
			3217 => "11111110011000010011001001001001",
			3218 => "0000001100000000001010111000001000",
			3219 => "0000000001000000001100011000000100",
			3220 => "11111110011011000011001011110101",
			3221 => "00000000000000000011001011110101",
			3222 => "0000001101000000001111100101001100",
			3223 => "0000001110000000000101000000111100",
			3224 => "0000000010000000001110000000100000",
			3225 => "0000000000000000000111000000010000",
			3226 => "0000001110000000001101101100001000",
			3227 => "0000000100000000001111101000000100",
			3228 => "00000000000000100011001011110101",
			3229 => "00000001011011000011001011110101",
			3230 => "0000000001000000001101111100000100",
			3231 => "00000000001111010011001011110101",
			3232 => "11111101111001100011001011110101",
			3233 => "0000001001000000001010100100001000",
			3234 => "0000000111000000000111010000000100",
			3235 => "11111110101000010011001011110101",
			3236 => "00000000110010000011001011110101",
			3237 => "0000001100000000000001101000000100",
			3238 => "00000010000100110011001011110101",
			3239 => "11111111111000110011001011110101",
			3240 => "0000001110000000001011110000010000",
			3241 => "0000000010000000001000110100001000",
			3242 => "0000000001000000000111101000000100",
			3243 => "00000000010111100011001011110101",
			3244 => "11111111010001010011001011110101",
			3245 => "0000001010000000001001000100000100",
			3246 => "00000000000000000011001011110101",
			3247 => "11111110001100010011001011110101",
			3248 => "0000001000000000001100000100000100",
			3249 => "11111110101110000011001011110101",
			3250 => "0000001000000000001001101000000100",
			3251 => "00000001000001100011001011110101",
			3252 => "11111110110111110011001011110101",
			3253 => "0000000001000000001100011000001100",
			3254 => "0000000000000000001011000100001000",
			3255 => "0000000101000000000011001000000100",
			3256 => "00000000000000000011001011110101",
			3257 => "00000001101011110011001011110101",
			3258 => "00000000000000000011001011110101",
			3259 => "11111111011011010011001011110101",
			3260 => "11111110011000110011001011110101",
			3261 => "0000001110000000001110110100000100",
			3262 => "11111110011010000011001110010011",
			3263 => "0000001101000000001111100101001000",
			3264 => "0000001110000000001100001100110100",
			3265 => "0000000111000000000101100100011100",
			3266 => "0000001000000000001100000100001100",
			3267 => "0000000110000000001011001100000100",
			3268 => "11111110101001000011001110010011",
			3269 => "0000000110000000001111000000000100",
			3270 => "00000010110101010011001110010011",
			3271 => "00000001001101100011001110010011",
			3272 => "0000001101000000001001100000001000",
			3273 => "0000001011000000001010010100000100",
			3274 => "11111110001010010011001110010011",
			3275 => "11111111011110100011001110010011",
			3276 => "0000000100000000001010110100000100",
			3277 => "00000010000000100011001110010011",
			3278 => "00000000000000000011001110010011",
			3279 => "0000001110000000001000011100001100",
			3280 => "0000000100000000001101001000001000",
			3281 => "0000001000000000000001110000000100",
			3282 => "11111110100010110011001110010011",
			3283 => "00000000110010110011001110010011",
			3284 => "11111101111011010011001110010011",
			3285 => "0000000000000000001000110000000100",
			3286 => "11111111000101110011001110010011",
			3287 => "0000000000000000000010011000000100",
			3288 => "00000001011100010011001110010011",
			3289 => "00000000000000000011001110010011",
			3290 => "0000001000000000000111000100010000",
			3291 => "0000000101000000000011001000000100",
			3292 => "11111111101110100011001110010011",
			3293 => "0000000111000000000101100100000100",
			3294 => "00000101100011000011001110010011",
			3295 => "0000001000000000001100000100000100",
			3296 => "11111111111100100011001110010011",
			3297 => "00000001110001000011001110010011",
			3298 => "11111111010001100011001110010011",
			3299 => "11111110010010010011001110010011",
			3300 => "00000000000000000011001110010101",
			3301 => "00000000000000000011001110011001",
			3302 => "00000000000000000011001110011101",
			3303 => "00000000000000000011001110100001",
			3304 => "00000000000000000011001110100101",
			3305 => "00000000000000000011001110101001",
			3306 => "00000000000000000011001110101101",
			3307 => "00000000000000000011001110110001",
			3308 => "00000000000000000011001110110101",
			3309 => "00000000000000000011001110111001",
			3310 => "00000000000000000011001110111101",
			3311 => "00000000000000000011001111000001",
			3312 => "00000000000000000011001111000101",
			3313 => "00000000000000000011001111001001",
			3314 => "00000000000000000011001111001101",
			3315 => "00000000000000000011001111010001",
			3316 => "00000000000000000011001111010101",
			3317 => "00000000000000000011001111011001",
			3318 => "00000000000000000011001111011101",
			3319 => "0000001001000000001010100100000100",
			3320 => "11111111111111000011001111101001",
			3321 => "00000000000000000011001111101001",
			3322 => "0000000110000000000100111100000100",
			3323 => "00000000000000000011001111111101",
			3324 => "0000000110000000001001111100000100",
			3325 => "00000000000100110011001111111101",
			3326 => "00000000000000000011001111111101",
			3327 => "0000000001000000000100110100001000",
			3328 => "0000000001000000000111101000000100",
			3329 => "00000000000000000011010000010001",
			3330 => "00000000010100010011010000010001",
			3331 => "00000000000000000011010000010001",
			3332 => "0000000001000000001100011000001000",
			3333 => "0000000000000000000001110000000100",
			3334 => "00000000000000000011010000100101",
			3335 => "11111111111001100011010000100101",
			3336 => "00000000000000000011010000100101",
			3337 => "0000001001000000001010100100001000",
			3338 => "0000000110000000001001111100000100",
			3339 => "11111111110011000011010000111001",
			3340 => "00000000000000000011010000111001",
			3341 => "00000000000000000011010000111001",
			3342 => "0000000111000000001111011100001000",
			3343 => "0000000111000000000001101000000100",
			3344 => "00000000000000000011010001010101",
			3345 => "11111111111010100011010001010101",
			3346 => "0000000111000000000100010000000100",
			3347 => "00000000001101100011010001010101",
			3348 => "00000000000000000011010001010101",
			3349 => "0000000000000000000010101000001100",
			3350 => "0000001000000000001010110000000100",
			3351 => "00000000000000000011010001110001",
			3352 => "0000001000000000000001010100000100",
			3353 => "00000000000111100011010001110001",
			3354 => "00000000000000000011010001110001",
			3355 => "11111111111101100011010001110001",
			3356 => "0000000100000000001000011100000100",
			3357 => "00000000000000000011010010001101",
			3358 => "0000000010000000000011110100001000",
			3359 => "0000000001000000000111101000000100",
			3360 => "00000000000000000011010010001101",
			3361 => "11111111110011000011010010001101",
			3362 => "00000000000000000011010010001101",
			3363 => "0000001001000000001010100000000100",
			3364 => "00000000000000000011010010101001",
			3365 => "0000000101000000000111011000001000",
			3366 => "0000001001000000000011101000000100",
			3367 => "00000000010011010011010010101001",
			3368 => "00000000000000000011010010101001",
			3369 => "00000000000000000011010010101001",
			3370 => "0000000000000000000010101000001100",
			3371 => "0000001001000000001010100100000100",
			3372 => "00000000000000000011010011010101",
			3373 => "0000001111000000000011000000000100",
			3374 => "00000000011000010011010011010101",
			3375 => "00000000000000000011010011010101",
			3376 => "0000000011000000001000110100001000",
			3377 => "0000000000000000001010101100000100",
			3378 => "00000000000000000011010011010101",
			3379 => "11111111101111100011010011010101",
			3380 => "00000000000000000011010011010101",
			3381 => "0000001011000000001011011100000100",
			3382 => "00000000000000000011010011111001",
			3383 => "0000000110000000001001111100001100",
			3384 => "0000000110000000000100111100000100",
			3385 => "00000000000000000011010011111001",
			3386 => "0000001011000000000110100000000100",
			3387 => "00000000001101010011010011111001",
			3388 => "00000000000000000011010011111001",
			3389 => "00000000000000000011010011111001",
			3390 => "0000001001000000001010100000000100",
			3391 => "00000000000000000011010100011101",
			3392 => "0000001011000000000010110100001100",
			3393 => "0000001001000000000011101000001000",
			3394 => "0000001001000000001010100000000100",
			3395 => "00000000000000000011010100011101",
			3396 => "00000000001011000011010100011101",
			3397 => "00000000000000000011010100011101",
			3398 => "00000000000000000011010100011101",
			3399 => "0000000000000000001000101100010000",
			3400 => "0000001010000000000011101000000100",
			3401 => "00000000000000000011010101001001",
			3402 => "0000000101000000000011001000001000",
			3403 => "0000000101000000001100100100000100",
			3404 => "00000000000000000011010101001001",
			3405 => "00000000010001000011010101001001",
			3406 => "00000000000000000011010101001001",
			3407 => "0000000010000000000011110100000100",
			3408 => "11111111111101010011010101001001",
			3409 => "00000000000000000011010101001001",
			3410 => "0000001001000000000111101100000100",
			3411 => "00000000000000000011010101110101",
			3412 => "0000000001000000000100110100001000",
			3413 => "0000001000000000001010110000000100",
			3414 => "00000000000000000011010101110101",
			3415 => "00000000001101100011010101110101",
			3416 => "0000000011000000001011101100000100",
			3417 => "00000000000000000011010101110101",
			3418 => "0000000011000000000011110000000100",
			3419 => "11111111110110110011010101110101",
			3420 => "00000000000000000011010101110101",
			3421 => "0000001001000000001010100100010100",
			3422 => "0000000111000000000111010000001000",
			3423 => "0000000100000000001111100100000100",
			3424 => "00000000000000000011010110110001",
			3425 => "11111111011011000011010110110001",
			3426 => "0000000111000000000100010000001000",
			3427 => "0000001011000000001011110100000100",
			3428 => "00000000000000000011010110110001",
			3429 => "00000000001000000011010110110001",
			3430 => "00000000000000000011010110110001",
			3431 => "0000000111000000001111011100001000",
			3432 => "0000001001000000000011101000000100",
			3433 => "00000000001100110011010110110001",
			3434 => "00000000000000000011010110110001",
			3435 => "00000000000000000011010110110001",
			3436 => "0000000000000000001101010000010100",
			3437 => "0000001010000000000011101000000100",
			3438 => "00000000000000000011010111011101",
			3439 => "0000001001000000001010100100001100",
			3440 => "0000001001000000001010011000000100",
			3441 => "00000000000000000011010111011101",
			3442 => "0000000000000000001011010100000100",
			3443 => "00000000000000000011010111011101",
			3444 => "00000000000100010011010111011101",
			3445 => "00000000000000000011010111011101",
			3446 => "11111111111100100011010111011101",
			3447 => "0000001000000000000001010100001100",
			3448 => "0000001001000000001010100100000100",
			3449 => "00000000000000000011011000100001",
			3450 => "0000000010000000000001011100000100",
			3451 => "00000000011110000011011000100001",
			3452 => "00000000000000000011011000100001",
			3453 => "0000001110000000001110000000001100",
			3454 => "0000000001000000001100011000001000",
			3455 => "0000000100000000000110111000000100",
			3456 => "00000000000000000011011000100001",
			3457 => "11111111100111110011011000100001",
			3458 => "00000000000000000011011000100001",
			3459 => "0000001101000000001111100100001000",
			3460 => "0000000111000000000111010000000100",
			3461 => "00000000000000000011011000100001",
			3462 => "00000000010001110011011000100001",
			3463 => "00000000000000000011011000100001",
			3464 => "0000001000000000000001010100010000",
			3465 => "0000000101000000001100100100000100",
			3466 => "00000000000000000011011001100101",
			3467 => "0000000000000000001111001000000100",
			3468 => "00000000000000000011011001100101",
			3469 => "0000000101000000000010011100000100",
			3470 => "00000000010111000011011001100101",
			3471 => "00000000000000000011011001100101",
			3472 => "0000001110000000001110000000010000",
			3473 => "0000000001000000001100011000001100",
			3474 => "0000000100000000001000110100000100",
			3475 => "00000000000000000011011001100101",
			3476 => "0000001001000000001001111100000100",
			3477 => "00000000000000000011011001100101",
			3478 => "11111111100001010011011001100101",
			3479 => "00000000000000000011011001100101",
			3480 => "00000000000000000011011001100101",
			3481 => "0000001001000000000111101100010000",
			3482 => "0000000111000000000111010000001100",
			3483 => "0000001110000000001000101000001000",
			3484 => "0000000110000000000100110100000100",
			3485 => "00000000000000000011011010111001",
			3486 => "11111111110100010011011010111001",
			3487 => "00000000000000000011011010111001",
			3488 => "00000000000000000011011010111001",
			3489 => "0000000001000000000100110100001100",
			3490 => "0000001010000000000011101000000100",
			3491 => "00000000000000000011011010111001",
			3492 => "0000001110000000000110010000000100",
			3493 => "00000000000000000011011010111001",
			3494 => "00000000010010110011011010111001",
			3495 => "0000000011000000001011101100000100",
			3496 => "00000000000000000011011010111001",
			3497 => "0000000011000000000011110000001000",
			3498 => "0000001100000000001000000000000100",
			3499 => "00000000000000000011011010111001",
			3500 => "11111111101110110011011010111001",
			3501 => "00000000000000000011011010111001",
			3502 => "0000000100000000001011110000011000",
			3503 => "0000001110000000001011101100010100",
			3504 => "0000001101000000001110101100000100",
			3505 => "00000000000000000011011011110101",
			3506 => "0000001000000000001000100100000100",
			3507 => "00000000000000000011011011110101",
			3508 => "0000001101000000001100010100001000",
			3509 => "0000000000000000001010101100000100",
			3510 => "00000000010110000011011011110101",
			3511 => "00000000000000000011011011110101",
			3512 => "00000000000000000011011011110101",
			3513 => "00000000000000000011011011110101",
			3514 => "0000001110000000000010010100000100",
			3515 => "11111111110011100011011011110101",
			3516 => "00000000000000000011011011110101",
			3517 => "0000001011000000000101110100011000",
			3518 => "0000001000000000000001110000010100",
			3519 => "0000001011000000001011011100000100",
			3520 => "00000000000000000011011101000001",
			3521 => "0000001111000000001111100100000100",
			3522 => "00000000000000000011011101000001",
			3523 => "0000001100000000000100011000000100",
			3524 => "00000000000000000011011101000001",
			3525 => "0000000100000000001000101000000100",
			3526 => "00000000000000000011011101000001",
			3527 => "00000000100011000011011101000001",
			3528 => "00000000000000000011011101000001",
			3529 => "0000001000000000000001110000001000",
			3530 => "0000001110000000000110111100000100",
			3531 => "00000000000000000011011101000001",
			3532 => "11111111110010100011011101000001",
			3533 => "0000001000000000001011010100000100",
			3534 => "00000000000101010011011101000001",
			3535 => "00000000000000000011011101000001",
			3536 => "0000000101000000001001010000000100",
			3537 => "00000000000000000011011101110101",
			3538 => "0000001101000000001011111000010100",
			3539 => "0000001001000000000010101100010000",
			3540 => "0000000000000000000010101000000100",
			3541 => "00000000000000000011011101110101",
			3542 => "0000001110000000001100111000000100",
			3543 => "00000000000000000011011101110101",
			3544 => "0000001000000000000111000100000100",
			3545 => "00000000011100100011011101110101",
			3546 => "00000000000000000011011101110101",
			3547 => "00000000000000000011011101110101",
			3548 => "00000000000000000011011101110101",
			3549 => "0000001001000000001010100000000100",
			3550 => "00000000000000000011011110101001",
			3551 => "0000000111000000000101100100010100",
			3552 => "0000000100000000001001001100010000",
			3553 => "0000001001000000001010100000000100",
			3554 => "00000000000000000011011110101001",
			3555 => "0000001001000000000011101000001000",
			3556 => "0000000101000000001100010100000100",
			3557 => "00000000010001000011011110101001",
			3558 => "00000000000000000011011110101001",
			3559 => "00000000000000000011011110101001",
			3560 => "00000000000000000011011110101001",
			3561 => "00000000000000000011011110101001",
			3562 => "0000000100000000001011110000011000",
			3563 => "0000000011000000001101101100010100",
			3564 => "0000001000000000001010110000000100",
			3565 => "00000000000000000011011111110101",
			3566 => "0000001000000000000001010100001100",
			3567 => "0000001011000000001011011100000100",
			3568 => "00000000000000000011011111110101",
			3569 => "0000000011000000001000001100000100",
			3570 => "00000000000000000011011111110101",
			3571 => "00000000010101110011011111110101",
			3572 => "00000000000000000011011111110101",
			3573 => "00000000000000000011011111110101",
			3574 => "0000000011000000001000000100000100",
			3575 => "11111111111010110011011111110101",
			3576 => "0000001011000000001001010000001000",
			3577 => "0000001011000000001011110100000100",
			3578 => "00000000000000000011011111110101",
			3579 => "00000000000100000011011111110101",
			3580 => "00000000000000000011011111110101",
			3581 => "0000001000000000000110011100010100",
			3582 => "0000001010000000000011101000000100",
			3583 => "00000000000000000011100001011001",
			3584 => "0000001010000000000111110100001100",
			3585 => "0000000110000000001111000000001000",
			3586 => "0000000110000000001011001100000100",
			3587 => "00000000000000000011100001011001",
			3588 => "00000000001000100011100001011001",
			3589 => "00000000000000000011100001011001",
			3590 => "00000000000000000011100001011001",
			3591 => "0000000110000000001000010000001000",
			3592 => "0000000001000000001100011000000100",
			3593 => "11111111001100110011100001011001",
			3594 => "00000000000000000011100001011001",
			3595 => "0000000000000000001101010000001100",
			3596 => "0000000010000000000110111000000100",
			3597 => "00000000000000000011100001011001",
			3598 => "0000001000000000000001110000000100",
			3599 => "00000000000000000011100001011001",
			3600 => "00000000011001010011100001011001",
			3601 => "0000000000000000000011111100001000",
			3602 => "0000001010000000001100011100000100",
			3603 => "11111111101000010011100001011001",
			3604 => "00000000000000000011100001011001",
			3605 => "00000000000000000011100001011001",
			3606 => "0000000110000000000100111100001100",
			3607 => "0000000100000000001011101100000100",
			3608 => "00000000000000000011100010100101",
			3609 => "0000001001000000000010101100000100",
			3610 => "11111111011110010011100010100101",
			3611 => "00000000000000000011100010100101",
			3612 => "0000001100000000000001011000011000",
			3613 => "0000000000000000000010101000000100",
			3614 => "00000000000000000011100010100101",
			3615 => "0000000000000000000010111100010000",
			3616 => "0000001011000000000010001000000100",
			3617 => "00000000000000000011100010100101",
			3618 => "0000001001000000000010101100001000",
			3619 => "0000001101000000000111111100000100",
			3620 => "00000000000000000011100010100101",
			3621 => "00000000100001000011100010100101",
			3622 => "00000000000000000011100010100101",
			3623 => "00000000000000000011100010100101",
			3624 => "00000000000000000011100010100101",
			3625 => "0000001100000000001011000000001000",
			3626 => "0000001111000000000110111000000100",
			3627 => "11111111010111000011100011101001",
			3628 => "00000000000000000011100011101001",
			3629 => "0000001101000000001111100100011000",
			3630 => "0000001011000000000010001000000100",
			3631 => "00000000000000000011100011101001",
			3632 => "0000000100000000001011110000000100",
			3633 => "00000000000000000011100011101001",
			3634 => "0000000111000000000100010000001100",
			3635 => "0000000100000000001001001100001000",
			3636 => "0000001101000000001010001000000100",
			3637 => "00000000000000000011100011101001",
			3638 => "00000000011011000011100011101001",
			3639 => "00000000000000000011100011101001",
			3640 => "00000000000000000011100011101001",
			3641 => "11111111111001110011100011101001",
			3642 => "0000001001000000001010100100010100",
			3643 => "0000001100000000001000000000001000",
			3644 => "0000000000000000000001110100000100",
			3645 => "00000000000000000011100101000101",
			3646 => "11111111101101110011100101000101",
			3647 => "0000001100000000000010001000001000",
			3648 => "0000000100000000001001000000000100",
			3649 => "00000000000101010011100101000101",
			3650 => "00000000000000000011100101000101",
			3651 => "00000000000000000011100101000101",
			3652 => "0000001100000000001000011000011000",
			3653 => "0000001001000000000011101000010100",
			3654 => "0000000000000000000010101000000100",
			3655 => "00000000000000000011100101000101",
			3656 => "0000001100000000000100011000000100",
			3657 => "00000000000000000011100101000101",
			3658 => "0000001000000000001001101000001000",
			3659 => "0000001000000000000101000100000100",
			3660 => "00000000000000000011100101000101",
			3661 => "00000000100110100011100101000101",
			3662 => "00000000000000000011100101000101",
			3663 => "00000000000000000011100101000101",
			3664 => "00000000000000000011100101000101",
			3665 => "0000001110000000001011111000011000",
			3666 => "0000000000000000000001110100010100",
			3667 => "0000000110000000000100110100000100",
			3668 => "00000000000000000011100110110001",
			3669 => "0000000101000000000101110000001100",
			3670 => "0000001100000000001101010100000100",
			3671 => "00000000000000000011100110110001",
			3672 => "0000001000000000001000100100000100",
			3673 => "00000000000000000011100110110001",
			3674 => "00000000100111100011100110110001",
			3675 => "00000000000000000011100110110001",
			3676 => "00000000000000000011100110110001",
			3677 => "0000001100000000000001101000001100",
			3678 => "0000000010000000000110111000001000",
			3679 => "0000000001000000001100011000000100",
			3680 => "11111111010001010011100110110001",
			3681 => "00000000000000000011100110110001",
			3682 => "00000000000000000011100110110001",
			3683 => "0000001101000000001111100100010000",
			3684 => "0000001110000000001100001100000100",
			3685 => "00000000000000000011100110110001",
			3686 => "0000001001000000000010101100001000",
			3687 => "0000000000000000000100000000000100",
			3688 => "00000000011011110011100110110001",
			3689 => "00000000000000000011100110110001",
			3690 => "00000000000000000011100110110001",
			3691 => "00000000000000000011100110110001",
			3692 => "0000001100000000001011000000001000",
			3693 => "0000001110000000001000101000000100",
			3694 => "11111111001111110011101000001101",
			3695 => "00000000000000000011101000001101",
			3696 => "0000000111000000000100010000011000",
			3697 => "0000001011000000000010001000000100",
			3698 => "00000000000000000011101000001101",
			3699 => "0000000100000000001110111000010000",
			3700 => "0000000100000000001011110000000100",
			3701 => "00000000000000000011101000001101",
			3702 => "0000001101000000001010001000000100",
			3703 => "00000000000000000011101000001101",
			3704 => "0000001101000000001100000000000100",
			3705 => "00000000100100100011101000001101",
			3706 => "00000000000000000011101000001101",
			3707 => "00000000000000000011101000001101",
			3708 => "0000000100000000001011100000001100",
			3709 => "0000001100000000001111011100000100",
			3710 => "00000000000000000011101000001101",
			3711 => "0000001011000000000010110100000100",
			3712 => "00000000000000000011101000001101",
			3713 => "11111111101011010011101000001101",
			3714 => "00000000000000000011101000001101",
			3715 => "0000001001000000000111101100010100",
			3716 => "0000001110000000000001011100001100",
			3717 => "0000000100000000001100010000000100",
			3718 => "00000000000000000011101010001001",
			3719 => "0000001100000000001111011100000100",
			3720 => "11111111001100100011101010001001",
			3721 => "00000000000000000011101010001001",
			3722 => "0000000101000000000010000100000100",
			3723 => "00000000000101000011101010001001",
			3724 => "00000000000000000011101010001001",
			3725 => "0000001110000000001011101100010000",
			3726 => "0000000101000000001100100100000100",
			3727 => "00000000000000000011101010001001",
			3728 => "0000000000000000000111000100000100",
			3729 => "00000000000000000011101010001001",
			3730 => "0000000000000000001010101100000100",
			3731 => "00000000101110010011101010001001",
			3732 => "00000000000000000011101010001001",
			3733 => "0000000000000000000111000000001000",
			3734 => "0000001000000000000001010100000100",
			3735 => "00000000000000000011101010001001",
			3736 => "11111111100111000011101010001001",
			3737 => "0000000101000000000110111100010000",
			3738 => "0000000110000000001000010000000100",
			3739 => "00000000000000000011101010001001",
			3740 => "0000000101000000001001010000000100",
			3741 => "00000000000000000011101010001001",
			3742 => "0000000110000000001001111100000100",
			3743 => "00000000100101010011101010001001",
			3744 => "00000000000000000011101010001001",
			3745 => "00000000000000000011101010001001",
			3746 => "0000001100000000001000000000010100",
			3747 => "0000001001000000000000001000001000",
			3748 => "0000001110000000000010010100000100",
			3749 => "11111111000110110011101011111101",
			3750 => "00000000000000000011101011111101",
			3751 => "0000000101000000000111100000001000",
			3752 => "0000000101000000000010110100000100",
			3753 => "00000000000000000011101011111101",
			3754 => "11111111111101100011101011111101",
			3755 => "00000000000010100011101011111101",
			3756 => "0000000101000000000110111100100100",
			3757 => "0000000011000000000011110000011000",
			3758 => "0000001111000000001000110100010000",
			3759 => "0000000110000000000101010000001100",
			3760 => "0000000000000000001111001000000100",
			3761 => "00000000000000000011101011111101",
			3762 => "0000001001000000000010101100000100",
			3763 => "00000000101111100011101011111101",
			3764 => "00000000000000000011101011111101",
			3765 => "00000000000000000011101011111101",
			3766 => "0000000011000000001110000000000100",
			3767 => "11111111100111100011101011111101",
			3768 => "00000000000000000011101011111101",
			3769 => "0000001001000000000010101100001000",
			3770 => "0000000000000000000111111000000100",
			3771 => "00000000110110010011101011111101",
			3772 => "00000000000000000011101011111101",
			3773 => "00000000000000000011101011111101",
			3774 => "11111111100000010011101011111101",
			3775 => "0000001110000000001011111000011000",
			3776 => "0000000000000000000001110100010100",
			3777 => "0000000110000000000100110100000100",
			3778 => "00000000000000000011101101111001",
			3779 => "0000001011000000001011110100001100",
			3780 => "0000001100000000001101010100000100",
			3781 => "00000000000000000011101101111001",
			3782 => "0000001000000000001000100100000100",
			3783 => "00000000000000000011101101111001",
			3784 => "00000000101010010011101101111001",
			3785 => "00000000000000000011101101111001",
			3786 => "00000000000000000011101101111001",
			3787 => "0000001100000000000001101000010000",
			3788 => "0000000100000000000110001100001100",
			3789 => "0000000111000000000110100100000100",
			3790 => "00000000000000000011101101111001",
			3791 => "0000000110000000000101010000000100",
			3792 => "11111111010110000011101101111001",
			3793 => "00000000000000000011101101111001",
			3794 => "00000000000000000011101101111001",
			3795 => "0000001101000000001111100100010100",
			3796 => "0000001110000000001100001100001000",
			3797 => "0000000100000000001101001000000100",
			3798 => "00000000000000000011101101111001",
			3799 => "11111111111111110011101101111001",
			3800 => "0000001001000000000010101100001000",
			3801 => "0000000000000000000100000000000100",
			3802 => "00000000011110010011101101111001",
			3803 => "00000000000000000011101101111001",
			3804 => "00000000000000000011101101111001",
			3805 => "00000000000000000011101101111001",
			3806 => "0000001001000000000111101100011000",
			3807 => "0000001100000000001000000000001000",
			3808 => "0000001110000000001000101000000100",
			3809 => "11111111000101110011110000000101",
			3810 => "00000000000000000011110000000101",
			3811 => "0000000101000000001110110100001000",
			3812 => "0000001101000000000011001000000100",
			3813 => "00000000000000000011110000000101",
			3814 => "00000000000001010011110000000101",
			3815 => "0000001101000000001111010100000100",
			3816 => "00000000000000000011110000000101",
			3817 => "11111111111010100011110000000101",
			3818 => "0000001100000000000100011000010000",
			3819 => "0000001000000000000001010100001100",
			3820 => "0000001001000000000000001000000100",
			3821 => "00000000000000000011110000000101",
			3822 => "0000001110000000000110010000000100",
			3823 => "00000000000000000011110000000101",
			3824 => "00000000111001110011110000000101",
			3825 => "00000000000000000011110000000101",
			3826 => "0000000110000000001000010000001000",
			3827 => "0000000010000000000110101100000100",
			3828 => "00000000000000000011110000000101",
			3829 => "11111111011011000011110000000101",
			3830 => "0000001011000000000001000000010100",
			3831 => "0000001011000000000101110100001000",
			3832 => "0000001111000000000011000000000100",
			3833 => "00000000000000000011110000000101",
			3834 => "11111111111101010011110000000101",
			3835 => "0000000000000000000111000000000100",
			3836 => "00000000000000000011110000000101",
			3837 => "0000001000000000000111000100000100",
			3838 => "00000000111010000011110000000101",
			3839 => "00000000000000000011110000000101",
			3840 => "11111111110111100011110000000101",
			3841 => "0000000100000000001000110100011100",
			3842 => "0000001101000000001100010100011000",
			3843 => "0000000110000000001000010000010100",
			3844 => "0000000000000000000010101000010000",
			3845 => "0000000110000000000100110100000100",
			3846 => "00000000000000000011110001111001",
			3847 => "0000000010000000001000101000001000",
			3848 => "0000000111000000000011100000000100",
			3849 => "00000000000000000011110001111001",
			3850 => "00000000100000010011110001111001",
			3851 => "00000000000000000011110001111001",
			3852 => "00000000000000000011110001111001",
			3853 => "00000000000000000011110001111001",
			3854 => "00000000000000000011110001111001",
			3855 => "0000001110000000001000110100001000",
			3856 => "0000000001000000001110010100000100",
			3857 => "00000000000000000011110001111001",
			3858 => "11111111010011110011110001111001",
			3859 => "0000001101000000001111100100010100",
			3860 => "0000000111000000000111010000000100",
			3861 => "00000000000000000011110001111001",
			3862 => "0000000001000000000001000100000100",
			3863 => "00000000000000000011110001111001",
			3864 => "0000000001000000001100011000001000",
			3865 => "0000001110000000001000011100000100",
			3866 => "00000000000000000011110001111001",
			3867 => "00000000110000100011110001111001",
			3868 => "00000000000000000011110001111001",
			3869 => "00000000000000000011110001111001",
			3870 => "0000001110000000001110110100010000",
			3871 => "0000000111000000000110100100000100",
			3872 => "11111110011011010011110011101101",
			3873 => "0000000111000000000110100100001000",
			3874 => "0000001101000000000001000000000100",
			3875 => "00000000111101110011110011101101",
			3876 => "00000000000000000011110011101101",
			3877 => "11111111000011110011110011101101",
			3878 => "0000001101000000001111100100101000",
			3879 => "0000001110000000000110001100011000",
			3880 => "0000000000000000000010011000010100",
			3881 => "0000001010000000000011101000000100",
			3882 => "11111110110100010011110011101101",
			3883 => "0000000010000000001000100000001000",
			3884 => "0000000001000000001101111100000100",
			3885 => "00000010010001000011110011101101",
			3886 => "00000000011101000011110011101101",
			3887 => "0000000000000000000111000000000100",
			3888 => "11111111001011110011110011101101",
			3889 => "00000000101110000011110011101101",
			3890 => "11111110100111100011110011101101",
			3891 => "0000001000000000000111000100001100",
			3892 => "0000000111000000000101100100000100",
			3893 => "00000100001000000011110011101101",
			3894 => "0000000001000000001100011000000100",
			3895 => "00000001101010110011110011101101",
			3896 => "00000000000000000011110011101101",
			3897 => "00000000000000000011110011101101",
			3898 => "11111110100100110011110011101101",
			3899 => "0000000000000000001101010000101100",
			3900 => "0000000110000000001011001100000100",
			3901 => "00000000000000000011110101010001",
			3902 => "0000000011000000001101101100010100",
			3903 => "0000000101000000001100100100000100",
			3904 => "00000000000000000011110101010001",
			3905 => "0000000110000000001001100100000100",
			3906 => "00000000000000000011110101010001",
			3907 => "0000000000000000001010101100001000",
			3908 => "0000000000000000000110001000000100",
			3909 => "00000000000000000011110101010001",
			3910 => "00000000110010010011110101010001",
			3911 => "00000000000000000011110101010001",
			3912 => "0000001111000000000110111000000100",
			3913 => "11111111110011100011110101010001",
			3914 => "0000000110000000001000010000000100",
			3915 => "00000000000000000011110101010001",
			3916 => "0000000011000000000010010100000100",
			3917 => "00000000000000000011110101010001",
			3918 => "0000001010000000001000010100000100",
			3919 => "00000000000000000011110101010001",
			3920 => "00000000011000110011110101010001",
			3921 => "0000000010000000000011110100000100",
			3922 => "11111111111000110011110101010001",
			3923 => "00000000000000000011110101010001",
			3924 => "0000001001000000001010100000101000",
			3925 => "0000001100000000001011000000001000",
			3926 => "0000000100000000000110101100000100",
			3927 => "00000000000000000011110111100101",
			3928 => "11111111001010010011110111100101",
			3929 => "0000000010000000000010010100010000",
			3930 => "0000000110000000000100110100000100",
			3931 => "00000000000000000011110111100101",
			3932 => "0000000100000000001000011100001000",
			3933 => "0000001000000000001000100100000100",
			3934 => "00000000000000000011110111100101",
			3935 => "00000000001000100011110111100101",
			3936 => "00000000000000000011110111100101",
			3937 => "0000001110000000001011110000000100",
			3938 => "11111111011111010011110111100101",
			3939 => "0000000011000000001110111000001000",
			3940 => "0000001110000000001000000100000100",
			3941 => "00000000000000000011110111100101",
			3942 => "00000000010000000011110111100101",
			3943 => "00000000000000000011110111100101",
			3944 => "0000001100000000001011011100100000",
			3945 => "0000001011000000001011011100001000",
			3946 => "0000000100000000000011000000000100",
			3947 => "00000000000000000011110111100101",
			3948 => "11111111101111110011110111100101",
			3949 => "0000000000000000000111000100000100",
			3950 => "00000000000000000011110111100101",
			3951 => "0000000001000000001010011000010000",
			3952 => "0000001110000000001111101000001000",
			3953 => "0000001101000000000110010000000100",
			3954 => "00000001000111010011110111100101",
			3955 => "00000000000000000011110111100101",
			3956 => "0000001110000000000110001100000100",
			3957 => "11111111110110110011110111100101",
			3958 => "00000000110100110011110111100101",
			3959 => "00000000000000000011110111100101",
			3960 => "11111111101111100011110111100101",
			3961 => "0000001001000000001010100000101100",
			3962 => "0000000111000000001111011100001000",
			3963 => "0000000100000000000110101100000100",
			3964 => "00000000000000000011111010011001",
			3965 => "11111110110000110011111010011001",
			3966 => "0000001011000000000010110100010100",
			3967 => "0000000100000000000011001100010000",
			3968 => "0000001111000000000000010000000100",
			3969 => "00000000000000000011111010011001",
			3970 => "0000001010000000000011101000000100",
			3971 => "00000000000000000011111010011001",
			3972 => "0000000101000000001100010100000100",
			3973 => "00000000101010000011111010011001",
			3974 => "00000000000000000011111010011001",
			3975 => "00000000000000000011111010011001",
			3976 => "0000000011000000001000001000001100",
			3977 => "0000001100000000001111011100000100",
			3978 => "00000000000000000011111010011001",
			3979 => "0000001100000000000001011000000100",
			3980 => "11111111100011010011111010011001",
			3981 => "00000000000000000011111010011001",
			3982 => "00000000000000000011111010011001",
			3983 => "0000001100000000001001110100011100",
			3984 => "0000000000000000001000101100011000",
			3985 => "0000000101000000001100100100001000",
			3986 => "0000001100000000001010111000000100",
			3987 => "00000000001101000011111010011001",
			3988 => "00000000000000000011111010011001",
			3989 => "0000001100000000000100011000000100",
			3990 => "00000000000000000011111010011001",
			3991 => "0000000001000000001101111100000100",
			3992 => "00000000000000000011111010011001",
			3993 => "0000001001000000001010100000000100",
			3994 => "00000000000000000011111010011001",
			3995 => "00000001001110100011111010011001",
			3996 => "00000000000000000011111010011001",
			3997 => "0000000001000000000100110100001100",
			3998 => "0000001110000000000011000000000100",
			3999 => "00000000000000000011111010011001",
			4000 => "0000000101000000000111111100000100",
			4001 => "00000000000000000011111010011001",
			4002 => "00000000100001000011111010011001",
			4003 => "0000001011000000000101110100000100",
			4004 => "00000000000000000011111010011001",
			4005 => "11111111001100100011111010011001",
			4006 => "0000000111000000000110100100001100",
			4007 => "0000000001000000001101111100000100",
			4008 => "11111110011001010011111100010101",
			4009 => "0000001101000000001110000100000100",
			4010 => "00000010011010110011111100010101",
			4011 => "11111110110110100011111100010101",
			4012 => "0000001101000000001111100100110000",
			4013 => "0000000001000000001010011000101000",
			4014 => "0000000101000000001111010000010000",
			4015 => "0000001101000000000110100000000100",
			4016 => "00000011010010100011111100010101",
			4017 => "0000000001000000001101111100000100",
			4018 => "11111110011001110011111100010101",
			4019 => "0000001110000000001011101100000100",
			4020 => "00000001001101110011111100010101",
			4021 => "11111110100100000011111100010101",
			4022 => "0000000100000000000011101100001100",
			4023 => "0000000001000000001001011000000100",
			4024 => "00000110100011000011111100010101",
			4025 => "0000000110000000000100111100000100",
			4026 => "11111110100010100011111100010101",
			4027 => "00000001011111000011111100010101",
			4028 => "0000001110000000001001001100000100",
			4029 => "11111101101100110011111100010101",
			4030 => "0000000111000000001010010100000100",
			4031 => "00000000111011010011111100010101",
			4032 => "00000100110000010011111100010101",
			4033 => "0000001100000000001000000000000100",
			4034 => "00000010000000000011111100010101",
			4035 => "11111110011100010011111100010101",
			4036 => "11111110001100100011111100010101",
			4037 => "0000000111000000000110100100001100",
			4038 => "0000000001000000001101111100000100",
			4039 => "11111110011001100011111110011001",
			4040 => "0000001101000000001110000100000100",
			4041 => "00000001111011110011111110011001",
			4042 => "11111111000000000011111110011001",
			4043 => "0000001101000000001111100100110100",
			4044 => "0000001110000000000110001100100000",
			4045 => "0000000000000000001111000100011000",
			4046 => "0000000001000000001010011000010000",
			4047 => "0000000110000000001000010000001000",
			4048 => "0000000001000000001101011100000100",
			4049 => "00000010011110100011111110011001",
			4050 => "11111111110101110011111110011001",
			4051 => "0000001101000000001001011100000100",
			4052 => "11111110101011110011111110011001",
			4053 => "00000001110010110011111110011001",
			4054 => "0000001101000000001110010000000100",
			4055 => "00000001101001110011111110011001",
			4056 => "11111110011110000011111110011001",
			4057 => "0000001110000000001100001100000100",
			4058 => "11111101111111100011111110011001",
			4059 => "00000000000000000011111110011001",
			4060 => "0000000111000000000000011100000100",
			4061 => "00000111100111010011111110011001",
			4062 => "0000001000000000000111000100001100",
			4063 => "0000000001000000001100011000001000",
			4064 => "0000000100000000000011101100000100",
			4065 => "00000001101010010011111110011001",
			4066 => "00000010110111010011111110011001",
			4067 => "11111111101101100011111110011001",
			4068 => "11111111000111100011111110011001",
			4069 => "11111110001111110011111110011001",
			4070 => "0000000000000000000010101000100100",
			4071 => "0000001001000000001010100100011000",
			4072 => "0000000110000000001001100100010100",
			4073 => "0000001101000000000101110000010000",
			4074 => "0000000110000000000100110100000100",
			4075 => "00000000000000000100000000111101",
			4076 => "0000000111000000000001101000001000",
			4077 => "0000000111000000001000000000000100",
			4078 => "00000000000000000100000000111101",
			4079 => "00000000100110000100000000111101",
			4080 => "00000000000000000100000000111101",
			4081 => "00000000000000000100000000111101",
			4082 => "11111111100111010100000000111101",
			4083 => "0000000111000000001111011100001000",
			4084 => "0000000011000000000001011100000100",
			4085 => "00000001001111010100000000111101",
			4086 => "00000000000000000100000000111101",
			4087 => "00000000000000000100000000111101",
			4088 => "0000001110000000000001011100000100",
			4089 => "11111110111100010100000000111101",
			4090 => "0000001110000000001100001100011000",
			4091 => "0000000100000000001010110100010100",
			4092 => "0000001001000000001010100100001100",
			4093 => "0000000111000000000100010000001000",
			4094 => "0000000101000000000101110000000100",
			4095 => "00000000000000000100000000111101",
			4096 => "00000000111010000100000000111101",
			4097 => "00000000000000000100000000111101",
			4098 => "0000001110000000000011000000000100",
			4099 => "00000000000000000100000000111101",
			4100 => "11111111100011010100000000111101",
			4101 => "11111111010011100100000000111101",
			4102 => "0000001011000000000001000000010000",
			4103 => "0000001011000000000000110100000100",
			4104 => "00000000000000000100000000111101",
			4105 => "0000001001000000000010101100001000",
			4106 => "0000000000000000001100001000000100",
			4107 => "00000001001010100100000000111101",
			4108 => "00000000000000000100000000111101",
			4109 => "00000000000000000100000000111101",
			4110 => "11111111110011110100000000111101",
			4111 => "0000001100000000001010111000001000",
			4112 => "0000001001000000000010101100000100",
			4113 => "11111110011010110100000010111001",
			4114 => "00000000000000000100000010111001",
			4115 => "0000001101000000001111100100110100",
			4116 => "0000001110000000000101000000100100",
			4117 => "0000000100000000001010110100011100",
			4118 => "0000001110000000001111101000010000",
			4119 => "0000001001000000001010100100001000",
			4120 => "0000000110000000001111000000000100",
			4121 => "00000000110101010100000010111001",
			4122 => "11111111000111010100000010111001",
			4123 => "0000001100000000001000000000000100",
			4124 => "00000010001000000100000010111001",
			4125 => "11111111111111100100000010111001",
			4126 => "0000001001000000000010101100001000",
			4127 => "0000000111000000000111010000000100",
			4128 => "11111111010101010100000010111001",
			4129 => "00000001000100000100000010111001",
			4130 => "11111101111110100100000010111001",
			4131 => "0000001110000000001000110100000100",
			4132 => "11111110001100010100000010111001",
			4133 => "00000000000000000100000010111001",
			4134 => "0000000001000000001100011000001100",
			4135 => "0000000000000000001011000100001000",
			4136 => "0000000011000000000101000000000100",
			4137 => "00000000000000000100000010111001",
			4138 => "00000001101101000100000010111001",
			4139 => "00000000000000000100000010111001",
			4140 => "11111111010110010100000010111001",
			4141 => "11111110010110000100000010111001",
			4142 => "0000000100000000000010010100101000",
			4143 => "0000001110000000001011111000100100",
			4144 => "0000000110000000001011001100010000",
			4145 => "0000000100000000001100010000001100",
			4146 => "0000000100000000000010000100000100",
			4147 => "00000000000000000100000101111101",
			4148 => "0000001001000000001011001100000100",
			4149 => "00000000000110110100000101111101",
			4150 => "00000000000000000100000101111101",
			4151 => "11111111110101000100000101111101",
			4152 => "0000001010000000001000100100010000",
			4153 => "0000001010000000000011101000000100",
			4154 => "00000000000000000100000101111101",
			4155 => "0000001110000000000110010000000100",
			4156 => "00000000000000000100000101111101",
			4157 => "0000000101000000001110101100000100",
			4158 => "00000000000000000100000101111101",
			4159 => "00000001001101110100000101111101",
			4160 => "00000000000000000100000101111101",
			4161 => "11111111100111100100000101111101",
			4162 => "0000001110000000001000101000010000",
			4163 => "0000001001000000000010101100001000",
			4164 => "0000000001000000001010011000000100",
			4165 => "11111110101000100100000101111101",
			4166 => "00000000000000000100000101111101",
			4167 => "0000000001000000001010011000000100",
			4168 => "00000000001100110100000101111101",
			4169 => "00000000000000000100000101111101",
			4170 => "0000001110000000000011000000010000",
			4171 => "0000000110000000001000010000001100",
			4172 => "0000000010000000000010010100000100",
			4173 => "00000000000000000100000101111101",
			4174 => "0000000110000000000100111100000100",
			4175 => "00000000000000000100000101111101",
			4176 => "00000000110100010100000101111101",
			4177 => "00000000000000000100000101111101",
			4178 => "0000000001000000001100011000011000",
			4179 => "0000001100000000000100000100001100",
			4180 => "0000000110000000001000010000000100",
			4181 => "00000000000000000100000101111101",
			4182 => "0000001100000000001001110100000100",
			4183 => "00000000000000000100000101111101",
			4184 => "00000000101010100100000101111101",
			4185 => "0000000110000000001001111100001000",
			4186 => "0000001001000000001001111100000100",
			4187 => "00000000000000000100000101111101",
			4188 => "11111111000110000100000101111101",
			4189 => "00000000000000000100000101111101",
			4190 => "11111110101101000100000101111101",
			4191 => "0000001011000000000001000001000000",
			4192 => "0000001110000000001100001100110000",
			4193 => "0000000000000000001101010000101000",
			4194 => "0000001111000000001111101000010000",
			4195 => "0000001101000000001100010100001100",
			4196 => "0000001001000000001010100000000100",
			4197 => "00000000000000000100001000000001",
			4198 => "0000001001000000001010100100000100",
			4199 => "00000000110101000100001000000001",
			4200 => "00000000000000000100001000000001",
			4201 => "00000000000000000100001000000001",
			4202 => "0000001011000000001011110100001000",
			4203 => "0000000111000000001111011100000100",
			4204 => "11111111000101100100001000000001",
			4205 => "00000000000000000100001000000001",
			4206 => "0000000000000000000111000000001000",
			4207 => "0000000011000000000010010100000100",
			4208 => "00000000000000000100001000000001",
			4209 => "11111111110111010100001000000001",
			4210 => "0000001110000000000011000000000100",
			4211 => "00000000000000000100001000000001",
			4212 => "00000000101111110100001000000001",
			4213 => "0000000000000000001111000100000100",
			4214 => "00000000000000000100001000000001",
			4215 => "11111111001000100100001000000001",
			4216 => "0000001100000000000110100100000100",
			4217 => "00000000000000000100001000000001",
			4218 => "0000001001000000000010101100001000",
			4219 => "0000000000000000000100000000000100",
			4220 => "00000001000010110100001000000001",
			4221 => "00000000000000000100001000000001",
			4222 => "00000000000000000100001000000001",
			4223 => "11111111010111000100001000000001",
			4224 => "0000000100000000000010010100101000",
			4225 => "0000001110000000001011111000100100",
			4226 => "0000001000000000000101000100100000",
			4227 => "0000001010000000000011101000010100",
			4228 => "0000001011000000000111010000001100",
			4229 => "0000001011000000001010011100000100",
			4230 => "00000000000000000100001011001101",
			4231 => "0000000100000000001000001100000100",
			4232 => "00000000100011000100001011001101",
			4233 => "00000000000000000100001011001101",
			4234 => "0000001011000000000100000100000100",
			4235 => "00000000000000000100001011001101",
			4236 => "11111111110000000100001011001101",
			4237 => "0000001101000000001100100100000100",
			4238 => "00000000000000000100001011001101",
			4239 => "0000001110000000001110110100000100",
			4240 => "00000000000000000100001011001101",
			4241 => "00000001001010100100001011001101",
			4242 => "00000000000000000100001011001101",
			4243 => "11111111110001100100001011001101",
			4244 => "0000001110000000001000101000010100",
			4245 => "0000001001000000000010101100001100",
			4246 => "0000000100000000001011110000000100",
			4247 => "00000000000000000100001011001101",
			4248 => "0000000001000000001010011000000100",
			4249 => "11111110100110100100001011001101",
			4250 => "00000000000000000100001011001101",
			4251 => "0000000001000000001010011000000100",
			4252 => "00000000001101100100001011001101",
			4253 => "00000000000000000100001011001101",
			4254 => "0000000001000000001100011000100000",
			4255 => "0000001011000000000010110100010000",
			4256 => "0000001101000000000011001000000100",
			4257 => "00000000000000000100001011001101",
			4258 => "0000000100000000001110111000001000",
			4259 => "0000000100000000001000011100000100",
			4260 => "00000000000000000100001011001101",
			4261 => "00000001000100110100001011001101",
			4262 => "00000000000000000100001011001101",
			4263 => "0000001110000000001110100100000100",
			4264 => "11111111001010010100001011001101",
			4265 => "0000001101000000000000010000001000",
			4266 => "0000001011000000000111100000000100",
			4267 => "00000000100100000100001011001101",
			4268 => "00000000000000000100001011001101",
			4269 => "11111111010110000100001011001101",
			4270 => "0000001110000000000011000000001000",
			4271 => "0000001100000000001001110100000100",
			4272 => "00000000010110000100001011001101",
			4273 => "00000000000000000100001011001101",
			4274 => "11111110110100000100001011001101",
			4275 => "0000000010000000001110100101000100",
			4276 => "0000000010000000001110000000101100",
			4277 => "0000001110000000000110010000001100",
			4278 => "0000001100000000001011000000000100",
			4279 => "10111111100011110100001110101001",
			4280 => "0000001100000000001011000000000100",
			4281 => "11000001100011000100001110101001",
			4282 => "10111111101001010100001110101001",
			4283 => "0000001101000000001001100000011100",
			4284 => "0000000001000000001100011000010000",
			4285 => "0000000111000000000111010000001000",
			4286 => "0000001001000000001010100000000100",
			4287 => "10111111101110110100001110101001",
			4288 => "11000010111101010100001110101001",
			4289 => "0000000000000000000001110100000100",
			4290 => "11000100111101000100001110101001",
			4291 => "11100110101011010100001110101001",
			4292 => "0000000010000000001100111000000100",
			4293 => "11111000000000000100001110101001",
			4294 => "0000000001000000001100011000000100",
			4295 => "11001010111111100100001110101001",
			4296 => "11000001010111010100001110101001",
			4297 => "10111111100100100100001110101001",
			4298 => "0000001001000000000111101100001000",
			4299 => "0000000000000000000010011000000100",
			4300 => "00001010101010010100001110101001",
			4301 => "11000000001000110100001110101001",
			4302 => "0000001001000000001010100100001100",
			4303 => "0000000101000000000101110000000100",
			4304 => "10111111100111010100001110101001",
			4305 => "0000000111000000000000011100000100",
			4306 => "11101101010000000100001110101001",
			4307 => "11000101010110100100001110101001",
			4308 => "10111111100101000100001110101001",
			4309 => "0000001000000000001111001000100100",
			4310 => "0000001001000000000000001000001000",
			4311 => "0000000011000000001000000100000100",
			4312 => "10111111111001000100001110101001",
			4313 => "00001111111110110100001110101001",
			4314 => "0000001110000000000010111000010100",
			4315 => "0000001001000000001010100100001000",
			4316 => "0000000101000000000111111100000100",
			4317 => "10111111101010110100001110101001",
			4318 => "11101100001101000100001110101001",
			4319 => "0000001001000000000010101100001000",
			4320 => "0000000010000000000110001100000100",
			4321 => "11000000000000110100001110101001",
			4322 => "11000101110011110100001110101001",
			4323 => "10111111100101100100001110101001",
			4324 => "0000000001000000001010011000000100",
			4325 => "11110110001011100100001110101001",
			4326 => "11000000000000110100001110101001",
			4327 => "0000001000000000000111000100000100",
			4328 => "11000101010110100100001110101001",
			4329 => "10111111100100010100001110101001",
			4330 => "0000001001000000000111101100101100",
			4331 => "0000001100000000001000000000001000",
			4332 => "0000001111000000001000000100000100",
			4333 => "11111110100110000100010010001101",
			4334 => "00000000000000000100010010001101",
			4335 => "0000001101000000001010000100011100",
			4336 => "0000000001000000000101011100001100",
			4337 => "0000000001000000001101011100001000",
			4338 => "0000001111000000001011110000000100",
			4339 => "00000000001011000100010010001101",
			4340 => "00000000000000000100010010001101",
			4341 => "11111111100000000100010010001101",
			4342 => "0000000000000000000010101000000100",
			4343 => "00000000000000000100010010001101",
			4344 => "0000000100000000000011010100001000",
			4345 => "0000001010000000001010110000000100",
			4346 => "00000001000001110100010010001101",
			4347 => "00000000000000000100010010001101",
			4348 => "00000000000000000100010010001101",
			4349 => "0000001110000000000101000000000100",
			4350 => "11111111001011010100010010001101",
			4351 => "00000000000000000100010010001101",
			4352 => "0000000100000000001011110000011100",
			4353 => "0000001011000000000010001000010100",
			4354 => "0000001001000000000000001000000100",
			4355 => "00000000000000000100010010001101",
			4356 => "0000000000000000000010101000001100",
			4357 => "0000001101000000001100100100000100",
			4358 => "00000000000000000100010010001101",
			4359 => "0000001010000000000011101000000100",
			4360 => "00000000000000000100010010001101",
			4361 => "00000001010111000100010010001101",
			4362 => "00000000000000000100010010001101",
			4363 => "0000000011000000001011101100000100",
			4364 => "00000000000000000100010010001101",
			4365 => "11111111100100010100010010001101",
			4366 => "0000000111000000001111011100001100",
			4367 => "0000000001000000001010011000000100",
			4368 => "11111110110010100100010010001101",
			4369 => "0000000000000000001000110000000100",
			4370 => "00000000011111110100010010001101",
			4371 => "00000000000000000100010010001101",
			4372 => "0000000111000000000101100100010000",
			4373 => "0000001000000000001001101000001100",
			4374 => "0000000000000000000111000000000100",
			4375 => "00000000000000000100010010001101",
			4376 => "0000001001000000000010101100000100",
			4377 => "00000001011010010100010010001101",
			4378 => "00000000000000000100010010001101",
			4379 => "00000000000000000100010010001101",
			4380 => "0000000001000000000100110100001100",
			4381 => "0000001010000000000110011000000100",
			4382 => "00000000000000000100010010001101",
			4383 => "0000001100000000000001011000000100",
			4384 => "00000000011101100100010010001101",
			4385 => "00000000000000000100010010001101",
			4386 => "11111111010101100100010010001101",
			4387 => "0000001100000000001101010100000100",
			4388 => "11111110110001010100010100110001",
			4389 => "0000000111000000000101100100111000",
			4390 => "0000001001000000001010100100100100",
			4391 => "0000000110000000001001100100010100",
			4392 => "0000001001000000000000001000001000",
			4393 => "0000000001000000001001011000000100",
			4394 => "00000000000000000100010100110001",
			4395 => "11111111110111010100010100110001",
			4396 => "0000001100000000000100011000001000",
			4397 => "0000001101000000001100100100000100",
			4398 => "00000000000000000100010100110001",
			4399 => "00000001001010100100010100110001",
			4400 => "00000000000000000100010100110001",
			4401 => "0000000111000000000111010000000100",
			4402 => "11111110101001100100010100110001",
			4403 => "0000000100000000001010110100001000",
			4404 => "0000001100000000001000011000000100",
			4405 => "00000001000001100100010100110001",
			4406 => "00000000000000000100010100110001",
			4407 => "00000000000000000100010100110001",
			4408 => "0000000110000000001000010000001000",
			4409 => "0000000111000000001111011100000100",
			4410 => "00000001000001010100010100110001",
			4411 => "00000000000000000100010100110001",
			4412 => "0000001011000000000101110100000100",
			4413 => "11111111010000010100010100110001",
			4414 => "0000001001000000000010101100000100",
			4415 => "00000000111101010100010100110001",
			4416 => "00000000000000000100010100110001",
			4417 => "0000001110000000001000000100001000",
			4418 => "0000000001000000000101011100000100",
			4419 => "00000000000000000100010100110001",
			4420 => "11111110111100100100010100110001",
			4421 => "0000000111000000001010010100001100",
			4422 => "0000000001000000000100110100001000",
			4423 => "0000000000000000000100000000000100",
			4424 => "00000000111010100100010100110001",
			4425 => "00000000000000000100010100110001",
			4426 => "00000000000000000100010100110001",
			4427 => "11111111001000010100010100110001",
			4428 => "0000001000000000000001010100101100",
			4429 => "0000001101000000001100010100101000",
			4430 => "0000000110000000000100110100000100",
			4431 => "00000000000000000100010111101101",
			4432 => "0000001011000000001011011100011000",
			4433 => "0000000011000000000110111100001100",
			4434 => "0000001000000000001100011100001000",
			4435 => "0000001011000000000100000100000100",
			4436 => "00000000110011100100010111101101",
			4437 => "00000000000000000100010111101101",
			4438 => "00000000000000000100010111101101",
			4439 => "0000001100000000001101010100000100",
			4440 => "00000000000000000100010111101101",
			4441 => "0000000101000000000111100000000100",
			4442 => "11111111111001000100010111101101",
			4443 => "00000000000000000100010111101101",
			4444 => "0000001000000000001100011100000100",
			4445 => "00000000000000000100010111101101",
			4446 => "0000000111000000000001101000000100",
			4447 => "00000000000000000100010111101101",
			4448 => "00000001010011100100010111101101",
			4449 => "11111111101011100100010111101101",
			4450 => "0000001101000000001100010100001000",
			4451 => "0000001011000000001011110100000100",
			4452 => "11111110110111010100010111101101",
			4453 => "00000000000000000100010111101101",
			4454 => "0000000111000000000100010000010000",
			4455 => "0000000100000000001110111000001100",
			4456 => "0000000110000000001000010000000100",
			4457 => "00000000000000000100010111101101",
			4458 => "0000001001000000000010101100000100",
			4459 => "00000001000111110100010111101101",
			4460 => "00000000000000000100010111101101",
			4461 => "00000000000000000100010111101101",
			4462 => "0000000110000000001001111100010000",
			4463 => "0000000111000000000100010000000100",
			4464 => "00000000000000000100010111101101",
			4465 => "0000001011000000000010110100000100",
			4466 => "00000000000000000100010111101101",
			4467 => "0000001100000000001111011100000100",
			4468 => "00000000000000000100010111101101",
			4469 => "11111111001010110100010111101101",
			4470 => "0000000001000000000100110100001000",
			4471 => "0000000100000000000111011100000100",
			4472 => "00000000110110110100010111101101",
			4473 => "00000000000000000100010111101101",
			4474 => "00000000000000000100010111101101",
			4475 => "0000000001000000000101011100011000",
			4476 => "0000000000000000000111000000010100",
			4477 => "0000001110000000001010000100001100",
			4478 => "0000001100000000001011000000000100",
			4479 => "11111110011001110100011010110001",
			4480 => "0000000101000000000110100000000100",
			4481 => "00001000101101100100011010110001",
			4482 => "11111110011100110100011010110001",
			4483 => "0000001011000000001011110100000100",
			4484 => "00001100001010010100011010110001",
			4485 => "00000000000000000100011010110001",
			4486 => "11111110010111100100011010110001",
			4487 => "0000001001000000000010101101000100",
			4488 => "0000000101000000001001010000100000",
			4489 => "0000000100000000000110111000011000",
			4490 => "0000001001000000001010100000001100",
			4491 => "0000001001000000000000001000000100",
			4492 => "11111110011011100100011010110001",
			4493 => "0000000100000000001111100100000100",
			4494 => "00001100110111000100011010110001",
			4495 => "11111111011110100100011010110001",
			4496 => "0000001110000000001000001100000100",
			4497 => "00000111111111100100011010110001",
			4498 => "0000001010000000001000100100000100",
			4499 => "11111101110100100100011010110001",
			4500 => "00000001011011000100011010110001",
			4501 => "0000000001000000001100011000000100",
			4502 => "11111110010010100100011010110001",
			4503 => "00000000011111000100011010110001",
			4504 => "0000001000000000000001010100010000",
			4505 => "0000001001000000000101010000001000",
			4506 => "0000001011000000001011110100000100",
			4507 => "11111111101110110100011010110001",
			4508 => "00000001010000100100011010110001",
			4509 => "0000000111000000000101110100000100",
			4510 => "11111110011011010100011010110001",
			4511 => "11111100101011110100011010110001",
			4512 => "0000000101000000000111011000010000",
			4513 => "0000001100000000001000000000001000",
			4514 => "0000001110000000001111101000000100",
			4515 => "00001101010111100100011010110001",
			4516 => "00000001000001100100011010110001",
			4517 => "0000000110000000000100111100000100",
			4518 => "11111111001001110100011010110001",
			4519 => "00000001111001010100011010110001",
			4520 => "11111110000100010100011010110001",
			4521 => "0000000100000000001011110000000100",
			4522 => "00000001011001010100011010110001",
			4523 => "11111110011001010100011010110001",
			4524 => "0000000001000000000101011100010100",
			4525 => "0000000000000000000111000000010000",
			4526 => "0000000011000000001000100000001100",
			4527 => "0000001100000000001011000000000100",
			4528 => "11111110011001100100011101101101",
			4529 => "0000001011000000000000011100000100",
			4530 => "00001111011100110100011101101101",
			4531 => "11111110011100010100011101101101",
			4532 => "00000111101011110100011101101101",
			4533 => "11111110010111100100011101101101",
			4534 => "0000001001000000000010101101000100",
			4535 => "0000000101000000000101110000101000",
			4536 => "0000001001000000001010100000011000",
			4537 => "0000000010000000000110111100001000",
			4538 => "0000001010000000000011101000000100",
			4539 => "11111110011101110100011101101101",
			4540 => "00001101001011100100011101101101",
			4541 => "0000001101000000000111111100001000",
			4542 => "0000000101000000000111100000000100",
			4543 => "11111110011010000100011101101101",
			4544 => "11111111001010110100011101101101",
			4545 => "0000000101000000000101001000000100",
			4546 => "11111101010010000100011101101101",
			4547 => "11111110100100000100011101101101",
			4548 => "0000000010000000001111100100000100",
			4549 => "00001000111000000100011101101101",
			4550 => "0000000001000000001100011000000100",
			4551 => "11111110010001010100011101101101",
			4552 => "0000001010000000001001000100000100",
			4553 => "00000011110010100100011101101101",
			4554 => "11111110110100110100011101101101",
			4555 => "0000001010000000001000010100001100",
			4556 => "0000000111000000000000011100000100",
			4557 => "00000010000110110100011101101101",
			4558 => "0000000111000000000101110100000100",
			4559 => "11111110011001010100011101101101",
			4560 => "11111100011101010100011101101101",
			4561 => "0000000101000000000111011000001100",
			4562 => "0000000010000000001011110000000100",
			4563 => "00000110010100110100011101101101",
			4564 => "0000001010000000001001000100000100",
			4565 => "11111100110100010100011101101101",
			4566 => "00000010000000110100011101101101",
			4567 => "11111101110010100100011101101101",
			4568 => "0000000011000000000011000000000100",
			4569 => "00000011010101000100011101101101",
			4570 => "11111110011001000100011101101101",
			4571 => "0000000000000000000010101000111000",
			4572 => "0000001001000000000000001000010000",
			4573 => "0000000110000000001001100100000100",
			4574 => "11111111011011110100100001000001",
			4575 => "0000001010000000000111110100001000",
			4576 => "0000000000000000000110001000000100",
			4577 => "00000000000000000100100001000001",
			4578 => "00000000000101000100100001000001",
			4579 => "00000000000000000100100001000001",
			4580 => "0000000011000000001101101100100000",
			4581 => "0000001011000000001011011100011000",
			4582 => "0000001010000000000111110100001100",
			4583 => "0000000111000000000110100100001000",
			4584 => "0000001110000000001110110100000100",
			4585 => "00000000000000000100100001000001",
			4586 => "00000000110001110100100001000001",
			4587 => "00000000000000000100100001000001",
			4588 => "0000001111000000001000001100000100",
			4589 => "00000000000000000100100001000001",
			4590 => "0000001011000000000000011100000100",
			4591 => "00000000000000000100100001000001",
			4592 => "11111111101110010100100001000001",
			4593 => "0000000000000000000111000100000100",
			4594 => "00000000000000000100100001000001",
			4595 => "00000001100100110100100001000001",
			4596 => "0000000000000000000010101000000100",
			4597 => "11111111110111110100100001000001",
			4598 => "00000000000000000100100001000001",
			4599 => "0000001110000000000001011100000100",
			4600 => "11111110101000010100100001000001",
			4601 => "0000000111000000000111110000101000",
			4602 => "0000001101000000001100010100010100",
			4603 => "0000000110000000001000010000001100",
			4604 => "0000001100000000001011000000000100",
			4605 => "00000000000000000100100001000001",
			4606 => "0000001101000000000111111100000100",
			4607 => "00000000000000000100100001000001",
			4608 => "00000000011010010100100001000001",
			4609 => "0000000111000000001000011000000100",
			4610 => "00000000000000000100100001000001",
			4611 => "11111111000011000100100001000001",
			4612 => "0000000110000000001000010000000100",
			4613 => "00000000000000000100100001000001",
			4614 => "0000000000000000000010011000001000",
			4615 => "0000001001000000000010101100000100",
			4616 => "00000001001100110100100001000001",
			4617 => "00000000000000000100100001000001",
			4618 => "0000001110000000000110001100000100",
			4619 => "11111111110110000100100001000001",
			4620 => "00000000000000000100100001000001",
			4621 => "0000001101000000001000001100000100",
			4622 => "00000000000000000100100001000001",
			4623 => "11111111011011110100100001000001",
			4624 => "0000001011000000001010011100000100",
			4625 => "11111110011010100100100010110101",
			4626 => "0000000101000000001111010100110100",
			4627 => "0000001110000000001100001100100100",
			4628 => "0000000100000000001001001100100000",
			4629 => "0000000111000000000101100100010000",
			4630 => "0000000111000000001111011100001000",
			4631 => "0000001100000000001000000000000100",
			4632 => "00000000100100110100100010110101",
			4633 => "11111110000101000100100010110101",
			4634 => "0000001010000000000001010000000100",
			4635 => "00000001101000110100100010110101",
			4636 => "11111111010000110100100010110101",
			4637 => "0000001000000000001100000100001000",
			4638 => "0000001010000000001001000100000100",
			4639 => "11111110100111110100100010110101",
			4640 => "00000000000000000100100010110101",
			4641 => "0000000001000000001100011000000100",
			4642 => "00000001011011010100100010110101",
			4643 => "11111111101101110100100010110101",
			4644 => "11111101111110010100100010110101",
			4645 => "0000000001000000001100011000001100",
			4646 => "0000000000000000001011000100001000",
			4647 => "0000000011000000000110001100000100",
			4648 => "00000000000000000100100010110101",
			4649 => "00000001110000010100100010110101",
			4650 => "11111111011101000100100010110101",
			4651 => "11111111001001110100100010110101",
			4652 => "11111110001100100100100010110101",
			4653 => "0000001001000000000111101100110100",
			4654 => "0000001100000000001000000000001000",
			4655 => "0000001111000000001000000100000100",
			4656 => "11111110100011100100100110110001",
			4657 => "00000000000000000100100110110001",
			4658 => "0000000101000000001110110100100100",
			4659 => "0000000001000000000101011100010100",
			4660 => "0000001100000000001001110100001100",
			4661 => "0000000101000000000010011100001000",
			4662 => "0000001000000000001000010100000100",
			4663 => "00000000000000000100100110110001",
			4664 => "00000000100000110100100110110001",
			4665 => "00000000000000000100100110110001",
			4666 => "0000000101000000000011001000000100",
			4667 => "11111111010101100100100110110001",
			4668 => "00000000000000000100100110110001",
			4669 => "0000000000000000000010101000000100",
			4670 => "00000000000000000100100110110001",
			4671 => "0000000100000000000011010100001000",
			4672 => "0000001000000000001011010100000100",
			4673 => "00000001000010110100100110110001",
			4674 => "00000000000000000100100110110001",
			4675 => "00000000000000000100100110110001",
			4676 => "0000000001000000001110010100000100",
			4677 => "11111111000011100100100110110001",
			4678 => "00000000000000000100100110110001",
			4679 => "0000000100000000001011110000100000",
			4680 => "0000001011000000000010001000011000",
			4681 => "0000001001000000000000001000000100",
			4682 => "00000000000000000100100110110001",
			4683 => "0000000000000000000010101000010000",
			4684 => "0000000101000000001100100100001000",
			4685 => "0000000011000000001111010100000100",
			4686 => "00000000110110010100100110110001",
			4687 => "00000000000000000100100110110001",
			4688 => "0000001010000000000111110100000100",
			4689 => "00000000000000000100100110110001",
			4690 => "00000001101111000100100110110001",
			4691 => "00000000000000000100100110110001",
			4692 => "0000000011000000001011101100000100",
			4693 => "00000000000000000100100110110001",
			4694 => "11111111011011010100100110110001",
			4695 => "0000000111000000001111011100001100",
			4696 => "0000000001000000001010011000000100",
			4697 => "11111110101110010100100110110001",
			4698 => "0000000000000000001000110000000100",
			4699 => "00000000100111000100100110110001",
			4700 => "00000000000000000100100110110001",
			4701 => "0000000111000000000101100100010000",
			4702 => "0000001000000000001001101000001100",
			4703 => "0000000000000000000111000000000100",
			4704 => "00000000000000000100100110110001",
			4705 => "0000001001000000000010101100000100",
			4706 => "00000001100000010100100110110001",
			4707 => "00000000000000000100100110110001",
			4708 => "00000000000000000100100110110001",
			4709 => "0000000001000000000100110100001100",
			4710 => "0000000110000000000101010000000100",
			4711 => "00000000000000000100100110110001",
			4712 => "0000001100000000000001011000000100",
			4713 => "00000000100110110100100110110001",
			4714 => "00000000000000000100100110110001",
			4715 => "11111111010001010100100110110001",
			4716 => "0000001100000000001101010100000100",
			4717 => "11111110100111110100101001101101",
			4718 => "0000000100000000000011001100111100",
			4719 => "0000001010000000001000010100100000",
			4720 => "0000000011000000001100111000010100",
			4721 => "0000001001000000001010100100010000",
			4722 => "0000000001000000001001011000001000",
			4723 => "0000000110000000000100110100000100",
			4724 => "00000000000000000100101001101101",
			4725 => "00000000100001010100101001101101",
			4726 => "0000001011000000000100000100000100",
			4727 => "00000000000000000100101001101101",
			4728 => "11111111000011100100101001101101",
			4729 => "00000000111100110100101001101101",
			4730 => "0000001100000000001000000000000100",
			4731 => "00000000000000000100101001101101",
			4732 => "0000001000000000000001010100000100",
			4733 => "11111111011011010100101001101101",
			4734 => "00000000000000000100101001101101",
			4735 => "0000001101000000000010000100010100",
			4736 => "0000000111000000001000011000001000",
			4737 => "0000001010000000001000010100000100",
			4738 => "00000000000000000100101001101101",
			4739 => "11111111110100000100101001101101",
			4740 => "0000001010000000000001010000001000",
			4741 => "0000001101000000001001011100000100",
			4742 => "00000000000000000100101001101101",
			4743 => "00000001010111110100101001101101",
			4744 => "00000000000000000100101001101101",
			4745 => "0000001000000000001100000100000100",
			4746 => "11111111111001000100101001101101",
			4747 => "00000000000000000100101001101101",
			4748 => "0000001110000000001000110100001000",
			4749 => "0000000100000000000011001100000100",
			4750 => "00000000000000000100101001101101",
			4751 => "11111110111001100100101001101101",
			4752 => "0000000101000000001100010000010000",
			4753 => "0000001001000000001010100100001100",
			4754 => "0000000101000000001110010000000100",
			4755 => "00000000000000000100101001101101",
			4756 => "0000000001000000001011111100000100",
			4757 => "00000000000000000100101001101101",
			4758 => "00000001000111100100101001101101",
			4759 => "00000000000000000100101001101101",
			4760 => "0000000110000000001001111100000100",
			4761 => "11111111000011010100101001101101",
			4762 => "00000000000000000100101001101101",
			4763 => "0000000001000000000101011100000100",
			4764 => "11111110011010000100101100001001",
			4765 => "0000000001000000001100011001000100",
			4766 => "0000000101000000001001010000100000",
			4767 => "0000001001000000001010100000001100",
			4768 => "0000000010000000000110111100001000",
			4769 => "0000001001000000000000001000000100",
			4770 => "11111110100101100100101100001001",
			4771 => "00000100110010100100101100001001",
			4772 => "11111110011000110100101100001001",
			4773 => "0000000100000000000011000000000100",
			4774 => "00000011100000110100101100001001",
			4775 => "0000001101000000001001011100001000",
			4776 => "0000000001000000001100011000000100",
			4777 => "11111110010010000100101100001001",
			4778 => "00000000000000000100101100001001",
			4779 => "0000001011000000000010001000000100",
			4780 => "00001100011011100100101100001001",
			4781 => "11111111001100110100101100001001",
			4782 => "0000000110000000001000010000001100",
			4783 => "0000001101000000001100010100001000",
			4784 => "0000000110000000001011001100000100",
			4785 => "11111111100010000100101100001001",
			4786 => "00000011000100010100101100001001",
			4787 => "11111101101100100100101100001001",
			4788 => "0000000100000000000101010100001100",
			4789 => "0000000001000000001101111100000100",
			4790 => "00000001110100000100101100001001",
			4791 => "0000000100000000000101000000000100",
			4792 => "00000000111110100100101100001001",
			4793 => "00000011110010110100101100001001",
			4794 => "0000001110000000001110100100000100",
			4795 => "11111101100110010100101100001001",
			4796 => "0000001100000000001011011100000100",
			4797 => "00000001101111010100101100001001",
			4798 => "11111111111100100100101100001001",
			4799 => "0000000011000000000001011100000100",
			4800 => "00000010011110110100101100001001",
			4801 => "11111110011010010100101100001001",
			4802 => "0000001001000000001000010000000100",
			4803 => "11111110011010010100101110110101",
			4804 => "0000001001000000000010101101001100",
			4805 => "0000000101000000001001010000101000",
			4806 => "0000001001000000001010100100010100",
			4807 => "0000000010000000000110111100001000",
			4808 => "0000001001000000000000001000000100",
			4809 => "11111110100111010100101110110101",
			4810 => "00000011010010000100101110110101",
			4811 => "0000001100000000001000000000000100",
			4812 => "11111110011010010100101110110101",
			4813 => "0000000111000000000001101000000100",
			4814 => "00000101111010010100101110110101",
			4815 => "11111110011110100100101110110101",
			4816 => "0000000101000000001110000100001100",
			4817 => "0000001101000000000111111100001000",
			4818 => "0000000100000000000110111000000100",
			4819 => "00000011001001100100101110110101",
			4820 => "11111110111000100100101110110101",
			4821 => "00001000111111010100101110110101",
			4822 => "0000001011000000000100010000000100",
			4823 => "11111110001101100100101110110101",
			4824 => "00000000000000000100101110110101",
			4825 => "0000000110000000001000010000001100",
			4826 => "0000001101000000001100010100001000",
			4827 => "0000000011000000001011101100000100",
			4828 => "11111111100010000100101110110101",
			4829 => "00000010111011010100101110110101",
			4830 => "11111110001000110100101110110101",
			4831 => "0000000000000000001101010000001100",
			4832 => "0000001001000000000010101100001000",
			4833 => "0000001001000000001010100000000100",
			4834 => "00000001101101100100101110110101",
			4835 => "00000010101111010100101110110101",
			4836 => "11111110110100100100101110110101",
			4837 => "0000001110000000001000011100000100",
			4838 => "11111101110010110100101110110101",
			4839 => "0000001010000000000001010000000100",
			4840 => "11111111101111010100101110110101",
			4841 => "00000001101100100100101110110101",
			4842 => "0000001100000000001010111000000100",
			4843 => "00000000001100000100101110110101",
			4844 => "11111110011011010100101110110101",
			4845 => "0000000001000000000101011100000100",
			4846 => "11111110011010100100110001011001",
			4847 => "0000000001000000001100011001001000",
			4848 => "0000000101000000001001010000101000",
			4849 => "0000001001000000001010100000001100",
			4850 => "0000000010000000001100000000001000",
			4851 => "0000001111000000000111011000000100",
			4852 => "11111110111000100100110001011001",
			4853 => "00000001001010100100110001011001",
			4854 => "11111110011010100100110001011001",
			4855 => "0000000100000000000011000000001100",
			4856 => "0000000110000000001111000000000100",
			4857 => "00000011111000000100110001011001",
			4858 => "0000000111000000000001101000000100",
			4859 => "11111110111110100100110001011001",
			4860 => "00000010000001000100110001011001",
			4861 => "0000001101000000001001011100001000",
			4862 => "0000000001000000001100011000000100",
			4863 => "11111110010110000100110001011001",
			4864 => "00000000000000000100110001011001",
			4865 => "0000000101000000001110000100000100",
			4866 => "00001010110011110100110001011001",
			4867 => "11111111000011000100110001011001",
			4868 => "0000000110000000000100111100000100",
			4869 => "11111110010110100100110001011001",
			4870 => "0000000100000000001010110100010000",
			4871 => "0000000000000000000010101000001000",
			4872 => "0000000100000000001110000000000100",
			4873 => "00000011010000100100110001011001",
			4874 => "11111110100010000100110001011001",
			4875 => "0000000111000000001011011100000100",
			4876 => "00000010100000110100110001011001",
			4877 => "00000001010011110100110001011001",
			4878 => "0000000011000000001100001100000100",
			4879 => "11111110000110100100110001011001",
			4880 => "0000001101000000000111010100000100",
			4881 => "00000001101010100100110001011001",
			4882 => "11111111111101010100110001011001",
			4883 => "0000000011000000000001011100000100",
			4884 => "00000001111001000100110001011001",
			4885 => "11111110011011000100110001011001",
			4886 => "0000000111000000000011100000000100",
			4887 => "11111110011100110100110100001101",
			4888 => "0000001110000000001011111000011100",
			4889 => "0000001010000000000011101000001000",
			4890 => "0000000001000000001111001100000100",
			4891 => "00000001000011010100110100001101",
			4892 => "11111110110011110100110100001101",
			4893 => "0000000000000000000001110100010000",
			4894 => "0000001110000000000110010000000100",
			4895 => "00000000000000000100110100001101",
			4896 => "0000000100000000000010010100001000",
			4897 => "0000000000000000001011010100000100",
			4898 => "00000000000000000100110100001101",
			4899 => "00000001101000000100110100001101",
			4900 => "00000000000000000100110100001101",
			4901 => "11111111000110110100110100001101",
			4902 => "0000000000000000000010101000000100",
			4903 => "11111110011001000100110100001101",
			4904 => "0000001100000000001000011000011100",
			4905 => "0000000001000000001100011000001100",
			4906 => "0000000101000000001001010000000100",
			4907 => "11111110011110100100110100001101",
			4908 => "0000001110000000000010010100000100",
			4909 => "11111111110111110100110100001101",
			4910 => "00000001000111110100110100001101",
			4911 => "0000001011000000000010001000001000",
			4912 => "0000001011000000000110110100000100",
			4913 => "00000000110000010100110100001101",
			4914 => "11111111100011000100110100001101",
			4915 => "0000001001000000000010101100000100",
			4916 => "00000001111000000100110100001101",
			4917 => "00000000000000000100110100001101",
			4918 => "0000001110000000001000011100001100",
			4919 => "0000000100000000001101001000001000",
			4920 => "0000001000000000000001110000000100",
			4921 => "11111111000010000100110100001101",
			4922 => "00000000011000110100110100001101",
			4923 => "11111110100000110100110100001101",
			4924 => "0000001011000000000001000000001000",
			4925 => "0000000001000000000100110100000100",
			4926 => "00000001011011100100110100001101",
			4927 => "11111111010001110100110100001101",
			4928 => "0000001101000000001111100100000100",
			4929 => "00000000000000000100110100001101",
			4930 => "11111110101011110100110100001101",
			4931 => "0000000111000000001000000000000100",
			4932 => "11111110100000000100111000000011",
			4933 => "0000000001000000001101111100101100",
			4934 => "0000000111000000000111010000010100",
			4935 => "0000001111000000001010001000001100",
			4936 => "0000001111000000001001011100000100",
			4937 => "00000000000000000100111000000011",
			4938 => "0000001000000000000011101000000100",
			4939 => "00000000000000000100111000000011",
			4940 => "00000000111011110100111000000011",
			4941 => "0000000111000000000111010000000100",
			4942 => "11111110100000010100111000000011",
			4943 => "00000000000000000100111000000011",
			4944 => "0000001101000000001111010100010000",
			4945 => "0000000001000000000001111000001100",
			4946 => "0000000110000000000100111100000100",
			4947 => "00000000000000000100111000000011",
			4948 => "0000000000000000000011010000000100",
			4949 => "00000001010011010100111000000011",
			4950 => "00000000000000000100111000000011",
			4951 => "11111111101110000100111000000011",
			4952 => "0000000001000000001110010100000100",
			4953 => "11111110101001010100111000000011",
			4954 => "00000000000000000100111000000011",
			4955 => "0000000001000000000100110100100000",
			4956 => "0000001101000000001001011100010000",
			4957 => "0000000110000000001111000000001100",
			4958 => "0000000001000000001101111100001000",
			4959 => "0000000001000000001101111100000100",
			4960 => "00000000000000000100111000000011",
			4961 => "00000001000110100100111000000011",
			4962 => "00000000000000000100111000000011",
			4963 => "11111111001000100100111000000011",
			4964 => "0000000110000000001000010000000100",
			4965 => "00000000000000000100111000000011",
			4966 => "0000000001000000001101111100000100",
			4967 => "00000000000000000100111000000011",
			4968 => "0000000111000000001000011000000100",
			4969 => "00000000000000000100111000000011",
			4970 => "00000010000001110100111000000011",
			4971 => "0000000001000000001100011000011100",
			4972 => "0000000011000000001100111000001100",
			4973 => "0000001011000000001011011100001000",
			4974 => "0000001011000000000000011100000100",
			4975 => "00000000000000000100111000000011",
			4976 => "11111111111001000100111000000011",
			4977 => "00000001001001110100111000000011",
			4978 => "0000000000000000000111000000001000",
			4979 => "0000001011000000000100010000000100",
			4980 => "00000000000000000100111000000011",
			4981 => "11111110101000010100111000000011",
			4982 => "0000001000000000000001110000000100",
			4983 => "00000000111110100100111000000011",
			4984 => "11111111101011110100111000000011",
			4985 => "0000000111000000000000011100001100",
			4986 => "0000001011000000001011011100000100",
			4987 => "00000000000000000100111000000011",
			4988 => "0000001000000000001001101000000100",
			4989 => "00000001100011110100111000000011",
			4990 => "00000000000000000100111000000011",
			4991 => "11111111100000010100111000000011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1652, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(3300, initial_addr_3'length));
	end generate gen_rom_10;

	gen_rom_11: if SELECT_ROM = 11 generate
		bank <= (
			0 => "00000000000000000000000000000101",
			1 => "00000000000000000000000000001001",
			2 => "00000000000000000000000000001101",
			3 => "00000000000000000000000000010001",
			4 => "00000000000000000000000000010101",
			5 => "00000000000000000000000000011001",
			6 => "00000000000000000000000000011101",
			7 => "00000000000000000000000000100001",
			8 => "00000000000000000000000000100101",
			9 => "00000000000000000000000000101001",
			10 => "00000000000000000000000000101101",
			11 => "00000000000000000000000000110001",
			12 => "00000000000000000000000000110101",
			13 => "00000000000000000000000000111001",
			14 => "00000000000000000000000000111101",
			15 => "00000000000000000000000001000001",
			16 => "00000000000000000000000001000101",
			17 => "00000000000000000000000001001001",
			18 => "00000000000000000000000001001101",
			19 => "00000000000000000000000001010001",
			20 => "00000000000000000000000001010101",
			21 => "00000000000000000000000001011001",
			22 => "00000000000000000000000001011101",
			23 => "00000000000000000000000001100001",
			24 => "00000000000000000000000001100101",
			25 => "00000000000000000000000001101001",
			26 => "00000000000000000000000001101101",
			27 => "00000000000000000000000001110001",
			28 => "0000000001000000001101111100000100",
			29 => "11111111111111110000000001111101",
			30 => "00000000000000000000000001111101",
			31 => "0000001000000000001100011100000100",
			32 => "00000000000000000000000010001001",
			33 => "11111111111110110000000010001001",
			34 => "0000000010000000001011111000001000",
			35 => "0000001110000000000110010000000100",
			36 => "00000000000000000000000010011101",
			37 => "11111111110111110000000010011101",
			38 => "00000000000000000000000010011101",
			39 => "0000001001000000000111101100001000",
			40 => "0000000000000000000110001000000100",
			41 => "00000000000000000000000010110001",
			42 => "11111111101000000000000010110001",
			43 => "00000000000000000000000010110001",
			44 => "0000000001000000000111101000001000",
			45 => "0000001001000000000111101100000100",
			46 => "11111111111010100000000011000101",
			47 => "00000000000000000000000011000101",
			48 => "00000000000000000000000011000101",
			49 => "0000001001000000000000001000001000",
			50 => "0000000001000000001101111100000100",
			51 => "11111111111110000000000011011001",
			52 => "00000000000000000000000011011001",
			53 => "00000000000000000000000011011001",
			54 => "0000001000000000000001010100001100",
			55 => "0000000001000000001011111100000100",
			56 => "00000000000000000000000011110101",
			57 => "0000000001000000001100011000000100",
			58 => "00000000001101010000000011110101",
			59 => "00000000000000000000000011110101",
			60 => "00000000000000000000000011110101",
			61 => "0000000001000000000100110100001100",
			62 => "0000001110000000000110010000000100",
			63 => "00000000000000000000000100010001",
			64 => "0000000100000000000011001100000100",
			65 => "11111111110010010000000100010001",
			66 => "00000000000000000000000100010001",
			67 => "00000000000000000000000100010001",
			68 => "0000001001000000001001111100001000",
			69 => "0000000100000000001100010000000100",
			70 => "00000000000000000000000100111101",
			71 => "11111111100110000000000100111101",
			72 => "0000001110000000001100000000001000",
			73 => "0000000100000000001111100100000100",
			74 => "00000000000000000000000100111101",
			75 => "00000000001111000000000100111101",
			76 => "0000000100000000001111101000000100",
			77 => "11111111100000000000000100111101",
			78 => "00000000000000000000000100111101",
			79 => "0000001110000000000110010000001100",
			80 => "0000001001000000000101010000000100",
			81 => "00000000000000000000000101101001",
			82 => "0000000000000000001100000100000100",
			83 => "00000000000000000000000101101001",
			84 => "00000000001011100000000101101001",
			85 => "0000001001000000000111101100001000",
			86 => "0000001101000000001110101100000100",
			87 => "00000000000000000000000101101001",
			88 => "11111111101010000000000101101001",
			89 => "00000000000000000000000101101001",
			90 => "0000000001000000001110010100000100",
			91 => "00000000000000000000000110001101",
			92 => "0000001001000000001010100100001100",
			93 => "0000001000000000000001110000001000",
			94 => "0000001000000000001010110000000100",
			95 => "00000000000000000000000110001101",
			96 => "00000000001010100000000110001101",
			97 => "00000000000000000000000110001101",
			98 => "00000000000000000000000110001101",
			99 => "0000001110000000000110010000000100",
			100 => "00000000000000000000000110110001",
			101 => "0000000001000000001101111100001100",
			102 => "0000001100000000001011000000001000",
			103 => "0000001100000000000100001000000100",
			104 => "00000000000000000000000110110001",
			105 => "11111111101111000000000110110001",
			106 => "00000000000000000000000110110001",
			107 => "00000000000000000000000110110001",
			108 => "0000001001000000000111101100001000",
			109 => "0000001011000000000100000100000100",
			110 => "00000000000000000000000111011101",
			111 => "11111111101000000000000111011101",
			112 => "0000001100000000001010111000000100",
			113 => "00000000000000000000000111011101",
			114 => "0000001101000000001111010000001000",
			115 => "0000001010000000001000010100000100",
			116 => "00000000011111110000000111011101",
			117 => "00000000000000000000000111011101",
			118 => "00000000000000000000000111011101",
			119 => "0000001001000000000111101100001100",
			120 => "0000000010000000001000001100001000",
			121 => "0000001000000000001010110000000100",
			122 => "00000000000000000000001000010001",
			123 => "11111111100111010000001000010001",
			124 => "00000000000000000000001000010001",
			125 => "0000000110000000001111000000001000",
			126 => "0000001100000000001011000000000100",
			127 => "00000000011010110000001000010001",
			128 => "00000000000000000000001000010001",
			129 => "0000000010000000001100111000000100",
			130 => "11111111111110110000001000010001",
			131 => "00000000000000000000001000010001",
			132 => "0000000001000000001110010100001000",
			133 => "0000000000000000001001101000000100",
			134 => "00000000000000000000001001000101",
			135 => "11111111111100010000001001000101",
			136 => "0000001101000000000111111100010000",
			137 => "0000000100000000000001011100000100",
			138 => "00000000000000000000001001000101",
			139 => "0000001110000000001011111000001000",
			140 => "0000000000000000000110001000000100",
			141 => "00000000000000000000001001000101",
			142 => "00000000011111000000001001000101",
			143 => "00000000000000000000001001000101",
			144 => "00000000000000000000001001000101",
			145 => "0000000010000000001010000100010000",
			146 => "0000001100000000001000000000001100",
			147 => "0000001110000000000010000000000100",
			148 => "00000000000000000000001010001001",
			149 => "0000000110000000001001100100000100",
			150 => "11111111101011110000001010001001",
			151 => "00000000000000000000001010001001",
			152 => "00000000000000000000001010001001",
			153 => "0000001111000000001000001100001100",
			154 => "0000000100000000001011101100000100",
			155 => "00000000000000000000001010001001",
			156 => "0000001010000000001000010100000100",
			157 => "00000000011100100000001010001001",
			158 => "00000000000000000000001010001001",
			159 => "0000000100000000000010010100000100",
			160 => "11111111110010010000001010001001",
			161 => "00000000000000000000001010001001",
			162 => "0000000001000000000100110100011000",
			163 => "0000001110000000000110010000010000",
			164 => "0000001110000000001110101000000100",
			165 => "00000000000000000000001010111101",
			166 => "0000000110000000001010011000000100",
			167 => "00000000000000000000001010111101",
			168 => "0000001111000000000000010000000100",
			169 => "00000000001110010000001010111101",
			170 => "00000000000000000000001010111101",
			171 => "0000000100000000000011001100000100",
			172 => "11111111100100100000001010111101",
			173 => "00000000000000000000001010111101",
			174 => "00000000000000000000001010111101",
			175 => "0000001100000000001010111000011000",
			176 => "0000001101000000001100100100001100",
			177 => "0000000001000000001011111100000100",
			178 => "11111111011110010000001100011001",
			179 => "0000001000000000000001110000000100",
			180 => "00000000010100000000001100011001",
			181 => "00000000000000000000001100011001",
			182 => "0000000100000000001101101100001000",
			183 => "0000000101000000000010110100000100",
			184 => "00000000000000000000001100011001",
			185 => "11111110111011010000001100011001",
			186 => "00000000000000000000001100011001",
			187 => "0000001101000000000010011100010000",
			188 => "0000001001000000001001111100000100",
			189 => "00000000000000000000001100011001",
			190 => "0000000100000000000001011100000100",
			191 => "00000000000000000000001100011001",
			192 => "0000001110000000001011111000000100",
			193 => "00000000110100000000001100011001",
			194 => "00000000000000000000001100011001",
			195 => "0000001110000000001111010100000100",
			196 => "00000000000000000000001100011001",
			197 => "11111111111001000000001100011001",
			198 => "0000000001000000001110010100001100",
			199 => "0000001001000000000100101100001000",
			200 => "0000000100000000001100010000000100",
			201 => "00000000000000000000001101011101",
			202 => "11111111111001010000001101011101",
			203 => "00000000000000000000001101011101",
			204 => "0000001101000000000111111100010100",
			205 => "0000000100000000000001011100000100",
			206 => "00000000000000000000001101011101",
			207 => "0000001110000000001011111000001100",
			208 => "0000000110000000000100111100001000",
			209 => "0000000000000000000110001000000100",
			210 => "00000000000000000000001101011101",
			211 => "00000000100100110000001101011101",
			212 => "00000000000000000000001101011101",
			213 => "00000000000000000000001101011101",
			214 => "00000000000000000000001101011101",
			215 => "0000000010000000001011111000011000",
			216 => "0000001010000000000111110100010100",
			217 => "0000000011000000001111010100010000",
			218 => "0000000100000000001111100100001000",
			219 => "0000000011000000001110110100000100",
			220 => "00000000000000000000001110110001",
			221 => "11111111110001000000001110110001",
			222 => "0000001111000000000110010000000100",
			223 => "00000000000000000000001110110001",
			224 => "00000000011110100000001110110001",
			225 => "00000000000000000000001110110001",
			226 => "11111110111001100000001110110001",
			227 => "0000000011000000001011111000001100",
			228 => "0000000110000000000100111100001000",
			229 => "0000000001000000000001000100000100",
			230 => "00000000000000000000001110110001",
			231 => "00000000111101100000001110110001",
			232 => "00000000000000000000001110110001",
			233 => "0000000001000000001101111100000100",
			234 => "11111111101011100000001110110001",
			235 => "00000000000000000000001110110001",
			236 => "0000000010000000001100000000000100",
			237 => "00000000000000000000001111100101",
			238 => "0000000010000000001111101000010100",
			239 => "0000000001000000000001000100000100",
			240 => "00000000000000000000001111100101",
			241 => "0000000001000000001100011000001100",
			242 => "0000000110000000001101011000000100",
			243 => "00000000000000000000001111100101",
			244 => "0000000110000000001000010000000100",
			245 => "00000000001011010000001111100101",
			246 => "00000000000000000000001111100101",
			247 => "00000000000000000000001111100101",
			248 => "00000000000000000000001111100101",
			249 => "0000001100000000001010111100001100",
			250 => "0000000001000000000111101000001000",
			251 => "0000001000000000000001010000000100",
			252 => "00000000000000000000010001000001",
			253 => "11111111100101010000010001000001",
			254 => "00000000000000000000010001000001",
			255 => "0000001110000000001110110100001100",
			256 => "0000001010000000001010100000000100",
			257 => "00000000000000000000010001000001",
			258 => "0000001001000000000101010000000100",
			259 => "00000000000000000000010001000001",
			260 => "00000000101001000000010001000001",
			261 => "0000000100000000000011000000001100",
			262 => "0000001001000000001010100000001000",
			263 => "0000000001000000000001111000000100",
			264 => "00000000000000000000010001000001",
			265 => "11111111100001010000010001000001",
			266 => "00000000000000000000010001000001",
			267 => "0000000011000000001111100100001000",
			268 => "0000000001000000000111101000000100",
			269 => "00000000000000000000010001000001",
			270 => "00000000011100110000010001000001",
			271 => "00000000000000000000010001000001",
			272 => "0000001100000000001010111000010000",
			273 => "0000001000000000001100011100000100",
			274 => "00000000000000000000010010100101",
			275 => "0000001001000000000000001000001000",
			276 => "0000000111000000001001001000000100",
			277 => "11111110010010010000010010100101",
			278 => "00000000000000000000010010100101",
			279 => "00000000000000000000010010100101",
			280 => "0000001100000000000100011000010000",
			281 => "0000000000000000001111001000000100",
			282 => "00000000000000000000010010100101",
			283 => "0000001000000000000001010100001000",
			284 => "0000001110000000001011111000000100",
			285 => "00000000110111010000010010100101",
			286 => "00000000000000000000010010100101",
			287 => "00000000000000000000010010100101",
			288 => "0000001110000000001100010000001000",
			289 => "0000000001000000001110010100000100",
			290 => "00000000000000000000010010100101",
			291 => "00000000000100110000010010100101",
			292 => "0000000100000000001011110000001000",
			293 => "0000001000000000001010110000000100",
			294 => "00000000000000000000010010100101",
			295 => "11111110111110000000010010100101",
			296 => "00000000000000000000010010100101",
			297 => "0000001100000000001010111100010000",
			298 => "0000000001000000000111101000001100",
			299 => "0000000000000000001011010100000100",
			300 => "00000000000000000000010100001001",
			301 => "0000000111000000001000000000000100",
			302 => "11111111011101000000010100001001",
			303 => "00000000000000000000010100001001",
			304 => "00000000000000000000010100001001",
			305 => "0000000111000000001001001000001100",
			306 => "0000001001000000001010100000001000",
			307 => "0000000001000000000001000100000100",
			308 => "00000000000000000000010100001001",
			309 => "00000000110000000000010100001001",
			310 => "00000000000000000000010100001001",
			311 => "0000001110000000001100010000001100",
			312 => "0000000010000000001100000000000100",
			313 => "00000000000000000000010100001001",
			314 => "0000000001000000001110010100000100",
			315 => "00000000000000000000010100001001",
			316 => "00000000010101110000010100001001",
			317 => "0000000001000000001101111100001000",
			318 => "0000001100000000001000000000000100",
			319 => "11111111010100000000010100001001",
			320 => "00000000000000000000010100001001",
			321 => "00000000000000000000010100001001",
			322 => "0000000010000000001010000100001100",
			323 => "0000001000000000001010110000000100",
			324 => "00000000000000000000010101100101",
			325 => "0000000110000000001001100100000100",
			326 => "11111111010010000000010101100101",
			327 => "00000000000000000000010101100101",
			328 => "0000001110000000001100010000001000",
			329 => "0000001001000000000101010000000100",
			330 => "00000000000000000000010101100101",
			331 => "00000000101011000000010101100101",
			332 => "0000001001000000000000001000010000",
			333 => "0000001100000000001000000000001100",
			334 => "0000001101000000000001000000000100",
			335 => "00000000000000000000010101100101",
			336 => "0000000001000000001101111100000100",
			337 => "11111111010100100000010101100101",
			338 => "00000000000000000000010101100101",
			339 => "00000000000000000000010101100101",
			340 => "0000001011000000000101100100001000",
			341 => "0000001010000000001000010100000100",
			342 => "00000000010010010000010101100101",
			343 => "00000000000000000000010101100101",
			344 => "00000000000000000000010101100101",
			345 => "0000000001000000001011111100001000",
			346 => "0000000110000000001001100100000100",
			347 => "11111111001110100000010111000001",
			348 => "00000000000000000000010111000001",
			349 => "0000001110000000001100000000001100",
			350 => "0000000100000000001111100100000100",
			351 => "00000000000000000000010111000001",
			352 => "0000001100000000001011000000000100",
			353 => "00000000101110010000010111000001",
			354 => "00000000000000000000010111000001",
			355 => "0000000100000000000010010100001100",
			356 => "0000000001000000001101111100001000",
			357 => "0000001111000000000111010100000100",
			358 => "00000000000000000000010111000001",
			359 => "11111111001011010000010111000001",
			360 => "00000000000000000000010111000001",
			361 => "0000001101000000000111111100001100",
			362 => "0000000000000000000111000000001000",
			363 => "0000001111000000001000101000000100",
			364 => "00000000011111000000010111000001",
			365 => "00000000000000000000010111000001",
			366 => "00000000000000000000010111000001",
			367 => "00000000000000000000010111000001",
			368 => "0000000010000000001011111000011000",
			369 => "0000001010000000000111110100010100",
			370 => "0000001110000000001100010000001100",
			371 => "0000000100000000001111100100000100",
			372 => "00000000000000000000011000101101",
			373 => "0000001111000000000110010000000100",
			374 => "00000000000000000000011000101101",
			375 => "00000000011110000000011000101101",
			376 => "0000000100000000001000101000000100",
			377 => "11111111110100110000011000101101",
			378 => "00000000000000000000011000101101",
			379 => "11111110110100110000011000101101",
			380 => "0000000011000000001011111000010100",
			381 => "0000000110000000000100111100010000",
			382 => "0000001101000000000010011100001100",
			383 => "0000000111000000000111001000000100",
			384 => "00000000000000000000011000101101",
			385 => "0000000110000000001011001100000100",
			386 => "00000000000000000000011000101101",
			387 => "00000001000011110000011000101101",
			388 => "00000000000000000000011000101101",
			389 => "00000000000000000000011000101101",
			390 => "0000001011000000000111010000000100",
			391 => "00000000000000000000011000101101",
			392 => "0000000111000000001000011000000100",
			393 => "11111111101100100000011000101101",
			394 => "00000000000000000000011000101101",
			395 => "0000000010000000000110111100010000",
			396 => "0000001111000000001111010100001100",
			397 => "0000000110000000001001100100001000",
			398 => "0000000100000000001100010000000100",
			399 => "00000000000000000000011010001001",
			400 => "11111111101001100000011010001001",
			401 => "00000000000000000000011010001001",
			402 => "00000000000000000000011010001001",
			403 => "0000000100000000000001011100001000",
			404 => "0000001111000000001000001100000100",
			405 => "00000000000000000000011010001001",
			406 => "11111111111111010000011010001001",
			407 => "0000001111000000000011000000010100",
			408 => "0000000110000000001101011000000100",
			409 => "00000000000000000000011010001001",
			410 => "0000001100000000000100001000000100",
			411 => "00000000000000000000011010001001",
			412 => "0000000110000000000100111100001000",
			413 => "0000000001000000000001000100000100",
			414 => "00000000000000000000011010001001",
			415 => "00000000101011010000011010001001",
			416 => "00000000000000000000011010001001",
			417 => "00000000000000000000011010001001",
			418 => "0000001100000000001010111000011000",
			419 => "0000001101000000001100100100001100",
			420 => "0000000001000000001011111100000100",
			421 => "11111111100000010000011011111101",
			422 => "0000000010000000000011000000000100",
			423 => "00000000010100000000011011111101",
			424 => "00000000000000000000011011111101",
			425 => "0000000100000000001101101100001000",
			426 => "0000000011000000001001100000000100",
			427 => "00000000000000000000011011111101",
			428 => "11111110111111000000011011111101",
			429 => "00000000000000000000011011111101",
			430 => "0000001101000000000010011100011100",
			431 => "0000001001000000001001111100000100",
			432 => "00000000000000000000011011111101",
			433 => "0000000010000000001010000100001100",
			434 => "0000001110000000000110010000000100",
			435 => "00000000000000000000011011111101",
			436 => "0000001000000000001010110000000100",
			437 => "00000000000000000000011011111101",
			438 => "11111111110010110000011011111101",
			439 => "0000001110000000001011111000001000",
			440 => "0000000000000000000110001000000100",
			441 => "00000000000000000000011011111101",
			442 => "00000000110010000000011011111101",
			443 => "00000000000000000000011011111101",
			444 => "0000001110000000001111010100000100",
			445 => "00000000000000000000011011111101",
			446 => "11111111111100000000011011111101",
			447 => "0000001001000000001001111100000100",
			448 => "00000000000000000000011100111001",
			449 => "0000001101000000000111111100011000",
			450 => "0000001100000000001010111000000100",
			451 => "00000000000000000000011100111001",
			452 => "0000000110000000000100111100010000",
			453 => "0000001110000000001011111000001100",
			454 => "0000001100000000001000000000001000",
			455 => "0000001001000000000111101100000100",
			456 => "00000000000000000000011100111001",
			457 => "00000000011111110000011100111001",
			458 => "00000000000000000000011100111001",
			459 => "00000000000000000000011100111001",
			460 => "00000000000000000000011100111001",
			461 => "00000000000000000000011100111001",
			462 => "0000000001000000000001000100000100",
			463 => "00000000000000000000011101110101",
			464 => "0000001011000000000101100100011000",
			465 => "0000001010000000001010100100000100",
			466 => "00000000000000000000011101110101",
			467 => "0000001100000000001011000000010000",
			468 => "0000000111000000000001101000001100",
			469 => "0000001001000000001010100100001000",
			470 => "0000001110000000001011111000000100",
			471 => "00000000100001000000011101110101",
			472 => "00000000000000000000011101110101",
			473 => "00000000000000000000011101110101",
			474 => "00000000000000000000011101110101",
			475 => "00000000000000000000011101110101",
			476 => "00000000000000000000011101110101",
			477 => "0000000001000000001011111100001000",
			478 => "0000001001000000001001111100000100",
			479 => "11111110011110110000011111100001",
			480 => "00000000000000000000011111100001",
			481 => "0000001110000000000110111100010000",
			482 => "0000000100000000001111100100001000",
			483 => "0000001110000000000110010000000100",
			484 => "00000000110001010000011111100001",
			485 => "11111110101101000000011111100001",
			486 => "0000001100000000001011000000000100",
			487 => "00000001011100010000011111100001",
			488 => "00000000000000000000011111100001",
			489 => "0000001001000000000000001000001000",
			490 => "0000001101000000001110101000000100",
			491 => "00000000000000000000011111100001",
			492 => "11111110010111110000011111100001",
			493 => "0000001101000000000101001000001000",
			494 => "0000000000000000000111000000000100",
			495 => "00000001000110100000011111100001",
			496 => "00000000000000000000011111100001",
			497 => "0000001001000000001010100000001000",
			498 => "0000001011000000000110110100000100",
			499 => "00000000000000000000011111100001",
			500 => "00000000001111110000011111100001",
			501 => "0000001011000000000000011100000100",
			502 => "00000000000000000000011111100001",
			503 => "11111110111110010000011111100001",
			504 => "0000001100000000001010111000010000",
			505 => "0000000000000000000111000100000100",
			506 => "00000000000000000000100001011101",
			507 => "0000001001000000000000001000001000",
			508 => "0000000111000000001001001000000100",
			509 => "11111110011010100000100001011101",
			510 => "00000000000000000000100001011101",
			511 => "00000000000000000000100001011101",
			512 => "0000000111000000000110100100010100",
			513 => "0000001101000000000101001000010000",
			514 => "0000000010000000001100000000000100",
			515 => "00000000000000000000100001011101",
			516 => "0000001001000000000100101100000100",
			517 => "00000000000000000000100001011101",
			518 => "0000001110000000001011111000000100",
			519 => "00000000111110000000100001011101",
			520 => "00000000000000000000100001011101",
			521 => "00000000000000000000100001011101",
			522 => "0000000111000000001000011000001100",
			523 => "0000001110000000001100010000000100",
			524 => "00000000000000000000100001011101",
			525 => "0000001011000000000110110100000100",
			526 => "11111111000101000000100001011101",
			527 => "00000000000000000000100001011101",
			528 => "0000000101000000001110000100001100",
			529 => "0000001111000000001100111000001000",
			530 => "0000000010000000001010000100000100",
			531 => "00000000000000000000100001011101",
			532 => "00000000001011000000100001011101",
			533 => "00000000000000000000100001011101",
			534 => "00000000000000000000100001011101",
			535 => "0000001001000000000101010000000100",
			536 => "11111110101000110000100011000001",
			537 => "0000000100000000000010010100100000",
			538 => "0000001110000000000110111100010100",
			539 => "0000000100000000001111100100001000",
			540 => "0000001110000000000010000000000100",
			541 => "00000000010000000000100011000001",
			542 => "11111111010001110000100011000001",
			543 => "0000001100000000001011000000000100",
			544 => "00000001000101010000100011000001",
			545 => "0000000000000000001111001000000100",
			546 => "00000000010001000000100011000001",
			547 => "11111111100111000000100011000001",
			548 => "0000001111000000000000010000000100",
			549 => "00000000000000000000100011000001",
			550 => "0000000100000000000010010100000100",
			551 => "11111110110000110000100011000001",
			552 => "00000000000000000000100011000001",
			553 => "0000001110000000001011111000001100",
			554 => "0000001101000000000010011100001000",
			555 => "0000000110000000001000010000000100",
			556 => "00000001011111000000100011000001",
			557 => "00000000000000000000100011000001",
			558 => "00000000000000000000100011000001",
			559 => "11111111101010010000100011000001",
			560 => "0000000001000000000001000100000100",
			561 => "11111110011000110000100100000101",
			562 => "0000001110000000001011111000011100",
			563 => "0000001000000000000001110000011000",
			564 => "0000001101000000001001010000010000",
			565 => "0000001010000000001010100100000100",
			566 => "11111101101010100000100100000101",
			567 => "0000000000000000000111000000001000",
			568 => "0000001100000000001011000000000100",
			569 => "00000001110011010000100100000101",
			570 => "00000000101000010000100100000101",
			571 => "00000011110110010000100100000101",
			572 => "0000000010000000001111100100000100",
			573 => "11111110100001100000100100000101",
			574 => "00000010011011110000100100000101",
			575 => "11111101111100000000100100000101",
			576 => "11111110011001010000100100000101",
			577 => "0000001000000000000001110000101100",
			578 => "0000000011000000001011111000100100",
			579 => "0000000100000000001100111000010100",
			580 => "0000001110000000000110010000001000",
			581 => "0000000001000000001011111100000100",
			582 => "00000000000000000000100101100001",
			583 => "00000000101011110000100101100001",
			584 => "0000001011000000001011011100001000",
			585 => "0000001011000000000111010000000100",
			586 => "00000000000000000000100101100001",
			587 => "11111111001000010000100101100001",
			588 => "00000000000000000000100101100001",
			589 => "0000000001000000000001000100000100",
			590 => "00000000000000000000100101100001",
			591 => "0000000110000000000100111100001000",
			592 => "0000001000000000001010110000000100",
			593 => "00000000000000000000100101100001",
			594 => "00000001010110110000100101100001",
			595 => "00000000000000000000100101100001",
			596 => "0000000001000000000100110100000100",
			597 => "11111111000100110000100101100001",
			598 => "00000000000000000000100101100001",
			599 => "11111110101100000000100101100001",
			600 => "0000001000000000000001110000101100",
			601 => "0000000011000000001011111000100100",
			602 => "0000000100000000001100111000010000",
			603 => "0000001110000000000110010000001000",
			604 => "0000000001000000001011111100000100",
			605 => "00000000000000000000100110111101",
			606 => "00000000101001100000100110111101",
			607 => "0000000000000000000110001000000100",
			608 => "11111111001101010000100110111101",
			609 => "00000000000000000000100110111101",
			610 => "0000000001000000000001000100000100",
			611 => "00000000000000000000100110111101",
			612 => "0000000110000000000100111100001100",
			613 => "0000001000000000001010110000000100",
			614 => "00000000000000000000100110111101",
			615 => "0000001101000000000010011100000100",
			616 => "00000001010101010000100110111101",
			617 => "00000000000000000000100110111101",
			618 => "00000000000000000000100110111101",
			619 => "0000000001000000000100110100000100",
			620 => "11111111001000000000100110111101",
			621 => "00000000000000000000100110111101",
			622 => "11111110101101110000100110111101",
			623 => "0000001100000000001010111000100100",
			624 => "0000000010000000001000001100010100",
			625 => "0000001010000000000111110100010000",
			626 => "0000001011000000001010001100000100",
			627 => "00000000000000000000101001001001",
			628 => "0000000111000000001000000000000100",
			629 => "00000000000000000000101001001001",
			630 => "0000001011000000000000011100000100",
			631 => "11111111110010110000101001001001",
			632 => "00000000000000000000101001001001",
			633 => "11111110100010010000101001001001",
			634 => "0000001110000000001010000100001100",
			635 => "0000001011000000001001001000000100",
			636 => "00000000000000000000101001001001",
			637 => "0000000010000000001100111000000100",
			638 => "00000000001000110000101001001001",
			639 => "00000000000000000000101001001001",
			640 => "00000000000000000000101001001001",
			641 => "0000001001000000000111101100001100",
			642 => "0000001100000000000100011000000100",
			643 => "00000000000000000000101001001001",
			644 => "0000001100000000001000000000000100",
			645 => "11111111011000110000101001001001",
			646 => "00000000000000000000101001001001",
			647 => "0000000010000000001111010100000100",
			648 => "00000000000000000000101001001001",
			649 => "0000001110000000001111010100000100",
			650 => "00000000111001010000101001001001",
			651 => "0000000100000000001011110000000100",
			652 => "11111111110100110000101001001001",
			653 => "0000000111000000000001101000001000",
			654 => "0000000100000000000101000000000100",
			655 => "00000000010000010000101001001001",
			656 => "00000000000000000000101001001001",
			657 => "00000000000000000000101001001001",
			658 => "0000000001000000001011111100000100",
			659 => "11111110011001010000101010010101",
			660 => "0000000011000000001111100100100000",
			661 => "0000001110000000000110010000000100",
			662 => "00000001101110100000101010010101",
			663 => "0000001010000000000011101000001000",
			664 => "0000000111000000001001001000000100",
			665 => "00000000000000000000101010010101",
			666 => "11111101101100000000101010010101",
			667 => "0000000001000000000111101000001000",
			668 => "0000000110000000001001100100000100",
			669 => "00000000100001110000101010010101",
			670 => "11111101111111010000101010010101",
			671 => "0000001001000000001010100100001000",
			672 => "0000000000000000000110001000000100",
			673 => "11111111101101110000101010010101",
			674 => "00000001100100000000101010010101",
			675 => "11111110010011100000101010010101",
			676 => "11111110011010000000101010010101",
			677 => "0000000001000000000001000100000100",
			678 => "11111110011010000000101100011001",
			679 => "0000001110000000000110111100100000",
			680 => "0000001011000000000100000100001100",
			681 => "0000000100000000001011101100001000",
			682 => "0000001110000000000110010000000100",
			683 => "00000001100100000000101100011001",
			684 => "11111110110010010000101100011001",
			685 => "00000001101110000000101100011001",
			686 => "0000000100000000000001011100001100",
			687 => "0000001110000000000110010000000100",
			688 => "00000001001000010000101100011001",
			689 => "0000000101000000000110100000000100",
			690 => "11111111100100010000101100011001",
			691 => "11111110000111010000101100011001",
			692 => "0000000010000000000110101100000100",
			693 => "00000001100101010000101100011001",
			694 => "00000000000000000000101100011001",
			695 => "0000000111000000000110100100001100",
			696 => "0000000100000000000010010100000100",
			697 => "11111110100011100000101100011001",
			698 => "0000001110000000001011111000000100",
			699 => "00000001101001000000101100011001",
			700 => "11111111001001110000101100011001",
			701 => "0000000100000000000011000000001000",
			702 => "0000001000000000000110011100000100",
			703 => "11111110100111000000101100011001",
			704 => "11111011011100010000101100011001",
			705 => "0000001111000000001100111000001000",
			706 => "0000000100000000000010010100000100",
			707 => "11111111011011110000101100011001",
			708 => "00000001100010000000101100011001",
			709 => "11111110011110000000101100011001",
			710 => "0000001001000000000101010000001100",
			711 => "0000001001000000000101010000000100",
			712 => "11111110010111110000101110001101",
			713 => "0000001001000000000101010000000100",
			714 => "00000000000000000000101110001101",
			715 => "11111110101101110000101110001101",
			716 => "0000001101000000001001010000100100",
			717 => "0000001000000000000001110000100000",
			718 => "0000000010000000001101101100011100",
			719 => "0000001101000000000101001000010000",
			720 => "0000001100000000000100011000001000",
			721 => "0000000010000000001100111000000100",
			722 => "00000010100010100000101110001101",
			723 => "00000011110000010000101110001101",
			724 => "0000000010000000000111010100000100",
			725 => "00000000011110100000101110001101",
			726 => "00000010001111000000101110001101",
			727 => "0000001010000000000011101000000100",
			728 => "11111110011000110000101110001101",
			729 => "0000001110000000000111010100000100",
			730 => "00000010111111110000101110001101",
			731 => "11111110101000010000101110001101",
			732 => "00000101110011110000101110001101",
			733 => "11111110010001100000101110001101",
			734 => "0000001110000000001111010100001000",
			735 => "0000001001000000000100101100000100",
			736 => "11111110010111110000101110001101",
			737 => "00000001100100100000101110001101",
			738 => "11111110011000000000101110001101",
			739 => "0000001001000000001001111100010100",
			740 => "0000000001000000000001000100000100",
			741 => "11111110011100100000110000110001",
			742 => "0000001000000000000001010100001100",
			743 => "0000001000000000001010110000001000",
			744 => "0000000001000000001011111100000100",
			745 => "11111111110010110000110000110001",
			746 => "00000000000000000000110000110001",
			747 => "00000000010100110000110000110001",
			748 => "11111110111010000000110000110001",
			749 => "0000000111000000000001101000100100",
			750 => "0000000011000000001011111000011000",
			751 => "0000001100000000001011000000010000",
			752 => "0000000001000000001101111100001000",
			753 => "0000001110000000001000001100000100",
			754 => "00000001011010100000110000110001",
			755 => "00000000000000000000110000110001",
			756 => "0000000001000000000100110100000100",
			757 => "11111111101110110000110000110001",
			758 => "00000000100010110000110000110001",
			759 => "0000000001000000000001111000000100",
			760 => "11111111011001000000110000110001",
			761 => "00000000000000000000110000110001",
			762 => "0000000001000000000100110100000100",
			763 => "11111110101010010000110000110001",
			764 => "0000000101000000001110101000000100",
			765 => "00000000100111000000110000110001",
			766 => "00000000000000000000110000110001",
			767 => "0000001000000000000110011100001000",
			768 => "0000000011000000001010000100000100",
			769 => "00000000100110000000110000110001",
			770 => "00000000000000000000110000110001",
			771 => "0000001100000000001010111000000100",
			772 => "00000000000000000000110000110001",
			773 => "0000000100000000000101000000000100",
			774 => "11111110010000110000110000110001",
			775 => "0000000001000000000001111000001000",
			776 => "0000000001000000000001111000000100",
			777 => "00000000000000000000110000110001",
			778 => "00000000000011000000110000110001",
			779 => "11111111010000100000110000110001",
			780 => "0000000001000000000001000100000100",
			781 => "11111110011011000000110010010101",
			782 => "0000001110000000000110010000001000",
			783 => "0000000110000000001010011000000100",
			784 => "00000000000000000000110010010101",
			785 => "00000001100101000000110010010101",
			786 => "0000000100000000001100111000010100",
			787 => "0000000100000000000110101100000100",
			788 => "11111110000111010000110010010101",
			789 => "0000000011000000001100000000000100",
			790 => "00000000011101010000110010010101",
			791 => "0000000110000000001001100100001000",
			792 => "0000000110000000001011001100000100",
			793 => "00000000000000000000110010010101",
			794 => "11111110011000000000110010010101",
			795 => "00000000000000000000110010010101",
			796 => "0000001110000000001011111000010000",
			797 => "0000000001000000000111101000000100",
			798 => "11111110110100110000110010010101",
			799 => "0000000100000000000010010100001000",
			800 => "0000001110000000001111010100000100",
			801 => "00000001010101110000110010010101",
			802 => "11111110100011100000110010010101",
			803 => "00000001110110000000110010010101",
			804 => "11111110100110000000110010010101",
			805 => "0000000001000000000001000100000100",
			806 => "11111110100111100000110100011001",
			807 => "0000000111000000001001001000010100",
			808 => "0000000100000000001100111000001100",
			809 => "0000000000000000001011010100000100",
			810 => "00000000000100010000110100011001",
			811 => "0000001000000000001010110000000100",
			812 => "00000000000000000000110100011001",
			813 => "11111111011011000000110100011001",
			814 => "0000001110000000001000001100000100",
			815 => "00000001100000010000110100011001",
			816 => "00000000000000000000110100011001",
			817 => "0000001001000000000000001000010100",
			818 => "0000001110000000001100010000001100",
			819 => "0000000000000000001001101000000100",
			820 => "11111111010101000000110100011001",
			821 => "0000000000000000001111001000000100",
			822 => "00000000100111010000110100011001",
			823 => "00000000000000000000110100011001",
			824 => "0000001100000000001101010100000100",
			825 => "00000000000000000000110100011001",
			826 => "11111110111011010000110100011001",
			827 => "0000001100000000000100011000010000",
			828 => "0000000000000000001111001000000100",
			829 => "00000000000000000000110100011001",
			830 => "0000001000000000000001010100001000",
			831 => "0000001110000000001011111000000100",
			832 => "00000001000000010000110100011001",
			833 => "00000000000000000000110100011001",
			834 => "00000000000000000000110100011001",
			835 => "0000001000000000000110011100000100",
			836 => "00000000000000000000110100011001",
			837 => "11111111111010000000110100011001",
			838 => "0000001001000000001001111100001000",
			839 => "0000000100000000001100000000000100",
			840 => "00000000000000000000110110001101",
			841 => "11111110100100110000110110001101",
			842 => "0000000100000000000010010100100100",
			843 => "0000001101000000001100100100000100",
			844 => "00000001000000010000110110001101",
			845 => "0000001100000000001010111000000100",
			846 => "11111110110101000000110110001101",
			847 => "0000001000000000000110011100010000",
			848 => "0000001110000000000110111100001000",
			849 => "0000001000000000001010110000000100",
			850 => "00000000000000000000110110001101",
			851 => "00000001000100100000110110001101",
			852 => "0000000100000000000011000000000100",
			853 => "11111111100100010000110110001101",
			854 => "00000000000000000000110110001101",
			855 => "0000000000000000001111001000000100",
			856 => "00000000000000000000110110001101",
			857 => "0000001100000000000100011000000100",
			858 => "00000000000000000000110110001101",
			859 => "11111111000101010000110110001101",
			860 => "0000001101000000000111111100001100",
			861 => "0000000001000000000111101000000100",
			862 => "00000000000000000000110110001101",
			863 => "0000001110000000001011111000000100",
			864 => "00000001101100100000110110001101",
			865 => "00000000000000000000110110001101",
			866 => "11111111011101100000110110001101",
			867 => "0000001000000000000001010101000000",
			868 => "0000001101000000001111010000100000",
			869 => "0000000110000000001010011000000100",
			870 => "11111110011001100000111000110001",
			871 => "0000001100000000001011000000011000",
			872 => "0000000100000000000011000000010000",
			873 => "0000001110000000001100000000001000",
			874 => "0000000011000000001100010000000100",
			875 => "00000010000110010000111000110001",
			876 => "00000001101101110000111000110001",
			877 => "0000000010000000001000001100000100",
			878 => "11111111111111100000111000110001",
			879 => "11111110000101010000111000110001",
			880 => "0000000010000000001100111000000100",
			881 => "00000010000110000000111000110001",
			882 => "00000010110001010000111000110001",
			883 => "00000000100101100000111000110001",
			884 => "0000000101000000000110100000001000",
			885 => "0000000000000000000001010100000100",
			886 => "11111110111011010000111000110001",
			887 => "00000010110000010000111000110001",
			888 => "0000001100000000000100011000001100",
			889 => "0000000000000000000111000100000100",
			890 => "11111110011100110000111000110001",
			891 => "0000000110000000001111000000000100",
			892 => "00000010111011010000111000110001",
			893 => "11111111000000000000111000110001",
			894 => "0000000101000000001100100100001000",
			895 => "0000000101000000001110101000000100",
			896 => "11111110011100100000111000110001",
			897 => "00000000111000010000111000110001",
			898 => "11111110011001010000111000110001",
			899 => "0000001000000000000001110000010000",
			900 => "0000001110000000001000001100001100",
			901 => "0000001100000000000100001000000100",
			902 => "11111110011101010000111000110001",
			903 => "0000000100000000000010110000000100",
			904 => "00000001010100000000111000110001",
			905 => "00000010110101000000111000110001",
			906 => "11111110011010000000111000110001",
			907 => "11111110011000000000111000110001",
			908 => "0000000001000000000001000100000100",
			909 => "11111110100110010000111010111101",
			910 => "0000000111000000001001001000010100",
			911 => "0000000100000000001100111000001100",
			912 => "0000000000000000001011010100000100",
			913 => "00000000000101010000111010111101",
			914 => "0000001000000000001010110000000100",
			915 => "00000000000000000000111010111101",
			916 => "11111111010110010000111010111101",
			917 => "0000001110000000001000001100000100",
			918 => "00000001100010110000111010111101",
			919 => "00000000000000000000111010111101",
			920 => "0000001001000000000000001000011000",
			921 => "0000001110000000001100010000010000",
			922 => "0000000000000000001001101000000100",
			923 => "11111111010010110000111010111101",
			924 => "0000000000000000001111001000001000",
			925 => "0000000010000000001100000000000100",
			926 => "00000000000000000000111010111101",
			927 => "00000000110000000000111010111101",
			928 => "00000000000000000000111010111101",
			929 => "0000001100000000001101010100000100",
			930 => "00000000000000000000111010111101",
			931 => "11111110110111000000111010111101",
			932 => "0000001100000000000100011000010000",
			933 => "0000000000000000001111001000000100",
			934 => "00000000000000000000111010111101",
			935 => "0000001000000000000001010100001000",
			936 => "0000001110000000001011111000000100",
			937 => "00000001000010110000111010111101",
			938 => "00000000000000000000111010111101",
			939 => "00000000000000000000111010111101",
			940 => "0000001000000000000110011100000100",
			941 => "00000000000000000000111010111101",
			942 => "11111111111000010000111010111101",
			943 => "0000000001000000000001000100000100",
			944 => "11111110011001100000111100011001",
			945 => "0000000011000000001011101100101000",
			946 => "0000000011000000001100010000000100",
			947 => "00000001101100000000111100011001",
			948 => "0000000100000000001011101100001100",
			949 => "0000001111000000000110111100001000",
			950 => "0000000010000000001100000000000100",
			951 => "11111110111010100000111100011001",
			952 => "00000000000000000000111100011001",
			953 => "11111101101011100000111100011001",
			954 => "0000000001000000000111101000001000",
			955 => "0000000101000000000010110100000100",
			956 => "00000000000000000000111100011001",
			957 => "11111110011000010000111100011001",
			958 => "0000000100000000000011000000001000",
			959 => "0000000110000000001001100100000100",
			960 => "00000000110111010000111100011001",
			961 => "11111101001000010000111100011001",
			962 => "0000000110000000001000010000000100",
			963 => "00000001110100010000111100011001",
			964 => "11111111001110000000111100011001",
			965 => "11111110011011110000111100011001",
			966 => "0000000001000000000001000100000100",
			967 => "11111110011010110000111110001101",
			968 => "0000001110000000000110010000001000",
			969 => "0000000110000000001010011000000100",
			970 => "00000000000000000000111110001101",
			971 => "00000001100110010000111110001101",
			972 => "0000000100000000001100111000011000",
			973 => "0000000100000000001111100100000100",
			974 => "11111110001100110000111110001101",
			975 => "0000000011000000001100000000001000",
			976 => "0000001001000000000000001000000100",
			977 => "00000000000000000000111110001101",
			978 => "00000000110001010000111110001101",
			979 => "0000000110000000001001100100001000",
			980 => "0000000110000000001011001100000100",
			981 => "00000000000000000000111110001101",
			982 => "11111110011100110000111110001101",
			983 => "00000000000000000000111110001101",
			984 => "0000001110000000001011111000010100",
			985 => "0000000001000000000111101000000100",
			986 => "11111110110000100000111110001101",
			987 => "0000000100000000000010010100001000",
			988 => "0000001110000000001111010100000100",
			989 => "00000001011000000000111110001101",
			990 => "11111110100000100000111110001101",
			991 => "0000000110000000000100111100000100",
			992 => "00000001111100100000111110001101",
			993 => "00000000000000000000111110001101",
			994 => "11111110100100100000111110001101",
			995 => "0000000001000000000001000100000100",
			996 => "11111110011010010001000000100001",
			997 => "0000000111000000001001001000011100",
			998 => "0000000100000000000011001100010100",
			999 => "0000000011000000001100010000000100",
			1000 => "00000001100101110001000000100001",
			1001 => "0000000100000000001011101100000100",
			1002 => "11111110010001100001000000100001",
			1003 => "0000001110000000001011111000001000",
			1004 => "0000000100000000001101101100000100",
			1005 => "00000000000000000001000000100001",
			1006 => "00000001100001010001000000100001",
			1007 => "11111111101111100001000000100001",
			1008 => "0000000100000000001010110100000100",
			1009 => "00000100011111010001000000100001",
			1010 => "00000000000000000001000000100001",
			1011 => "0000001110000000000110111100010100",
			1012 => "0000001010000000000011101000001000",
			1013 => "0000000011000000001100010000000100",
			1014 => "00000000010111100001000000100001",
			1015 => "11111110010111100001000000100001",
			1016 => "0000001001000000000100101100000100",
			1017 => "11111111000000110001000000100001",
			1018 => "0000000010000000000111011000000100",
			1019 => "00000000000100110001000000100001",
			1020 => "00000001100111110001000000100001",
			1021 => "0000000011000000000111010100000100",
			1022 => "11111101100010010001000000100001",
			1023 => "0000000101000000001100100100010000",
			1024 => "0000000111000000000110100100001000",
			1025 => "0000000011000000001111100100000100",
			1026 => "00000000100101000001000000100001",
			1027 => "00000000000000000001000000100001",
			1028 => "0000001011000000001011011100000100",
			1029 => "11111111010000010001000000100001",
			1030 => "00000000000000000001000000100001",
			1031 => "11111110100011000001000000100001",
			1032 => "0000000001000000000001000100000100",
			1033 => "11111110011011110001000010101101",
			1034 => "0000001110000000000110010000001000",
			1035 => "0000000110000000001010011000000100",
			1036 => "00000000000000000001000010101101",
			1037 => "00000001100010100001000010101101",
			1038 => "0000000001000000000111101000010000",
			1039 => "0000001001000000000111101100001100",
			1040 => "0000000111000000000110100100000100",
			1041 => "11111110100000010001000010101101",
			1042 => "0000001100000000000100011000000100",
			1043 => "00000000000000000001000010101101",
			1044 => "11111111011001100001000010101101",
			1045 => "00000000000000000001000010101101",
			1046 => "0000000111000000000001101000010100",
			1047 => "0000000100000000000010010100001100",
			1048 => "0000001110000000000110111100001000",
			1049 => "0000000100000000001111100100000100",
			1050 => "11111110111001100001000010101101",
			1051 => "00000001001101010001000010101101",
			1052 => "11111110100001110001000010101101",
			1053 => "0000001110000000001011111000000100",
			1054 => "00000001101111100001000010101101",
			1055 => "11111111100100100001000010101101",
			1056 => "0000001100000000000100011000001100",
			1057 => "0000000000000000001111001000000100",
			1058 => "00000000000000000001000010101101",
			1059 => "0000001001000000001010100100000100",
			1060 => "00000001000010010001000010101101",
			1061 => "00000000000000000001000010101101",
			1062 => "0000001000000000001100011100000100",
			1063 => "00000000000000000001000010101101",
			1064 => "0000000100000000000101000000000100",
			1065 => "11111110000011010001000010101101",
			1066 => "11111111100010110001000010101101",
			1067 => "0000000001000000000001000100000100",
			1068 => "11111110011000110001000100100011",
			1069 => "0000001110000000001011111000110100",
			1070 => "0000001000000000000001110000110000",
			1071 => "0000000100000000000001011100011100",
			1072 => "0000001110000000001110110100001100",
			1073 => "0000000001000000001011111100000100",
			1074 => "11111101100110010001000100100011",
			1075 => "0000000001000000001101111100000100",
			1076 => "00000001110110100001000100100011",
			1077 => "00000000111001000001000100100011",
			1078 => "0000000100000000001011101100001000",
			1079 => "0000001010000000000011101000000100",
			1080 => "11111110100100100001000100100011",
			1081 => "11111100111001010001000100100011",
			1082 => "0000001100000000000100011000000100",
			1083 => "00000001001101110001000100100011",
			1084 => "11111101100010110001000100100011",
			1085 => "0000000010000000001101101100010000",
			1086 => "0000001101000000001111010000001000",
			1087 => "0000001111000000001111100100000100",
			1088 => "00000001111001100001000100100011",
			1089 => "00000001010000100001000100100011",
			1090 => "0000001111000000001111100100000100",
			1091 => "00000000000101110001000100100011",
			1092 => "11111111000011000001000100100011",
			1093 => "00000011101111110001000100100011",
			1094 => "11111101111111010001000100100011",
			1095 => "11111110011001100001000100100011",
			1096 => "00000000000000000001000100100101",
			1097 => "00000000000000000001000100101001",
			1098 => "00000000000000000001000100101101",
			1099 => "00000000000000000001000100110001",
			1100 => "00000000000000000001000100110101",
			1101 => "00000000000000000001000100111001",
			1102 => "00000000000000000001000100111101",
			1103 => "00000000000000000001000101000001",
			1104 => "00000000000000000001000101000101",
			1105 => "00000000000000000001000101001001",
			1106 => "00000000000000000001000101001101",
			1107 => "00000000000000000001000101010001",
			1108 => "00000000000000000001000101010101",
			1109 => "00000000000000000001000101011001",
			1110 => "00000000000000000001000101011101",
			1111 => "00000000000000000001000101100001",
			1112 => "00000000000000000001000101100101",
			1113 => "00000000000000000001000101101001",
			1114 => "00000000000000000001000101101101",
			1115 => "00000000000000000001000101110001",
			1116 => "00000000000000000001000101110101",
			1117 => "00000000000000000001000101111001",
			1118 => "00000000000000000001000101111101",
			1119 => "00000000000000000001000110000001",
			1120 => "00000000000000000001000110000101",
			1121 => "00000000000000000001000110001001",
			1122 => "00000000000000000001000110001101",
			1123 => "0000001000000000000001010100000100",
			1124 => "00000000000000000001000110011001",
			1125 => "11111111101101110001000110011001",
			1126 => "0000001000000000001100011100000100",
			1127 => "00000000000000000001000110100101",
			1128 => "11111111111011010001000110100101",
			1129 => "0000000001000000001101111100000100",
			1130 => "11111111111110010001000110110001",
			1131 => "00000000000000000001000110110001",
			1132 => "0000001110000000000110010000001000",
			1133 => "0000001110000000000101001000000100",
			1134 => "00000000000000000001000111000101",
			1135 => "00000000001010110001000111000101",
			1136 => "11111111111101010001000111000101",
			1137 => "0000001000000000000001010100001000",
			1138 => "0000000100000000000011000000000100",
			1139 => "00000000000000000001000111011001",
			1140 => "00000000001001010001000111011001",
			1141 => "11111111101011000001000111011001",
			1142 => "0000001110000000001100000000000100",
			1143 => "00000000000000000001000111101101",
			1144 => "0000001111000000001000001100000100",
			1145 => "00000000000000000001000111101101",
			1146 => "11111111111110000001000111101101",
			1147 => "0000000001000000001011111100000100",
			1148 => "11111111110001000001001000001001",
			1149 => "0000000001000000001100011000001000",
			1150 => "0000000001000000001110010100000100",
			1151 => "00000000000000000001001000001001",
			1152 => "00000000000010010001001000001001",
			1153 => "00000000000000000001001000001001",
			1154 => "0000001000000000000001010100001100",
			1155 => "0000000001000000001011111100000100",
			1156 => "00000000000000000001001000100101",
			1157 => "0000001001000000001010100100000100",
			1158 => "00000000001110000001001000100101",
			1159 => "00000000000000000001001000100101",
			1160 => "00000000000000000001001000100101",
			1161 => "0000000001000000000111101000001000",
			1162 => "0000001001000000000111101100000100",
			1163 => "11111111111000010001001001001001",
			1164 => "00000000000000000001001001001001",
			1165 => "0000000010000000001010000100000100",
			1166 => "00000000000000000001001001001001",
			1167 => "0000000010000000001111101000000100",
			1168 => "00000000000111000001001001001001",
			1169 => "00000000000000000001001001001001",
			1170 => "0000001110000000000110010000001100",
			1171 => "0000001001000000000101010000000100",
			1172 => "00000000000000000001001001110101",
			1173 => "0000000000000000001100000100000100",
			1174 => "00000000000000000001001001110101",
			1175 => "00000000001101010001001001110101",
			1176 => "0000000001000000000100110100001000",
			1177 => "0000001100000000000100001000000100",
			1178 => "00000000000000000001001001110101",
			1179 => "11111111101011010001001001110101",
			1180 => "00000000000000000001001001110101",
			1181 => "0000001001000000001001111100000100",
			1182 => "11111111101010010001001010011001",
			1183 => "0000000110000000000100111100001100",
			1184 => "0000000110000000001010011000000100",
			1185 => "00000000000000000001001010011001",
			1186 => "0000001001000000001010100100000100",
			1187 => "00000000001100000001001010011001",
			1188 => "00000000000000000001001010011001",
			1189 => "00000000000000000001001010011001",
			1190 => "0000000001000000001110010100000100",
			1191 => "00000000000000000001001010111101",
			1192 => "0000001001000000001010100100001100",
			1193 => "0000001000000000000001110000001000",
			1194 => "0000001000000000001010110000000100",
			1195 => "00000000000000000001001010111101",
			1196 => "00000000001001100001001010111101",
			1197 => "00000000000000000001001010111101",
			1198 => "00000000000000000001001010111101",
			1199 => "0000001001000000000000001000010000",
			1200 => "0000001110000000000110010000000100",
			1201 => "00000000000000000001001011100001",
			1202 => "0000000100000000000011110000001000",
			1203 => "0000000011000000001100010000000100",
			1204 => "00000000000000000001001011100001",
			1205 => "11111111110010000001001011100001",
			1206 => "00000000000000000001001011100001",
			1207 => "00000000000000000001001011100001",
			1208 => "0000001001000000000111101100001000",
			1209 => "0000001011000000000100000100000100",
			1210 => "00000000000000000001001100001101",
			1211 => "11111111101010000001001100001101",
			1212 => "0000001100000000001010111000000100",
			1213 => "00000000000000000001001100001101",
			1214 => "0000001101000000001111010000001000",
			1215 => "0000001010000000001000010100000100",
			1216 => "00000000011110000001001100001101",
			1217 => "00000000000000000001001100001101",
			1218 => "00000000000000000001001100001101",
			1219 => "0000001110000000000110010000010000",
			1220 => "0000001110000000000101001000000100",
			1221 => "00000000000000000001001101000001",
			1222 => "0000001101000000000001000000001000",
			1223 => "0000000010000000001011101100000100",
			1224 => "00000000010000000001001101000001",
			1225 => "00000000000000000001001101000001",
			1226 => "00000000000000000001001101000001",
			1227 => "0000000100000000000011000000001000",
			1228 => "0000001101000000001110101000000100",
			1229 => "00000000000000000001001101000001",
			1230 => "11111111101101100001001101000001",
			1231 => "00000000000000000001001101000001",
			1232 => "0000001001000000001001111100000100",
			1233 => "11111111101011110001001101101101",
			1234 => "0000000110000000000100111100010000",
			1235 => "0000000110000000001010011000000100",
			1236 => "00000000000000000001001101101101",
			1237 => "0000001001000000001010100100001000",
			1238 => "0000000001000000001110010100000100",
			1239 => "00000000000000000001001101101101",
			1240 => "00000000001010110001001101101101",
			1241 => "00000000000000000001001101101101",
			1242 => "00000000000000000001001101101101",
			1243 => "0000001001000000000111101100001100",
			1244 => "0000001000000000001010110000000100",
			1245 => "00000000000000000001001110101001",
			1246 => "0000001100000000001010111100000100",
			1247 => "11111111111000100001001110101001",
			1248 => "00000000000000000001001110101001",
			1249 => "0000001000000000000101000100010000",
			1250 => "0000001100000000001010111000000100",
			1251 => "00000000000000000001001110101001",
			1252 => "0000001001000000001010100100001000",
			1253 => "0000001100000000001011000000000100",
			1254 => "00000000011010000001001110101001",
			1255 => "00000000000000000001001110101001",
			1256 => "00000000000000000001001110101001",
			1257 => "00000000000000000001001110101001",
			1258 => "0000001001000000001001111100001000",
			1259 => "0000000100000000001100010000000100",
			1260 => "00000000000000000001001111101101",
			1261 => "11111111101001100001001111101101",
			1262 => "0000001110000000001100000000010000",
			1263 => "0000000100000000001111100100000100",
			1264 => "00000000000000000001001111101101",
			1265 => "0000001010000000000011101000000100",
			1266 => "00000000000000000001001111101101",
			1267 => "0000001010000000000111110100000100",
			1268 => "00000000101001000001001111101101",
			1269 => "00000000000000000001001111101101",
			1270 => "0000000100000000001111101000001000",
			1271 => "0000001111000000001000001100000100",
			1272 => "00000000000000000001001111101101",
			1273 => "11111111100010000001001111101101",
			1274 => "00000000000000000001001111101101",
			1275 => "0000000010000000001000001100011100",
			1276 => "0000001110000000000110010000001100",
			1277 => "0000000001000000001011111100001000",
			1278 => "0000000010000000000111011000000100",
			1279 => "11111111101110010001010001001001",
			1280 => "00000000000000000001010001001001",
			1281 => "00000000010111100001010001001001",
			1282 => "0000000100000000001101101100001100",
			1283 => "0000001011000000000101100100001000",
			1284 => "0000001100000000001000000000000100",
			1285 => "11111111001010000001010001001001",
			1286 => "00000000000000000001010001001001",
			1287 => "00000000000000000001010001001001",
			1288 => "00000000000000000001010001001001",
			1289 => "0000001110000000000111010100001100",
			1290 => "0000001001000000000101010000000100",
			1291 => "00000000000000000001010001001001",
			1292 => "0000000100000000001000101000000100",
			1293 => "00000000000000000001010001001001",
			1294 => "00000000101101110001010001001001",
			1295 => "0000000001000000001101111100000100",
			1296 => "11111111110001010001010001001001",
			1297 => "00000000000000000001010001001001",
			1298 => "0000001001000000001001111100001000",
			1299 => "0000000110000000001001100100000100",
			1300 => "11111111010000110001010010010101",
			1301 => "00000000000000000001010010010101",
			1302 => "0000001110000000001100000000010000",
			1303 => "0000000001000000001101111100001100",
			1304 => "0000000101000000000110100000001000",
			1305 => "0000001110000000001100010000000100",
			1306 => "00000000110011100001010010010101",
			1307 => "00000000000000000001010010010101",
			1308 => "00000000000000000001010010010101",
			1309 => "00000000000000000001010010010101",
			1310 => "0000000001000000001101111100001100",
			1311 => "0000001010000000001000100100001000",
			1312 => "0000001111000000000111010100000100",
			1313 => "00000000000000000001010010010101",
			1314 => "11111111010001000001010010010101",
			1315 => "00000000000000000001010010010101",
			1316 => "00000000000000000001010010010101",
			1317 => "0000001100000000001010111100000100",
			1318 => "00000000000000000001010011001001",
			1319 => "0000001101000000000010011100010100",
			1320 => "0000001010000000000011101000000100",
			1321 => "00000000000000000001010011001001",
			1322 => "0000000110000000000100111100001100",
			1323 => "0000000100000000001101101100000100",
			1324 => "00000000000000000001010011001001",
			1325 => "0000001001000000000101010000000100",
			1326 => "00000000000000000001010011001001",
			1327 => "00000000101100110001010011001001",
			1328 => "00000000000000000001010011001001",
			1329 => "00000000000000000001010011001001",
			1330 => "0000001100000000001010111000010000",
			1331 => "0000001110000000000110010000000100",
			1332 => "00000000000000000001010100010101",
			1333 => "0000001011000000001000011000000100",
			1334 => "00000000000000000001010100010101",
			1335 => "0000001101000000000101001000000100",
			1336 => "11111111110111000001010100010101",
			1337 => "00000000000000000001010100010101",
			1338 => "0000001101000000000010011100010100",
			1339 => "0000001100000000001011000000010000",
			1340 => "0000000110000000000100111100001100",
			1341 => "0000000001000000001011111100000100",
			1342 => "00000000000000000001010100010101",
			1343 => "0000001101000000001001010000000100",
			1344 => "00000000101000000001010100010101",
			1345 => "00000000000000000001010100010101",
			1346 => "00000000000000000001010100010101",
			1347 => "00000000000000000001010100010101",
			1348 => "00000000000000000001010100010101",
			1349 => "0000000010000000001010000100010000",
			1350 => "0000001110000000000110010000000100",
			1351 => "00000000000000000001010101110001",
			1352 => "0000000110000000001001100100001000",
			1353 => "0000001111000000001010000100000100",
			1354 => "11111111101001010001010101110001",
			1355 => "00000000000000000001010101110001",
			1356 => "00000000000000000001010101110001",
			1357 => "0000001111000000001000001100010000",
			1358 => "0000000100000000001011101100000100",
			1359 => "00000000000000000001010101110001",
			1360 => "0000001010000000001000010100001000",
			1361 => "0000000110000000001101011000000100",
			1362 => "00000000000000000001010101110001",
			1363 => "00000000100000100001010101110001",
			1364 => "00000000000000000001010101110001",
			1365 => "0000000100000000001000000100001100",
			1366 => "0000001110000000001100010000000100",
			1367 => "00000000000000000001010101110001",
			1368 => "0000001101000000001110101000000100",
			1369 => "00000000000000000001010101110001",
			1370 => "11111111101111000001010101110001",
			1371 => "00000000000000000001010101110001",
			1372 => "0000001100000000001010111000010000",
			1373 => "0000001010000000000111110100000100",
			1374 => "00000000000000000001010111010101",
			1375 => "0000000001000000001101111100001000",
			1376 => "0000000111000000001001001000000100",
			1377 => "11111110111000100001010111010101",
			1378 => "00000000000000000001010111010101",
			1379 => "00000000000000000001010111010101",
			1380 => "0000000111000000001001001000001100",
			1381 => "0000000010000000001100000000000100",
			1382 => "00000000000000000001010111010101",
			1383 => "0000001010000000001001000100000100",
			1384 => "00000000110100000001010111010101",
			1385 => "00000000000000000001010111010101",
			1386 => "0000001100000000000100011000001100",
			1387 => "0000001101000000000101001000001000",
			1388 => "0000000001000000001110010100000100",
			1389 => "00000000000000000001010111010101",
			1390 => "00000000010111010001010111010101",
			1391 => "00000000000000000001010111010101",
			1392 => "0000001000000000000110011100000100",
			1393 => "00000000000000000001010111010101",
			1394 => "0000000100000000000101000000000100",
			1395 => "11111111001110100001010111010101",
			1396 => "00000000000000000001010111010101",
			1397 => "0000001100000000001010111000011000",
			1398 => "0000001101000000001100100100001100",
			1399 => "0000001001000000000101010000000100",
			1400 => "11111111101010110001011001001001",
			1401 => "0000001110000000000110111100000100",
			1402 => "00000000100100010001011001001001",
			1403 => "00000000000000000001011001001001",
			1404 => "0000001011000000000100000100000100",
			1405 => "00000000000000000001011001001001",
			1406 => "0000000111000000001000000000000100",
			1407 => "00000000000000000001011001001001",
			1408 => "11111111001101110001011001001001",
			1409 => "0000000111000000000110100100001100",
			1410 => "0000001001000000000100101100000100",
			1411 => "00000000000000000001011001001001",
			1412 => "0000001110000000001011111000000100",
			1413 => "00000000101101000001011001001001",
			1414 => "00000000000000000001011001001001",
			1415 => "0000001000000000000101000100001100",
			1416 => "0000001000000000001010110000000100",
			1417 => "00000000000000000001011001001001",
			1418 => "0000001100000000001000000000000100",
			1419 => "00000000010110110001011001001001",
			1420 => "00000000000000000001011001001001",
			1421 => "0000001100000000001010111000000100",
			1422 => "00000000000000000001011001001001",
			1423 => "0000001001000000000000001000000100",
			1424 => "00000000000000000001011001001001",
			1425 => "11111111100101100001011001001001",
			1426 => "0000001100000000001010111000010000",
			1427 => "0000001010000000000111110100000100",
			1428 => "00000000000000000001011010110101",
			1429 => "0000000001000000001101111100001000",
			1430 => "0000000111000000001001001000000100",
			1431 => "11111110110101000001011010110101",
			1432 => "00000000000000000001011010110101",
			1433 => "00000000000000000001011010110101",
			1434 => "0000000111000000001001001000010000",
			1435 => "0000000010000000001100000000000100",
			1436 => "00000000000000000001011010110101",
			1437 => "0000001010000000001001000100001000",
			1438 => "0000000001000000001110010100000100",
			1439 => "00000000000000000001011010110101",
			1440 => "00000000110110100001011010110101",
			1441 => "00000000000000000001011010110101",
			1442 => "0000001100000000000100011000001100",
			1443 => "0000001101000000000101001000001000",
			1444 => "0000000001000000001110010100000100",
			1445 => "00000000000000000001011010110101",
			1446 => "00000000011000100001011010110101",
			1447 => "00000000000000000001011010110101",
			1448 => "0000001000000000000110011100000100",
			1449 => "00000000000000000001011010110101",
			1450 => "0000000100000000000101000000000100",
			1451 => "11111111001011010001011010110101",
			1452 => "00000000000000000001011010110101",
			1453 => "0000000010000000000110111100001100",
			1454 => "0000000110000000001001100100001000",
			1455 => "0000000100000000001100010000000100",
			1456 => "00000000000000000001011100000001",
			1457 => "11111111101110010001011100000001",
			1458 => "00000000000000000001011100000001",
			1459 => "0000000100000000000001011100000100",
			1460 => "00000000000000000001011100000001",
			1461 => "0000000110000000000100111100010100",
			1462 => "0000001100000000000100001000000100",
			1463 => "00000000000000000001011100000001",
			1464 => "0000001010000000000011101000000100",
			1465 => "00000000000000000001011100000001",
			1466 => "0000000010000000001111101000001000",
			1467 => "0000000001000000000001000100000100",
			1468 => "00000000000000000001011100000001",
			1469 => "00000000101001010001011100000001",
			1470 => "00000000000000000001011100000001",
			1471 => "00000000000000000001011100000001",
			1472 => "0000001111000000001000001100100000",
			1473 => "0000000111000000001110110000001100",
			1474 => "0000000001000000001011111100001000",
			1475 => "0000001101000000001110101100000100",
			1476 => "11111111100010000001011101101101",
			1477 => "00000000000000000001011101101101",
			1478 => "00000000000000000001011101101101",
			1479 => "0000000100000000001111100100001100",
			1480 => "0000000011000000001110110100000100",
			1481 => "00000000000000000001011101101101",
			1482 => "0000001110000000000110010000000100",
			1483 => "00000000000000000001011101101101",
			1484 => "11111111110010010001011101101101",
			1485 => "0000000001000000000001000100000100",
			1486 => "00000000000000000001011101101101",
			1487 => "00000000110011100001011101101101",
			1488 => "0000001100000000001011000000010100",
			1489 => "0000000001000000001101111100010000",
			1490 => "0000001110000000001100010000000100",
			1491 => "00000000000000000001011101101101",
			1492 => "0000001101000000001110101000000100",
			1493 => "00000000000000000001011101101101",
			1494 => "0000001001000000000000001000000100",
			1495 => "11111111001001010001011101101101",
			1496 => "00000000000000000001011101101101",
			1497 => "00000000000000000001011101101101",
			1498 => "00000000000000000001011101101101",
			1499 => "0000001000000000000001110000101000",
			1500 => "0000000100000000000011000000011000",
			1501 => "0000001110000000001100010000010000",
			1502 => "0000001010000000001010100100000100",
			1503 => "00000000000000000001011111000001",
			1504 => "0000001101000000001110000100001000",
			1505 => "0000000001000000001011111100000100",
			1506 => "00000000000000000001011111000001",
			1507 => "00000000101110110001011111000001",
			1508 => "00000000000000000001011111000001",
			1509 => "0000001001000000001010100000000100",
			1510 => "11111111000011010001011111000001",
			1511 => "00000000000000000001011111000001",
			1512 => "0000001101000000000111111100001100",
			1513 => "0000000001000000000001000100000100",
			1514 => "00000000000000000001011111000001",
			1515 => "0000001110000000001011111000000100",
			1516 => "00000000111010100001011111000001",
			1517 => "00000000000000000001011111000001",
			1518 => "00000000000000000001011111000001",
			1519 => "11111111011111000001011111000001",
			1520 => "0000001100000000001010111100001100",
			1521 => "0000000001000000000111101000001000",
			1522 => "0000001000000000000001010000000100",
			1523 => "00000000000000000001100000101101",
			1524 => "11111111100010100001100000101101",
			1525 => "00000000000000000001100000101101",
			1526 => "0000001110000000001110110100001100",
			1527 => "0000001010000000001010100000000100",
			1528 => "00000000000000000001100000101101",
			1529 => "0000001001000000000101010000000100",
			1530 => "00000000000000000001100000101101",
			1531 => "00000000101011000001100000101101",
			1532 => "0000000100000000000011000000010000",
			1533 => "0000001001000000001010100000001100",
			1534 => "0000001100000000000111001000000100",
			1535 => "00000000000000000001100000101101",
			1536 => "0000000001000000000001111000000100",
			1537 => "00000000000000000001100000101101",
			1538 => "11111111011101010001100000101101",
			1539 => "00000000000000000001100000101101",
			1540 => "0000000011000000001111100100001100",
			1541 => "0000000001000000000111101000000100",
			1542 => "00000000000000000001100000101101",
			1543 => "0000001100000000001010111000000100",
			1544 => "00000000000000000001100000101101",
			1545 => "00000000100001110001100000101101",
			1546 => "00000000000000000001100000101101",
			1547 => "0000001001000000001001111100000100",
			1548 => "00000000000000000001100001101001",
			1549 => "0000000101000000000001000000011000",
			1550 => "0000000000000000001001101000000100",
			1551 => "00000000000000000001100001101001",
			1552 => "0000000110000000000100111100010000",
			1553 => "0000001110000000001011111000001100",
			1554 => "0000000111000000000011100000000100",
			1555 => "00000000000000000001100001101001",
			1556 => "0000000111000000001000011000000100",
			1557 => "00000000010010110001100001101001",
			1558 => "00000000000000000001100001101001",
			1559 => "00000000000000000001100001101001",
			1560 => "00000000000000000001100001101001",
			1561 => "00000000000000000001100001101001",
			1562 => "0000001100000000001010111000011000",
			1563 => "0000000000000000000111000100010000",
			1564 => "0000001101000000001100100100000100",
			1565 => "00000000000000000001100011011101",
			1566 => "0000000101000000000010110100001000",
			1567 => "0000000101000000000010110100000100",
			1568 => "00000000000000000001100011011101",
			1569 => "11111111110100000001100011011101",
			1570 => "00000000000000000001100011011101",
			1571 => "0000000010000000001000001100000100",
			1572 => "11111111001010110001100011011101",
			1573 => "00000000000000000001100011011101",
			1574 => "0000001101000000000010011100011100",
			1575 => "0000001001000000001001111100000100",
			1576 => "00000000000000000001100011011101",
			1577 => "0000000010000000001010000100001100",
			1578 => "0000001110000000000110010000000100",
			1579 => "00000000000000000001100011011101",
			1580 => "0000000001000000000001111000000100",
			1581 => "00000000000000000001100011011101",
			1582 => "11111111110010110001100011011101",
			1583 => "0000001110000000001011111000001000",
			1584 => "0000000000000000000110001000000100",
			1585 => "00000000000000000001100011011101",
			1586 => "00000000101111100001100011011101",
			1587 => "00000000000000000001100011011101",
			1588 => "0000001110000000001111010100000100",
			1589 => "00000000000000000001100011011101",
			1590 => "11111111111111100001100011011101",
			1591 => "0000001001000000001001111100001100",
			1592 => "0000000110000000001001100100001000",
			1593 => "0000000100000000001100010000000100",
			1594 => "00000000000000000001100101001001",
			1595 => "11111111010010000001100101001001",
			1596 => "00000000000000000001100101001001",
			1597 => "0000001110000000001100000000010000",
			1598 => "0000000100000000001111100100000100",
			1599 => "00000000000000000001100101001001",
			1600 => "0000001000000000000110011100001000",
			1601 => "0000001000000000001010110000000100",
			1602 => "00000000000000000001100101001001",
			1603 => "00000000101001010001100101001001",
			1604 => "00000000000000000001100101001001",
			1605 => "0000000100000000000011000000001000",
			1606 => "0000001111000000000111010100000100",
			1607 => "00000000000000000001100101001001",
			1608 => "11111111001011000001100101001001",
			1609 => "0000001000000000000001010100010000",
			1610 => "0000000100000000000010010100000100",
			1611 => "00000000000000000001100101001001",
			1612 => "0000001101000000000111111100001000",
			1613 => "0000001111000000001000101000000100",
			1614 => "00000000100011000001100101001001",
			1615 => "00000000000000000001100101001001",
			1616 => "00000000000000000001100101001001",
			1617 => "00000000000000000001100101001001",
			1618 => "0000001100000000001010111000010000",
			1619 => "0000001010000000000111110100000100",
			1620 => "00000000000000000001100111000101",
			1621 => "0000001001000000000000001000001000",
			1622 => "0000000111000000001001001000000100",
			1623 => "11111110011110100001100111000101",
			1624 => "00000000000000000001100111000101",
			1625 => "00000000000000000001100111000101",
			1626 => "0000000111000000000110100100010100",
			1627 => "0000001101000000000101001000010000",
			1628 => "0000000010000000001100000000000100",
			1629 => "00000000000000000001100111000101",
			1630 => "0000001001000000000100101100000100",
			1631 => "00000000000000000001100111000101",
			1632 => "0000001110000000001011111000000100",
			1633 => "00000000111100100001100111000101",
			1634 => "00000000000000000001100111000101",
			1635 => "00000000000000000001100111000101",
			1636 => "0000000111000000001000011000001100",
			1637 => "0000001110000000001100010000000100",
			1638 => "00000000000000000001100111000101",
			1639 => "0000000101000000000111100000000100",
			1640 => "11111111001011010001100111000101",
			1641 => "00000000000000000001100111000101",
			1642 => "0000000101000000001110000100001100",
			1643 => "0000001111000000001100111000001000",
			1644 => "0000000010000000001010000100000100",
			1645 => "00000000000000000001100111000101",
			1646 => "00000000001010110001100111000101",
			1647 => "00000000000000000001100111000101",
			1648 => "00000000000000000001100111000101",
			1649 => "0000001001000000000101010000000100",
			1650 => "11111110011001110001101000011001",
			1651 => "0000001110000000001111010100011000",
			1652 => "0000001110000000000110010000000100",
			1653 => "00000001101001110001101000011001",
			1654 => "0000000100000000001111100100000100",
			1655 => "11111101110100000001101000011001",
			1656 => "0000001001000000000111101100000100",
			1657 => "11111110101101110001101000011001",
			1658 => "0000000110000000001111000000001000",
			1659 => "0000001000000000001010110000000100",
			1660 => "00000000011000010001101000011001",
			1661 => "00000001101101110001101000011001",
			1662 => "00000000011000100001101000011001",
			1663 => "0000001110000000001011111000001100",
			1664 => "0000001001000000001010100000000100",
			1665 => "11111110011011000001101000011001",
			1666 => "0000000100000000000010010100000100",
			1667 => "11111110100111110001101000011001",
			1668 => "00000001110011100001101000011001",
			1669 => "11111110011100110001101000011001",
			1670 => "0000000010000000001011111000100100",
			1671 => "0000001010000000000111110100100000",
			1672 => "0000001000000000001010110000010100",
			1673 => "0000001011000000000111010000000100",
			1674 => "00000000000000000001101010000101",
			1675 => "0000000111000000000001101000001100",
			1676 => "0000000011000000001110110100000100",
			1677 => "00000000000000000001101010000101",
			1678 => "0000001110000000000010000000000100",
			1679 => "00000000000000000001101010000101",
			1680 => "11111111011001110001101010000101",
			1681 => "00000000000000000001101010000101",
			1682 => "0000001110000000001111010100001000",
			1683 => "0000000001000000001011111100000100",
			1684 => "00000000000000000001101010000101",
			1685 => "00000000110000100001101010000101",
			1686 => "00000000000000000001101010000101",
			1687 => "11111111000100100001101010000101",
			1688 => "0000001101000000000111111100010000",
			1689 => "0000001000000000000001110000001100",
			1690 => "0000000100000000001011110000000100",
			1691 => "00000000000000000001101010000101",
			1692 => "0000001110000000001011111000000100",
			1693 => "00000001000001110001101010000101",
			1694 => "00000000000000000001101010000101",
			1695 => "00000000000000000001101010000101",
			1696 => "00000000000000000001101010000101",
			1697 => "0000001000000000000001110000110100",
			1698 => "0000001110000000001110110100010100",
			1699 => "0000000010000000000010000100001000",
			1700 => "0000000001000000001011111100000100",
			1701 => "11111111010010100001101011110001",
			1702 => "00000000000000000001101011110001",
			1703 => "0000000011000000001100000000001000",
			1704 => "0000000001000000000001000100000100",
			1705 => "00000000000000000001101011110001",
			1706 => "00000001010110000001101011110001",
			1707 => "00000000000000000001101011110001",
			1708 => "0000000001000000001101111100010000",
			1709 => "0000001011000000000111010000000100",
			1710 => "00000000000000000001101011110001",
			1711 => "0000000111000000000001101000001000",
			1712 => "0000000110000000001011001100000100",
			1713 => "00000000000000000001101011110001",
			1714 => "11111110101101010001101011110001",
			1715 => "00000000000000000001101011110001",
			1716 => "0000001000000000000101000100001100",
			1717 => "0000000100000000001101101100000100",
			1718 => "00000000000000000001101011110001",
			1719 => "0000001011000000000101100100000100",
			1720 => "00000001000111000001101011110001",
			1721 => "00000000000000000001101011110001",
			1722 => "11111111101011100001101011110001",
			1723 => "11111110100001000001101011110001",
			1724 => "0000000001000000001011111100001000",
			1725 => "0000001001000000001001111100000100",
			1726 => "11111110011111100001101101100101",
			1727 => "00000000000000000001101101100101",
			1728 => "0000001110000000000110111100010000",
			1729 => "0000000100000000001111100100001000",
			1730 => "0000001110000000000110010000000100",
			1731 => "00000000101110100001101101100101",
			1732 => "11111110110010010001101101100101",
			1733 => "0000001100000000001011000000000100",
			1734 => "00000001011011000001101101100101",
			1735 => "00000000000000000001101101100101",
			1736 => "0000001001000000000000001000001000",
			1737 => "0000000101000000000000110100000100",
			1738 => "00000000000000000001101101100101",
			1739 => "11111110011011010001101101100101",
			1740 => "0000001011000000000101100100001100",
			1741 => "0000001100000000000100011000001000",
			1742 => "0000000110000000001000010000000100",
			1743 => "00000001000001000001101101100101",
			1744 => "00000000000000000001101101100101",
			1745 => "00000000000000000001101101100101",
			1746 => "0000000001000000001101111100001100",
			1747 => "0000000111000000001000011000000100",
			1748 => "00000000000000000001101101100101",
			1749 => "0000001011000000000010001000000100",
			1750 => "00000000001111110001101101100101",
			1751 => "00000000000000000001101101100101",
			1752 => "11111111001000110001101101100101",
			1753 => "0000001001000000001001111100010100",
			1754 => "0000000000000000001010101100010000",
			1755 => "0000001001000000000101010000000100",
			1756 => "11111111000100100001101111101001",
			1757 => "0000001000000000001010110000001000",
			1758 => "0000000000000000001001101000000100",
			1759 => "00000000000000000001101111101001",
			1760 => "11111111111100110001101111101001",
			1761 => "00000000001111000001101111101001",
			1762 => "11111110011011110001101111101001",
			1763 => "0000000011000000001011111000100100",
			1764 => "0000000100000000000010010100011100",
			1765 => "0000001110000000000110111100010100",
			1766 => "0000001100000000001011000000001100",
			1767 => "0000001001000000001010100000001000",
			1768 => "0000000101000000001101000100000100",
			1769 => "00000001011000000001101111101001",
			1770 => "00000000000000000001101111101001",
			1771 => "00000000000000000001101111101001",
			1772 => "0000001000000000001010110000000100",
			1773 => "00000000000000000001101111101001",
			1774 => "11111111100110100001101111101001",
			1775 => "0000001111000000001000001100000100",
			1776 => "00000000000000000001101111101001",
			1777 => "11111110010110110001101111101001",
			1778 => "0000000110000000000100111100000100",
			1779 => "00000001100111010001101111101001",
			1780 => "00000000000000000001101111101001",
			1781 => "0000000101000000000110100000001000",
			1782 => "0000001001000000001010100100000100",
			1783 => "11111111001000100001101111101001",
			1784 => "00000000100100000001101111101001",
			1785 => "11111110101100110001101111101001",
			1786 => "0000000001000000000001000100000100",
			1787 => "11111110010111000001110001010101",
			1788 => "0000001101000000001111010000100000",
			1789 => "0000001110000000001011111000011100",
			1790 => "0000000001000000001101111100010100",
			1791 => "0000001101000000001110000100001100",
			1792 => "0000001000000000000110011000000100",
			1793 => "00000101100011000001110001010101",
			1794 => "0000001011000000000101100100000100",
			1795 => "00000011010001110001110001010101",
			1796 => "00000100110101000001110001010101",
			1797 => "0000000100000000001101101100000100",
			1798 => "11111111011100000001110001010101",
			1799 => "00000011010101000001110001010101",
			1800 => "0000001001000000001010100000000100",
			1801 => "00000101111010010001110001010101",
			1802 => "00000011001011110001110001010101",
			1803 => "11111110100000100001110001010101",
			1804 => "0000001110000000000111010100001000",
			1805 => "0000000001000000000001111000000100",
			1806 => "11111110010011000001110001010101",
			1807 => "00000011001000000001110001010101",
			1808 => "0000001110000000001011111000001000",
			1809 => "0000001111000000001011101100000100",
			1810 => "11111110011111000001110001010101",
			1811 => "00000001001000110001110001010101",
			1812 => "11111110010111010001110001010101",
			1813 => "0000000001000000001011111100000100",
			1814 => "11111110011001010001110010100001",
			1815 => "0000000011000000001111100100100000",
			1816 => "0000001110000000000110010000000100",
			1817 => "00000001101100110001110010100001",
			1818 => "0000000100000000001011101100001000",
			1819 => "0000000011000000001100010000000100",
			1820 => "11111111101001000001110010100001",
			1821 => "11111101101011100001110010100001",
			1822 => "0000001001000000000111101100000100",
			1823 => "11111111000001100001110010100001",
			1824 => "0000001110000000001000001100001000",
			1825 => "0000000111000000000001101000000100",
			1826 => "00000001100111110001110010100001",
			1827 => "00000000001101000001110010100001",
			1828 => "0000000100000000001110000000000100",
			1829 => "11111110011111110001110010100001",
			1830 => "00000001101001100001110010100001",
			1831 => "11111110011010100001110010100001",
			1832 => "0000001000000000000001110000111000",
			1833 => "0000000100000000001000000100101000",
			1834 => "0000001110000000001100010000011000",
			1835 => "0000000110000000001010011000001000",
			1836 => "0000000010000000000010000100000100",
			1837 => "11111111101011010001110100010101",
			1838 => "00000000000000000001110100010101",
			1839 => "0000001010000000000111110100001100",
			1840 => "0000001001000000001010100000001000",
			1841 => "0000001001000000001001111100000100",
			1842 => "00000000000000000001110100010101",
			1843 => "00000001000000110001110100010101",
			1844 => "00000000000000000001110100010101",
			1845 => "00000000000000000001110100010101",
			1846 => "0000001001000000000000001000001100",
			1847 => "0000000101000000001110101000001000",
			1848 => "0000001101000000001100100100000100",
			1849 => "00000000000000000001110100010101",
			1850 => "11111110101110100001110100010101",
			1851 => "00000000000000000001110100010101",
			1852 => "00000000000000000001110100010101",
			1853 => "0000000101000000000001000000001100",
			1854 => "0000001001000000000101010000000100",
			1855 => "00000000000000000001110100010101",
			1856 => "0000001110000000001111100100000100",
			1857 => "00000001010000010001110100010101",
			1858 => "00000000000000000001110100010101",
			1859 => "00000000000000000001110100010101",
			1860 => "11111110110001000001110100010101",
			1861 => "0000001001000000001001111100010100",
			1862 => "0000000000000000001010101100010000",
			1863 => "0000000001000000000001000100000100",
			1864 => "11111110111100010001110111000001",
			1865 => "0000000000000000001111001000001000",
			1866 => "0000000001000000001011111100000100",
			1867 => "11111111110010110001110111000001",
			1868 => "00000000000000000001110111000001",
			1869 => "00000000010101100001110111000001",
			1870 => "11111110011011000001110111000001",
			1871 => "0000000111000000000001101000100100",
			1872 => "0000000011000000001011111000011000",
			1873 => "0000001100000000001011000000010000",
			1874 => "0000000001000000001101111100001000",
			1875 => "0000001110000000001000001100000100",
			1876 => "00000001011101010001110111000001",
			1877 => "00000000000000000001110111000001",
			1878 => "0000000001000000000100110100000100",
			1879 => "11111111101001000001110111000001",
			1880 => "00000000100100110001110111000001",
			1881 => "0000001100000000001000000000000100",
			1882 => "11111111011101100001110111000001",
			1883 => "00000000000000000001110111000001",
			1884 => "0000000001000000000100110100000100",
			1885 => "11111110100111000001110111000001",
			1886 => "0000000101000000001110101000000100",
			1887 => "00000000101001010001110111000001",
			1888 => "00000000000000000001110111000001",
			1889 => "0000001010000000000111110100001100",
			1890 => "0000000011000000001000001100001000",
			1891 => "0000000000000000001001101000000100",
			1892 => "00000000000000000001110111000001",
			1893 => "00000000101110010001110111000001",
			1894 => "00000000000000000001110111000001",
			1895 => "0000000100000000000101000000000100",
			1896 => "11111110001100100001110111000001",
			1897 => "0000000000000000000111000000001000",
			1898 => "0000001001000000000010101100000100",
			1899 => "00000000001001100001110111000001",
			1900 => "00000000000000000001110111000001",
			1901 => "0000001100000000001010111000000100",
			1902 => "00000000000000000001110111000001",
			1903 => "11111111001001000001110111000001",
			1904 => "0000001000000000000001110000111000",
			1905 => "0000001110000000000110010000001100",
			1906 => "0000000110000000001010011000000100",
			1907 => "11111111010011110001111000110101",
			1908 => "0000000001000000000001000100000100",
			1909 => "00000000000000000001111000110101",
			1910 => "00000001010111100001111000110101",
			1911 => "0000001100000000000100011000011100",
			1912 => "0000000100000000001100111000001100",
			1913 => "0000001000000000001010110000001000",
			1914 => "0000000110000000001011001100000100",
			1915 => "00000000000000000001111000110101",
			1916 => "11111110111100110001111000110101",
			1917 => "00000000000000000001111000110101",
			1918 => "0000001110000000001010000100000100",
			1919 => "00000001001010010001111000110101",
			1920 => "0000000001000000001101111100000100",
			1921 => "11111110111011100001111000110101",
			1922 => "0000000100000000001011110000000100",
			1923 => "00000000000000000001111000110101",
			1924 => "00000000101001110001111000110101",
			1925 => "0000000111000000000110100100000100",
			1926 => "00000000000000000001111000110101",
			1927 => "0000000100000000000110001100001000",
			1928 => "0000000110000000001011001100000100",
			1929 => "00000000000000000001111000110101",
			1930 => "11111110100000010001111000110101",
			1931 => "00000000000000000001111000110101",
			1932 => "11111110100000010001111000110101",
			1933 => "0000000001000000000001000100000100",
			1934 => "11111110101010010001111011001001",
			1935 => "0000000111000000001001001000100000",
			1936 => "0000000100000000000010010100010100",
			1937 => "0000000011000000000111011000001000",
			1938 => "0000000001000000001101111100000100",
			1939 => "00000000101111010001111011001001",
			1940 => "00000000000000000001111011001001",
			1941 => "0000001100000000000100011000001000",
			1942 => "0000001101000000001100100100000100",
			1943 => "00000000000000000001111011001001",
			1944 => "11111111011011000001111011001001",
			1945 => "00000000000000000001111011001001",
			1946 => "0000001110000000001011111000001000",
			1947 => "0000001100000000000000001100000100",
			1948 => "00000000000000000001111011001001",
			1949 => "00000001011011000001111011001001",
			1950 => "00000000000000000001111011001001",
			1951 => "0000001100000000000100011000010000",
			1952 => "0000001000000000001100011100001000",
			1953 => "0000000011000000001100000000000100",
			1954 => "00000000000000000001111011001001",
			1955 => "11111111110011100001111011001001",
			1956 => "0000001000000000000001010100000100",
			1957 => "00000000110100100001111011001001",
			1958 => "00000000000000000001111011001001",
			1959 => "0000001110000000001100010000001100",
			1960 => "0000001101000000001110000100000100",
			1961 => "00000000010010010001111011001001",
			1962 => "0000001010000000000011101000000100",
			1963 => "11111111111000110001111011001001",
			1964 => "00000000000000000001111011001001",
			1965 => "0000000111000000000110100100000100",
			1966 => "00000000000000000001111011001001",
			1967 => "0000001000000000000110011100000100",
			1968 => "00000000000000000001111011001001",
			1969 => "11111110110010110001111011001001",
			1970 => "0000000001000000001011111100000100",
			1971 => "11111110011001000001111100011101",
			1972 => "0000000011000000001111100100100100",
			1973 => "0000001110000000000110010000000100",
			1974 => "00000001110000110001111100011101",
			1975 => "0000000100000000001011101100001100",
			1976 => "0000000011000000001100010000000100",
			1977 => "11111111100101000001111100011101",
			1978 => "0000000011000000000110111100000100",
			1979 => "11111101000010010001111100011101",
			1980 => "11111110100101100001111100011101",
			1981 => "0000001001000000000111101100000100",
			1982 => "11111110110100100001111100011101",
			1983 => "0000001110000000001000001100001000",
			1984 => "0000000111000000000001101000000100",
			1985 => "00000001110000000001111100011101",
			1986 => "00000000011101000001111100011101",
			1987 => "0000000100000000001110000000000100",
			1988 => "11111110011110100001111100011101",
			1989 => "00000001111100110001111100011101",
			1990 => "11111110011001110001111100011101",
			1991 => "0000000001000000000001000100000100",
			1992 => "11111110011000000001111110000001",
			1993 => "0000001101000000001001010000100100",
			1994 => "0000001000000000000001110000100000",
			1995 => "0000000010000000001101101100011100",
			1996 => "0000001101000000000101001000010000",
			1997 => "0000001100000000000100011000001000",
			1998 => "0000000100000000001101101100000100",
			1999 => "00000010001001100001111110000001",
			2000 => "00000010011011000001111110000001",
			2001 => "0000000010000000000111010100000100",
			2002 => "00000000011000000001111110000001",
			2003 => "00000001111100100001111110000001",
			2004 => "0000000000000000001111001000000100",
			2005 => "11111110011101000001111110000001",
			2006 => "0000000110000000001111000000000100",
			2007 => "00000010011011010001111110000001",
			2008 => "11111110110000110001111110000001",
			2009 => "00000100011100010001111110000001",
			2010 => "11111110010001100001111110000001",
			2011 => "0000000011000000001011111000001000",
			2012 => "0000000001000000000001111000000100",
			2013 => "11111110011000010001111110000001",
			2014 => "00000001000011100001111110000001",
			2015 => "11111110011000010001111110000001",
			2016 => "0000000001000000000001000100000100",
			2017 => "11111110011001100001111111100101",
			2018 => "0000001110000000001011111000101100",
			2019 => "0000000011000000001100010000001000",
			2020 => "0000000001000000001011111100000100",
			2021 => "00000010110001110001111111100101",
			2022 => "00000001101011110001111111100101",
			2023 => "0000000100000000001011101100001100",
			2024 => "0000001110000000001110110100000100",
			2025 => "11111111010111000001111111100101",
			2026 => "0000000111000000000110100100000100",
			2027 => "11111100110110100001111111100101",
			2028 => "11111110010010100001111111100101",
			2029 => "0000001001000000000111101100001000",
			2030 => "0000000110000000001011001100000100",
			2031 => "00000000110110100001111111100101",
			2032 => "11111110010101010001111111100101",
			2033 => "0000000100000000000011000000001000",
			2034 => "0000001010000000000111110100000100",
			2035 => "00000001010011110001111111100101",
			2036 => "11111100011011000001111111100101",
			2037 => "0000000010000000001101101100000100",
			2038 => "00000001100111110001111111100101",
			2039 => "00000010111010010001111111100101",
			2040 => "11111110011011000001111111100101",
			2041 => "0000000001000000000001000100000100",
			2042 => "11111110011001000010000000111001",
			2043 => "0000001110000000001011111000100100",
			2044 => "0000001000000000000001110000100000",
			2045 => "0000001110000000000110010000000100",
			2046 => "00000001110101000010000000111001",
			2047 => "0000000010000000001111010100001100",
			2048 => "0000000011000000001100010000000100",
			2049 => "11111111110100100010000000111001",
			2050 => "0000001010000000000010101100000100",
			2051 => "11111110100101100010000000111001",
			2052 => "11111101000101010010000000111001",
			2053 => "0000001001000000000111101100001000",
			2054 => "0000001100000000000100011000000100",
			2055 => "00000000111000100010000000111001",
			2056 => "11111101101000010010000000111001",
			2057 => "0000001001000000000111101100000100",
			2058 => "00001000011001110010000000111001",
			2059 => "00000001101100000010000000111001",
			2060 => "11111110000010110010000000111001",
			2061 => "11111110011001110010000000111001",
			2062 => "0000001000000000000001110000111000",
			2063 => "0000000110000000001010011000000100",
			2064 => "11111110101011010010000010101101",
			2065 => "0000001101000000000111100000010100",
			2066 => "0000000111000000001110110000001100",
			2067 => "0000000001000000001011111100001000",
			2068 => "0000000010000000000110111100000100",
			2069 => "11111111110000100010000010101101",
			2070 => "00000000000000000010000010101101",
			2071 => "00000000101100110010000010101101",
			2072 => "0000000110000000001111000000000100",
			2073 => "00000001011101010010000010101101",
			2074 => "00000000000000000010000010101101",
			2075 => "0000000100000000001000000100010100",
			2076 => "0000001110000000000111010100010000",
			2077 => "0000000010000000000111010100001000",
			2078 => "0000001110000000000010000100000100",
			2079 => "00000000100101010010000010101101",
			2080 => "11111110110001010010000010101101",
			2081 => "0000001101000000001111010000000100",
			2082 => "00000001010000110010000010101101",
			2083 => "11111111101001110010000010101101",
			2084 => "11111110100010000010000010101101",
			2085 => "0000000101000000000001000000001000",
			2086 => "0000001110000000001111100100000100",
			2087 => "00000001101100110010000010101101",
			2088 => "00000000000000000010000010101101",
			2089 => "11111111000111100010000010101101",
			2090 => "11111110011100000010000010101101",
			2091 => "0000001000000000000001110000110100",
			2092 => "0000000110000000001010011000000100",
			2093 => "11111110110000000010000100011001",
			2094 => "0000001101000000000111100000010100",
			2095 => "0000000001000000000001000100000100",
			2096 => "00000000000000000010000100011001",
			2097 => "0000000110000000001111000000001100",
			2098 => "0000001100000000000100001000001000",
			2099 => "0000001100000000000100001000000100",
			2100 => "00000000100010000010000100011001",
			2101 => "00000000000000000010000100011001",
			2102 => "00000001011010000010000100011001",
			2103 => "00000000000000000010000100011001",
			2104 => "0000001100000000001010111000000100",
			2105 => "11111110101111110010000100011001",
			2106 => "0000001001000000000111101100001100",
			2107 => "0000001100000000000100011000000100",
			2108 => "00000000000000000010000100011001",
			2109 => "0000000010000000001111010100000100",
			2110 => "00000000000000000010000100011001",
			2111 => "11111110111010100010000100011001",
			2112 => "0000001101000000000111111100001000",
			2113 => "0000000100000000001110000000000100",
			2114 => "00000000000011100010000100011001",
			2115 => "00000001100101000010000100011001",
			2116 => "11111111001011000010000100011001",
			2117 => "11111110011101000010000100011001",
			2118 => "0000000001000000000001000100000100",
			2119 => "11111110011010000010000110010101",
			2120 => "0000001110000000000110010000000100",
			2121 => "00000001101100000010000110010101",
			2122 => "0000001100000000000100011000011100",
			2123 => "0000000100000000000110101100000100",
			2124 => "11111101111110100010000110010101",
			2125 => "0000001110000000001100000000001000",
			2126 => "0000000010000000000110111100000100",
			2127 => "00000000000000000010000110010101",
			2128 => "00000001100111000010000110010101",
			2129 => "0000000100000000000010010100001000",
			2130 => "0000001100000000000100011000000100",
			2131 => "11111110011010000010000110010101",
			2132 => "00000000000011010010000110010101",
			2133 => "0000001110000000001011111000000100",
			2134 => "00000001011101010010000110010101",
			2135 => "11111110110110110010000110010101",
			2136 => "0000000111000000000110100100001000",
			2137 => "0000000011000000000000010000000100",
			2138 => "00000001000001000010000110010101",
			2139 => "00000000000000000010000110010101",
			2140 => "0000001100000000000100011000001000",
			2141 => "0000000001000000001101111100000100",
			2142 => "11111011110000110010000110010101",
			2143 => "00000000000000000010000110010101",
			2144 => "0000001110000000000111010100001000",
			2145 => "0000001001000000000111101100000100",
			2146 => "11111110011000110010000110010101",
			2147 => "00000001001010110010000110010101",
			2148 => "11111110011110100010000110010101",
			2149 => "0000000001000000000001000100000100",
			2150 => "11111110011011100010001000111011",
			2151 => "0000001110000000000110010000001000",
			2152 => "0000000110000000001010011000000100",
			2153 => "00000000000000000010001000111011",
			2154 => "00000001100100000010001000111011",
			2155 => "0000001100000000001010111000010100",
			2156 => "0000001101000000001100100100001100",
			2157 => "0000000001000000000111101000000100",
			2158 => "11111111001011010010001000111011",
			2159 => "0000000100000000001110100100000100",
			2160 => "00000001000000100010001000111011",
			2161 => "00000000000000000010001000111011",
			2162 => "0000000001000000001101111100000100",
			2163 => "11111110010100110010001000111011",
			2164 => "00000000000000000010001000111011",
			2165 => "0000000111000000000001101000011100",
			2166 => "0000001010000000000011101000001100",
			2167 => "0000000010000000001100000000000100",
			2168 => "11111111000001000010001000111011",
			2169 => "0000001101000000001110000100000100",
			2170 => "00000001000011010010001000111011",
			2171 => "11111111100100110010001000111011",
			2172 => "0000000110000000000100111100001000",
			2173 => "0000000100000000001100111000000100",
			2174 => "00000000000000000010001000111011",
			2175 => "00000001101101110010001000111011",
			2176 => "0000001101000000000101001000000100",
			2177 => "00000000000000000010001000111011",
			2178 => "11111111001010000010001000111011",
			2179 => "0000001100000000000100011000001100",
			2180 => "0000001010000000000011101000000100",
			2181 => "00000000000000000010001000111011",
			2182 => "0000000110000000001000010000000100",
			2183 => "00000001000110110010001000111011",
			2184 => "00000000000000000010001000111011",
			2185 => "0000001000000000001100011100000100",
			2186 => "00000000000000000010001000111011",
			2187 => "0000000100000000000101000000000100",
			2188 => "11111101111000110010001000111011",
			2189 => "11111111010011100010001000111011",
			2190 => "00000000000000000010001000111101",
			2191 => "00000000000000000010001001000001",
			2192 => "00000000000000000010001001000101",
			2193 => "00000000000000000010001001001001",
			2194 => "00000000000000000010001001001101",
			2195 => "00000000000000000010001001010001",
			2196 => "00000000000000000010001001010101",
			2197 => "00000000000000000010001001011001",
			2198 => "00000000000000000010001001011101",
			2199 => "00000000000000000010001001100001",
			2200 => "00000000000000000010001001100101",
			2201 => "00000000000000000010001001101001",
			2202 => "00000000000000000010001001101101",
			2203 => "00000000000000000010001001110001",
			2204 => "00000000000000000010001001110101",
			2205 => "00000000000000000010001001111001",
			2206 => "00000000000000000010001001111101",
			2207 => "00000000000000000010001010000001",
			2208 => "00000000000000000010001010000101",
			2209 => "00000000000000000010001010001001",
			2210 => "00000000000000000010001010001101",
			2211 => "00000000000000000010001010010001",
			2212 => "00000000000000000010001010010101",
			2213 => "00000000000000000010001010011001",
			2214 => "00000000000000000010001010011101",
			2215 => "00000000000000000010001010100001",
			2216 => "00000000000000000010001010100101",
			2217 => "0000001110000000001100000000000100",
			2218 => "00000000000000000010001010110001",
			2219 => "11111111111111000010001010110001",
			2220 => "0000001000000000001100011100000100",
			2221 => "00000000000000000010001010111101",
			2222 => "11111111111101010010001010111101",
			2223 => "0000001001000000000000001000000100",
			2224 => "11111111111111010010001011001001",
			2225 => "00000000000000000010001011001001",
			2226 => "0000001110000000000110010000001000",
			2227 => "0000001110000000000101001000000100",
			2228 => "00000000000000000010001011011101",
			2229 => "00000000001010000010001011011101",
			2230 => "11111111111110110010001011011101",
			2231 => "0000000001000000000111101000001000",
			2232 => "0000001001000000000111101100000100",
			2233 => "11111111111001000010001011110001",
			2234 => "00000000000000000010001011110001",
			2235 => "00000000000000000010001011110001",
			2236 => "0000000001000000001011111100000100",
			2237 => "00000000000000000010001100000101",
			2238 => "0000001001000000001010100100000100",
			2239 => "00000000000110010010001100000101",
			2240 => "00000000000000000010001100000101",
			2241 => "0000001110000000000110010000001100",
			2242 => "0000001110000000000101001000000100",
			2243 => "00000000000000000010001100100001",
			2244 => "0000000011000000001100000000000100",
			2245 => "00000000001100110010001100100001",
			2246 => "00000000000000000010001100100001",
			2247 => "11111111111100110010001100100001",
			2248 => "0000000001000000001101111100001100",
			2249 => "0000001100000000001011000000001000",
			2250 => "0000001000000000001010110000000100",
			2251 => "00000000000000000010001100111101",
			2252 => "11111111110011000010001100111101",
			2253 => "00000000000000000010001100111101",
			2254 => "00000000000000000010001100111101",
			2255 => "0000001110000000001100000000001100",
			2256 => "0000001111000000001100010000000100",
			2257 => "00000000000000000010001101100001",
			2258 => "0000001111000000001000001100000100",
			2259 => "00000000000001010010001101100001",
			2260 => "00000000000000000010001101100001",
			2261 => "0000001111000000001000001100000100",
			2262 => "00000000000000000010001101100001",
			2263 => "11111111111110110010001101100001",
			2264 => "0000001110000000000110010000001100",
			2265 => "0000001001000000000101010000000100",
			2266 => "00000000000000000010001110001101",
			2267 => "0000000000000000001100000100000100",
			2268 => "00000000000000000010001110001101",
			2269 => "00000000001100010010001110001101",
			2270 => "0000000001000000000100110100001000",
			2271 => "0000001100000000000100001000000100",
			2272 => "00000000000000000010001110001101",
			2273 => "11111111101110110010001110001101",
			2274 => "00000000000000000010001110001101",
			2275 => "0000000001000000001110010100000100",
			2276 => "00000000000000000010001110110001",
			2277 => "0000001001000000001010100100001100",
			2278 => "0000001000000000000001110000001000",
			2279 => "0000001000000000001010110000000100",
			2280 => "00000000000000000010001110110001",
			2281 => "00000000001010100010001110110001",
			2282 => "00000000000000000010001110110001",
			2283 => "00000000000000000010001110110001",
			2284 => "0000001000000000000001010100010000",
			2285 => "0000001101000000001111010000001100",
			2286 => "0000001000000000001000010100000100",
			2287 => "00000000000000000010001111010101",
			2288 => "0000001101000000000101110100000100",
			2289 => "00000000000000000010001111010101",
			2290 => "00000000001100010010001111010101",
			2291 => "00000000000000000010001111010101",
			2292 => "00000000000000000010001111010101",
			2293 => "0000001001000000000000001000010000",
			2294 => "0000001110000000000110010000000100",
			2295 => "00000000000000000010001111111001",
			2296 => "0000000010000000000011000000001000",
			2297 => "0000000011000000001100010000000100",
			2298 => "00000000000000000010001111111001",
			2299 => "11111111110111010010001111111001",
			2300 => "00000000000000000010001111111001",
			2301 => "00000000000000000010001111111001",
			2302 => "0000001110000000000110010000010000",
			2303 => "0000001110000000000101001000000100",
			2304 => "00000000000000000010010000100101",
			2305 => "0000000010000000001110010000000100",
			2306 => "00000000000000000010010000100101",
			2307 => "0000000010000000001100111000000100",
			2308 => "00000000001100010010010000100101",
			2309 => "00000000000000000010010000100101",
			2310 => "0000000100000000000011000000000100",
			2311 => "11111111110001010010010000100101",
			2312 => "00000000000000000010010000100101",
			2313 => "0000001001000000000111101100001000",
			2314 => "0000001011000000000100000100000100",
			2315 => "00000000000000000010010001011001",
			2316 => "11111111100101100010010001011001",
			2317 => "0000000100000000001101101100000100",
			2318 => "00000000000000000010010001011001",
			2319 => "0000001111000000001100111000001100",
			2320 => "0000001100000000001000000000001000",
			2321 => "0000001010000000001000010100000100",
			2322 => "00000000011110110010010001011001",
			2323 => "00000000000000000010010001011001",
			2324 => "00000000000000000010010001011001",
			2325 => "00000000000000000010010001011001",
			2326 => "0000001110000000000110010000000100",
			2327 => "00000000000000000010010010000101",
			2328 => "0000001001000000000000001000010000",
			2329 => "0000001100000000001011000000001100",
			2330 => "0000001100000000000100001000000100",
			2331 => "00000000000000000010010010000101",
			2332 => "0000000001000000001101111100000100",
			2333 => "11111111110000000010010010000101",
			2334 => "00000000000000000010010010000101",
			2335 => "00000000000000000010010010000101",
			2336 => "00000000000000000010010010000101",
			2337 => "0000000010000000001000001100010100",
			2338 => "0000001110000000000110010000001000",
			2339 => "0000000001000000001011111100000100",
			2340 => "11111111101101110010010011010001",
			2341 => "00000000011001010010010011010001",
			2342 => "0000000100000000001101101100001000",
			2343 => "0000001100000000001000000000000100",
			2344 => "11111111001011010010010011010001",
			2345 => "00000000000000000010010011010001",
			2346 => "00000000000000000010010011010001",
			2347 => "0000001110000000000111010100001100",
			2348 => "0000000000000000001111000100001000",
			2349 => "0000000001000000000001000100000100",
			2350 => "00000000000000000010010011010001",
			2351 => "00000000101111100010010011010001",
			2352 => "00000000000000000010010011010001",
			2353 => "0000000001000000001101111100000100",
			2354 => "11111111110000110010010011010001",
			2355 => "00000000000000000010010011010001",
			2356 => "0000000010000000001010000100010000",
			2357 => "0000001100000000001000000000001100",
			2358 => "0000000110000000001001100100001000",
			2359 => "0000001110000000000010000000000100",
			2360 => "00000000000000000010010100011101",
			2361 => "11111111101101110010010100011101",
			2362 => "00000000000000000010010100011101",
			2363 => "00000000000000000010010100011101",
			2364 => "0000001110000000001100000000010000",
			2365 => "0000000110000000001101011000000100",
			2366 => "00000000000000000010010100011101",
			2367 => "0000001100000000001011000000001000",
			2368 => "0000001010000000001000010100000100",
			2369 => "00000000011111100010010100011101",
			2370 => "00000000000000000010010100011101",
			2371 => "00000000000000000010010100011101",
			2372 => "0000000100000000000010010100000100",
			2373 => "11111111110010000010010100011101",
			2374 => "00000000000000000010010100011101",
			2375 => "0000000001000000001110010100001100",
			2376 => "0000001001000000000100101100001000",
			2377 => "0000000100000000001100010000000100",
			2378 => "00000000000000000010010101100001",
			2379 => "11111111110111000010010101100001",
			2380 => "00000000000000000010010101100001",
			2381 => "0000001101000000000111111100010100",
			2382 => "0000000100000000000001011100000100",
			2383 => "00000000000000000010010101100001",
			2384 => "0000001110000000001011111000001100",
			2385 => "0000000110000000000100111100001000",
			2386 => "0000000000000000000110001000000100",
			2387 => "00000000000000000010010101100001",
			2388 => "00000000100110100010010101100001",
			2389 => "00000000000000000010010101100001",
			2390 => "00000000000000000010010101100001",
			2391 => "00000000000000000010010101100001",
			2392 => "0000001100000000001010111100001100",
			2393 => "0000001000000000001010110000000100",
			2394 => "00000000000000000010010110101101",
			2395 => "0000000001000000000111101000000100",
			2396 => "11111111110110010010010110101101",
			2397 => "00000000000000000010010110101101",
			2398 => "0000000100000000000011000000001000",
			2399 => "0000001000000000001100011100000100",
			2400 => "00000000000000000010010110101101",
			2401 => "11111111110100110010010110101101",
			2402 => "0000000110000000000100111100010000",
			2403 => "0000001000000000000001110000001100",
			2404 => "0000000010000000001111101000001000",
			2405 => "0000001100000000001001110100000100",
			2406 => "00000000101110110010010110101101",
			2407 => "00000000000000000010010110101101",
			2408 => "00000000000000000010010110101101",
			2409 => "00000000000000000010010110101101",
			2410 => "00000000000000000010010110101101",
			2411 => "0000001100000000001010111000000100",
			2412 => "00000000000000000010010111100001",
			2413 => "0000001101000000000010011100010100",
			2414 => "0000001100000000001011000000010000",
			2415 => "0000001110000000001011111000001100",
			2416 => "0000000001000000001011111100000100",
			2417 => "00000000000000000010010111100001",
			2418 => "0000001101000000001001010000000100",
			2419 => "00000000100001110010010111100001",
			2420 => "00000000000000000010010111100001",
			2421 => "00000000000000000010010111100001",
			2422 => "00000000000000000010010111100001",
			2423 => "00000000000000000010010111100001",
			2424 => "0000000001000000000111101000010000",
			2425 => "0000001100000000001010111100001100",
			2426 => "0000000111000000001000000000001000",
			2427 => "0000000100000000000110101100000100",
			2428 => "00000000000000000010011000110101",
			2429 => "11111111101101010010011000110101",
			2430 => "00000000000000000010011000110101",
			2431 => "00000000000000000010011000110101",
			2432 => "0000000100000000000001011100001000",
			2433 => "0000000001000000000001111000000100",
			2434 => "00000000000000000010011000110101",
			2435 => "11111111111110110010011000110101",
			2436 => "0000001111000000000011000000010000",
			2437 => "0000000110000000000100111100001100",
			2438 => "0000000001000000001100011000001000",
			2439 => "0000001100000000001000000000000100",
			2440 => "00000000100111010010011000110101",
			2441 => "00000000000000000010011000110101",
			2442 => "00000000000000000010011000110101",
			2443 => "00000000000000000010011000110101",
			2444 => "00000000000000000010011000110101",
			2445 => "0000000001000000001011111100001000",
			2446 => "0000000001000000000001000100000100",
			2447 => "11001000111111000010011010010001",
			2448 => "11001011111110000010011010010001",
			2449 => "0000000011000000001111010100010100",
			2450 => "0000001011000000000101100100001100",
			2451 => "0000001000000000000110011000000100",
			2452 => "11100100101000000010011010010001",
			2453 => "0000000001000000001101111100000100",
			2454 => "11110110111001000010011010010001",
			2455 => "11100110001101010010011010010001",
			2456 => "0000000000000000001011010100000100",
			2457 => "11001001010001100010011010010001",
			2458 => "11100111111110010010011010010001",
			2459 => "0000001110000000000111010100001000",
			2460 => "0000000100000000000011000000000100",
			2461 => "11001001000010010010011010010001",
			2462 => "11110100000011000010011010010001",
			2463 => "0000001110000000001011111000001000",
			2464 => "0000000001000000001101111100000100",
			2465 => "11001001000100000010011010010001",
			2466 => "11010100111001010010011010010001",
			2467 => "11001000111111000010011010010001",
			2468 => "0000000010000000001011111000100000",
			2469 => "0000001010000000000111110100011000",
			2470 => "0000001110000000001100010000010000",
			2471 => "0000001001000000001010100000001100",
			2472 => "0000000001000000001110010100000100",
			2473 => "00000000000000000010011011110101",
			2474 => "0000000101000000000110100000000100",
			2475 => "00000000101110010010011011110101",
			2476 => "00000000000000000010011011110101",
			2477 => "00000000000000000010011011110101",
			2478 => "0000000001000000001101111100000100",
			2479 => "11111111110111100010011011110101",
			2480 => "00000000000000000010011011110101",
			2481 => "0000000010000000000000010000000100",
			2482 => "11111110110000110010011011110101",
			2483 => "00000000000000000010011011110101",
			2484 => "0000000011000000001011111000001100",
			2485 => "0000000110000000000100111100001000",
			2486 => "0000000001000000000001000100000100",
			2487 => "00000000000000000010011011110101",
			2488 => "00000001000100110010011011110101",
			2489 => "00000000000000000010011011110101",
			2490 => "0000000001000000001101111100000100",
			2491 => "11111111100110000010011011110101",
			2492 => "00000000000000000010011011110101",
			2493 => "0000001100000000001010111000001100",
			2494 => "0000001000000000001100011100000100",
			2495 => "00000000000000000010011101011001",
			2496 => "0000001001000000000000001000000100",
			2497 => "11111110110011000010011101011001",
			2498 => "00000000000000000010011101011001",
			2499 => "0000000111000000001001001000010000",
			2500 => "0000000100000000000110101100000100",
			2501 => "00000000000000000010011101011001",
			2502 => "0000001110000000001111100100001000",
			2503 => "0000000001000000001011111100000100",
			2504 => "00000000000000000010011101011001",
			2505 => "00000000111001000010011101011001",
			2506 => "00000000000000000010011101011001",
			2507 => "0000001100000000000100011000001100",
			2508 => "0000001101000000000101001000001000",
			2509 => "0000000001000000001110010100000100",
			2510 => "00000000000000000010011101011001",
			2511 => "00000000011001010010011101011001",
			2512 => "00000000000000000010011101011001",
			2513 => "0000001000000000000110011100000100",
			2514 => "00000000000000000010011101011001",
			2515 => "0000000100000000000101000000000100",
			2516 => "11111111000111100010011101011001",
			2517 => "00000000000000000010011101011001",
			2518 => "0000001100000000001010111100001100",
			2519 => "0000000001000000000111101000001000",
			2520 => "0000000000000000001001101000000100",
			2521 => "00000000000000000010011110111101",
			2522 => "11111111100000100010011110111101",
			2523 => "00000000000000000010011110111101",
			2524 => "0000000111000000001001001000001100",
			2525 => "0000000110000000000100111100001000",
			2526 => "0000000001000000000001000100000100",
			2527 => "00000000000000000010011110111101",
			2528 => "00000000101101010010011110111101",
			2529 => "00000000000000000010011110111101",
			2530 => "0000001001000000000000001000010000",
			2531 => "0000001110000000001110110100000100",
			2532 => "00000000000000000010011110111101",
			2533 => "0000000110000000001011001100000100",
			2534 => "00000000000000000010011110111101",
			2535 => "0000000001000000001101111100000100",
			2536 => "11111111010000110010011110111101",
			2537 => "00000000000000000010011110111101",
			2538 => "0000001100000000000100011000001000",
			2539 => "0000001110000000001011111000000100",
			2540 => "00000000011110000010011110111101",
			2541 => "00000000000000000010011110111101",
			2542 => "00000000000000000010011110111101",
			2543 => "0000000001000000000111101000100000",
			2544 => "0000001000000000000110011100011000",
			2545 => "0000001000000000001001000100001000",
			2546 => "0000001010000000001010100100000100",
			2547 => "11111111100000000010100000110001",
			2548 => "00000000000000000010100000110001",
			2549 => "0000001110000000001100000000001100",
			2550 => "0000001001000000000101010000000100",
			2551 => "00000000000000000010100000110001",
			2552 => "0000000101000000001101000100000100",
			2553 => "00000000100011100010100000110001",
			2554 => "00000000000000000010100000110001",
			2555 => "00000000000000000010100000110001",
			2556 => "0000000001000000000111101000000100",
			2557 => "11111110111100010010100000110001",
			2558 => "00000000000000000010100000110001",
			2559 => "0000001110000000001000001100010100",
			2560 => "0000001010000000000011101000001100",
			2561 => "0000000011000000000111011000001000",
			2562 => "0000000001000000001101111100000100",
			2563 => "00000000011101100010100000110001",
			2564 => "00000000000000000010100000110001",
			2565 => "11111111100010110010100000110001",
			2566 => "0000000011000000000000010000000100",
			2567 => "00000001001010100010100000110001",
			2568 => "00000000000000000010100000110001",
			2569 => "0000000101000000000110100000000100",
			2570 => "00000000000000000010100000110001",
			2571 => "11111111100111110010100000110001",
			2572 => "0000001100000000001010111100010000",
			2573 => "0000000001000000000111101000001100",
			2574 => "0000001000000000000001010000000100",
			2575 => "00000000000000000010100010011101",
			2576 => "0000000111000000001000000000000100",
			2577 => "11111111011111110010100010011101",
			2578 => "00000000000000000010100010011101",
			2579 => "00000000000000000010100010011101",
			2580 => "0000000111000000001001001000001100",
			2581 => "0000001001000000001010100000001000",
			2582 => "0000000001000000000001000100000100",
			2583 => "00000000000000000010100010011101",
			2584 => "00000000101101110010100010011101",
			2585 => "00000000000000000010100010011101",
			2586 => "0000001111000000001000001100010000",
			2587 => "0000001010000000000010101100000100",
			2588 => "00000000000000000010100010011101",
			2589 => "0000001000000000000110011100001000",
			2590 => "0000000010000000001100000000000100",
			2591 => "00000000000000000010100010011101",
			2592 => "00000000011111110010100010011101",
			2593 => "00000000000000000010100010011101",
			2594 => "0000000001000000001101111100001000",
			2595 => "0000001110000000001100010000000100",
			2596 => "00000000000000000010100010011101",
			2597 => "11111111011111000010100010011101",
			2598 => "00000000000000000010100010011101",
			2599 => "0000001100000000001010111000011100",
			2600 => "0000000010000000001000001100010000",
			2601 => "0000001011000000000101100100001100",
			2602 => "0000001101000000000101001000001000",
			2603 => "0000000111000000001001001000000100",
			2604 => "11111110110111110010100100011001",
			2605 => "00000000000000000010100100011001",
			2606 => "00000000000000000010100100011001",
			2607 => "00000000000000000010100100011001",
			2608 => "0000001110000000001010000100001000",
			2609 => "0000001101000000001011110100000100",
			2610 => "00000000000000000010100100011001",
			2611 => "00000000000100010010100100011001",
			2612 => "00000000000000000010100100011001",
			2613 => "0000001101000000000101001000010100",
			2614 => "0000001100000000000100011000010000",
			2615 => "0000000010000000001100000000000100",
			2616 => "00000000000000000010100100011001",
			2617 => "0000001110000000001011111000001000",
			2618 => "0000000110000000001101011000000100",
			2619 => "00000000000000000010100100011001",
			2620 => "00000000110101100010100100011001",
			2621 => "00000000000000000010100100011001",
			2622 => "00000000000000000010100100011001",
			2623 => "0000000100000000001011110000001100",
			2624 => "0000001100000000001010111000000100",
			2625 => "00000000000000000010100100011001",
			2626 => "0000001011000000000100000100000100",
			2627 => "00000000000000000010100100011001",
			2628 => "11111111011100100010100100011001",
			2629 => "00000000000000000010100100011001",
			2630 => "0000001001000000001001111100000100",
			2631 => "00000000000000000010100101010101",
			2632 => "0000000101000000000001000000011000",
			2633 => "0000000000000000001001101000000100",
			2634 => "00000000000000000010100101010101",
			2635 => "0000000110000000000100111100010000",
			2636 => "0000001110000000001011111000001100",
			2637 => "0000000111000000000011100000000100",
			2638 => "00000000000000000010100101010101",
			2639 => "0000001010000000000011101000000100",
			2640 => "00000000000000000010100101010101",
			2641 => "00000000011001100010100101010101",
			2642 => "00000000000000000010100101010101",
			2643 => "00000000000000000010100101010101",
			2644 => "00000000000000000010100101010101",
			2645 => "0000000010000000001100000000000100",
			2646 => "00000000000000000010100110010001",
			2647 => "0000001011000000000101100100011000",
			2648 => "0000001000000000001010110000000100",
			2649 => "00000000000000000010100110010001",
			2650 => "0000000111000000000001101000010000",
			2651 => "0000000100000000001011101100000100",
			2652 => "00000000000000000010100110010001",
			2653 => "0000001000000000000001110000001000",
			2654 => "0000001110000000001011111000000100",
			2655 => "00000000100110110010100110010001",
			2656 => "00000000000000000010100110010001",
			2657 => "00000000000000000010100110010001",
			2658 => "00000000000000000010100110010001",
			2659 => "00000000000000000010100110010001",
			2660 => "0000001001000000000101010000001100",
			2661 => "0000001001000000000101010000000100",
			2662 => "11111110010110100010100111111101",
			2663 => "0000001001000000000101010000000100",
			2664 => "11111111111101100010100111111101",
			2665 => "11111110100011100010100111111101",
			2666 => "0000001101000000001111010000011000",
			2667 => "0000001110000000001011111000010100",
			2668 => "0000001111000000001001100000000100",
			2669 => "00000101110111110010100111111101",
			2670 => "0000000000000000001001101000000100",
			2671 => "00000001011001100010100111111101",
			2672 => "0000001111000000001011101100001000",
			2673 => "0000001001000000001010100000000100",
			2674 => "00000100000101010010100111111101",
			2675 => "00000010010000110010100111111101",
			2676 => "00000110101010110010100111111101",
			2677 => "11111110011110110010100111111101",
			2678 => "0000001110000000000111010100001000",
			2679 => "0000001001000000000000001000000100",
			2680 => "11111110010001110010100111111101",
			2681 => "00000011100101100010100111111101",
			2682 => "0000001110000000001011111000001000",
			2683 => "0000001100000000000100011000000100",
			2684 => "00000001010111010010100111111101",
			2685 => "11111110011110010010100111111101",
			2686 => "11111110010110110010100111111101",
			2687 => "0000001001000000000101010000000100",
			2688 => "11111110011001110010101001010001",
			2689 => "0000001110000000001111010100010100",
			2690 => "0000001110000000000110010000000100",
			2691 => "00000001101010100010101001010001",
			2692 => "0000000100000000001111100100000100",
			2693 => "11111101101010100010101001010001",
			2694 => "0000001001000000000111101100000100",
			2695 => "11111110101000010010101001010001",
			2696 => "0000000110000000001111000000000100",
			2697 => "00000001101011110010101001010001",
			2698 => "00000000011111000010101001010001",
			2699 => "0000001100000000000100011000010000",
			2700 => "0000000100000000000010010100000100",
			2701 => "11111110010101100010101001010001",
			2702 => "0000001110000000001011111000001000",
			2703 => "0000000010000000001100111000000100",
			2704 => "00000000100010010010101001010001",
			2705 => "00000010000011000010101001010001",
			2706 => "11111110101111000010101001010001",
			2707 => "11111110011100010010101001010001",
			2708 => "0000001100000000001010111000100000",
			2709 => "0000000010000000001000001100010000",
			2710 => "0000001011000000000101100100001100",
			2711 => "0000001101000000000101001000001000",
			2712 => "0000000111000000001001001000000100",
			2713 => "11111110101101000010101011100101",
			2714 => "00000000000000000010101011100101",
			2715 => "00000000000000000010101011100101",
			2716 => "00000000000000000010101011100101",
			2717 => "0000001110000000001010000100001100",
			2718 => "0000001011000000001001001000000100",
			2719 => "00000000000000000010101011100101",
			2720 => "0000000010000000001100111000000100",
			2721 => "00000000001001100010101011100101",
			2722 => "00000000000000000010101011100101",
			2723 => "00000000000000000010101011100101",
			2724 => "0000001001000000000111101100001100",
			2725 => "0000001100000000000100011000000100",
			2726 => "00000000000000000010101011100101",
			2727 => "0000001100000000001000000000000100",
			2728 => "11111111010101000010101011100101",
			2729 => "00000000000000000010101011100101",
			2730 => "0000001101000000000101001000001100",
			2731 => "0000000010000000001100000000000100",
			2732 => "00000000000000000010101011100101",
			2733 => "0000001110000000001011111000000100",
			2734 => "00000000111111100010101011100101",
			2735 => "00000000000000000010101011100101",
			2736 => "0000000100000000001011110000001100",
			2737 => "0000000001000000000001111000000100",
			2738 => "00000000000000000010101011100101",
			2739 => "0000000111000000000110100100000100",
			2740 => "00000000000000000010101011100101",
			2741 => "11111111101110110010101011100101",
			2742 => "0000001110000000001111100100000100",
			2743 => "00000000000010110010101011100101",
			2744 => "00000000000000000010101011100101",
			2745 => "0000000001000000000001000100000100",
			2746 => "11111110011011010010101100111001",
			2747 => "0000001110000000000110010000001000",
			2748 => "0000001011000000000000011100000100",
			2749 => "00000001100101000010101100111001",
			2750 => "00000000000000000010101100111001",
			2751 => "0000000100000000001100111000001100",
			2752 => "0000000100000000000110101100000100",
			2753 => "11111110001111000010101100111001",
			2754 => "0000000011000000001100000000000100",
			2755 => "00000000011001110010101100111001",
			2756 => "11111110101111000010101100111001",
			2757 => "0000001110000000001011111000010000",
			2758 => "0000000001000000000111101000000100",
			2759 => "11111110111000010010101100111001",
			2760 => "0000000100000000000010010100001000",
			2761 => "0000001110000000001111010100000100",
			2762 => "00000001010010100010101100111001",
			2763 => "11111110100110010010101100111001",
			2764 => "00000001110011100010101100111001",
			2765 => "11111110100111110010101100111001",
			2766 => "0000000001000000000001000100000100",
			2767 => "11111110010111010010101110010101",
			2768 => "0000001101000000001111010000011000",
			2769 => "0000001000000000000001110000010100",
			2770 => "0000000010000000001101101100010000",
			2771 => "0000001100000000001011000000001100",
			2772 => "0000000010000000001100111000001000",
			2773 => "0000000011000000001000001100000100",
			2774 => "00000010110110110010101110010101",
			2775 => "00000001001101000010101110010101",
			2776 => "00000100001010100010101110010101",
			2777 => "00000001001101000010101110010101",
			2778 => "00000111010110100010101110010101",
			2779 => "11111110001101100010101110010101",
			2780 => "0000000101000000000110100000001000",
			2781 => "0000000000000000001000110000000100",
			2782 => "00000011111001000010101110010101",
			2783 => "11111111001100000010101110010101",
			2784 => "0000001110000000001111010100001000",
			2785 => "0000000001000000000111101000000100",
			2786 => "11111110010010110010101110010101",
			2787 => "00000010101010000010101110010101",
			2788 => "11111110010111100010101110010101",
			2789 => "0000001000000000000001110000101100",
			2790 => "0000000100000000001000000100011100",
			2791 => "0000001110000000000111010100011000",
			2792 => "0000000001000000001011111100001000",
			2793 => "0000001001000000001001111100000100",
			2794 => "11111110101101110010101111110001",
			2795 => "00000000000000000010101111110001",
			2796 => "0000000100000000000001011100001100",
			2797 => "0000000101000000000010110100000100",
			2798 => "00000001000111010010101111110001",
			2799 => "0000001110000000000110010000000100",
			2800 => "00000000101011100010101111110001",
			2801 => "11111111001101010010101111110001",
			2802 => "00000001010011110010101111110001",
			2803 => "11111110100100100010101111110001",
			2804 => "0000000101000000000001000000001100",
			2805 => "0000000001000000000001000100000100",
			2806 => "00000000000000000010101111110001",
			2807 => "0000001110000000001111100100000100",
			2808 => "00000001101100110010101111110001",
			2809 => "00000000000000000010101111110001",
			2810 => "11111111001011110010101111110001",
			2811 => "11111110011100100010101111110001",
			2812 => "0000001000000000000001110000111000",
			2813 => "0000001110000000001110110100011000",
			2814 => "0000000010000000000010000100001100",
			2815 => "0000000000000000001011010100001000",
			2816 => "0000000001000000001011111100000100",
			2817 => "11111111111010000010110001100101",
			2818 => "00000000001010010010110001100101",
			2819 => "11111111001010100010110001100101",
			2820 => "0000000011000000001100000000001000",
			2821 => "0000000001000000000001000100000100",
			2822 => "00000000000000000010110001100101",
			2823 => "00000001011010100010110001100101",
			2824 => "00000000000000000010110001100101",
			2825 => "0000000001000000001101111100010000",
			2826 => "0000001101000000001100100100000100",
			2827 => "00000000000000000010110001100101",
			2828 => "0000000111000000000001101000001000",
			2829 => "0000000110000000001011001100000100",
			2830 => "00000000000000000010110001100101",
			2831 => "11111110100100010010110001100101",
			2832 => "00000000000000000010110001100101",
			2833 => "0000001101000000000101001000001000",
			2834 => "0000000010000000001000001100000100",
			2835 => "00000000000000000010110001100101",
			2836 => "00000001001000000010110001100101",
			2837 => "0000001110000000000111010100000100",
			2838 => "00000000000000000010110001100101",
			2839 => "11111111001110010010110001100101",
			2840 => "11111110011111010010110001100101",
			2841 => "0000000001000000001011111100001000",
			2842 => "0000001001000000001001111100000100",
			2843 => "11111110100000010010110011101001",
			2844 => "00000000000000000010110011101001",
			2845 => "0000001111000000000000010000011100",
			2846 => "0000000100000000001111100100001100",
			2847 => "0000000011000000001110110100000100",
			2848 => "00000000101101000010110011101001",
			2849 => "0000001100000000000100011000000100",
			2850 => "11111110110000100010110011101001",
			2851 => "00000000000000000010110011101001",
			2852 => "0000001100000000001011000000001000",
			2853 => "0000000011000000001010000100000100",
			2854 => "00000001011000100010110011101001",
			2855 => "00000000000000000010110011101001",
			2856 => "0000001001000000000111101100000100",
			2857 => "11111111101101010010110011101001",
			2858 => "00000000000010010010110011101001",
			2859 => "0000001001000000000000001000001000",
			2860 => "0000001011000000000111010000000100",
			2861 => "00000000000000000010110011101001",
			2862 => "11111110100001100010110011101001",
			2863 => "0000001101000000000101001000001000",
			2864 => "0000000000000000000111000000000100",
			2865 => "00000001000110010010110011101001",
			2866 => "00000000000000000010110011101001",
			2867 => "0000001001000000001010100000001000",
			2868 => "0000001011000000000110110100000100",
			2869 => "00000000000000000010110011101001",
			2870 => "00000000001011100010110011101001",
			2871 => "0000001011000000000000011100000100",
			2872 => "00000000000000000010110011101001",
			2873 => "11111111000100010010110011101001",
			2874 => "0000001001000000000101010000000100",
			2875 => "11111110011010000010110101010101",
			2876 => "0000001110000000001111010100011000",
			2877 => "0000001110000000000110010000000100",
			2878 => "00000001101000110010110101010101",
			2879 => "0000000100000000001111100100000100",
			2880 => "11111101111100100010110101010101",
			2881 => "0000001001000000000111101100000100",
			2882 => "11111110110011010010110101010101",
			2883 => "0000000110000000001111000000001000",
			2884 => "0000001001000000000111101100000100",
			2885 => "00000000001111100010110101010101",
			2886 => "00000001101100010010110101010101",
			2887 => "00000000010110110010110101010101",
			2888 => "0000001100000000000100011000010000",
			2889 => "0000000100000000000010010100000100",
			2890 => "11111110011010100010110101010101",
			2891 => "0000001110000000001011111000001000",
			2892 => "0000000010000000001100111000000100",
			2893 => "00000000011000010010110101010101",
			2894 => "00000001110110010010110101010101",
			2895 => "11111110110110100010110101010101",
			2896 => "0000001111000000001111100100001000",
			2897 => "0000000110000000001001100100000100",
			2898 => "11111111111011010010110101010101",
			2899 => "00000000000000000010110101010101",
			2900 => "11111110011011110010110101010101",
			2901 => "0000001000000000000001110000110000",
			2902 => "0000000100000000001000000100100000",
			2903 => "0000001110000000001010000100011100",
			2904 => "0000000010000000000111010100010100",
			2905 => "0000001110000000000010000100010000",
			2906 => "0000000110000000001010011000001000",
			2907 => "0000000010000000000010000100000100",
			2908 => "11111111001100010010110110111001",
			2909 => "00000000000000000010110110111001",
			2910 => "0000000111000000001110110000000100",
			2911 => "00000000000000000010110110111001",
			2912 => "00000000110101000010110110111001",
			2913 => "11111110110100110010110110111001",
			2914 => "0000000101000000001101000100000100",
			2915 => "00000001001110110010110110111001",
			2916 => "00000000000000000010110110111001",
			2917 => "11111110111000110010110110111001",
			2918 => "0000001101000000000111111100001100",
			2919 => "0000000110000000001101011000000100",
			2920 => "00000000000000000010110110111001",
			2921 => "0000001110000000001111100100000100",
			2922 => "00000001101110100010110110111001",
			2923 => "00000000000000000010110110111001",
			2924 => "11111111110111110010110110111001",
			2925 => "11111110100011000010110110111001",
			2926 => "0000001000000000000001110000111000",
			2927 => "0000000100000000001000000100101000",
			2928 => "0000001000000000000110011100011100",
			2929 => "0000001101000000001100100100001000",
			2930 => "0000001001000000000101010000000100",
			2931 => "00000000000000000010111000101101",
			2932 => "00000000101110000010111000101101",
			2933 => "0000000100000000001111100100001000",
			2934 => "0000001110000000000010000000000100",
			2935 => "00000000000000000010111000101101",
			2936 => "11111111001101110010111000101101",
			2937 => "0000000011000000001111010100000100",
			2938 => "00000000101101110010111000101101",
			2939 => "0000001010000000000111110100000100",
			2940 => "11111111101001010010111000101101",
			2941 => "00000000000000000010111000101101",
			2942 => "0000001001000000000000001000001000",
			2943 => "0000000101000000001110101000000100",
			2944 => "11111110110001100010111000101101",
			2945 => "00000000000000000010111000101101",
			2946 => "00000000000000000010111000101101",
			2947 => "0000000101000000000001000000001100",
			2948 => "0000001001000000000101010000000100",
			2949 => "00000000000000000010111000101101",
			2950 => "0000001110000000001111100100000100",
			2951 => "00000001001101100010111000101101",
			2952 => "00000000000000000010111000101101",
			2953 => "00000000000000000010111000101101",
			2954 => "11111110110011000010111000101101",
			2955 => "0000001001000000000101010000000100",
			2956 => "11111110011000010010111010000001",
			2957 => "0000001110000000001011111000100100",
			2958 => "0000001101000000001001010000011100",
			2959 => "0000000010000000001101101100011000",
			2960 => "0000001101000000001111010000010000",
			2961 => "0000000011000000001100010000001000",
			2962 => "0000001000000000000110011000000100",
			2963 => "00000011000001100010111010000001",
			2964 => "00000010001100110010111010000001",
			2965 => "0000000100000000001011101100000100",
			2966 => "11111101011001000010111010000001",
			2967 => "00000010000111010010111010000001",
			2968 => "0000000001000000000001111000000100",
			2969 => "11111110011010100010111010000001",
			2970 => "00000001010011010010111010000001",
			2971 => "00000100011100000010111010000001",
			2972 => "0000001111000000001011101100000100",
			2973 => "11111110011011100010111010000001",
			2974 => "00000010011010110010111010000001",
			2975 => "11111110011000100010111010000001",
			2976 => "0000000001000000000001000100000100",
			2977 => "11111110101011110010111011111101",
			2978 => "0000000100000000000010010100101100",
			2979 => "0000001111000000000000010000100000",
			2980 => "0000000100000000001111100100001100",
			2981 => "0000000011000000001110110100000100",
			2982 => "00000000010010110010111011111101",
			2983 => "0000000111000000000001101000000100",
			2984 => "11111111001101010010111011111101",
			2985 => "00000000000000000010111011111101",
			2986 => "0000001100000000001011000000001000",
			2987 => "0000000011000000001000001100000100",
			2988 => "00000001000010010010111011111101",
			2989 => "00000000000000000010111011111101",
			2990 => "0000000000000000001111001000001000",
			2991 => "0000000011000000001010000100000100",
			2992 => "00000000001110000010111011111101",
			2993 => "00000000000000000010111011111101",
			2994 => "11111111100111100010111011111101",
			2995 => "0000000100000000000010010100001000",
			2996 => "0000001001000000001010100100000100",
			2997 => "11111110110111100010111011111101",
			2998 => "00000000000000000010111011111101",
			2999 => "00000000000000000010111011111101",
			3000 => "0000000011000000001111100100001000",
			3001 => "0000000110000000001000010000000100",
			3002 => "00000001011001000010111011111101",
			3003 => "00000000000000000010111011111101",
			3004 => "0000001000000000000101000100000100",
			3005 => "00000000000000000010111011111101",
			3006 => "11111111100001010010111011111101",
			3007 => "0000000001000000001011111100001000",
			3008 => "0000001001000000001001111100000100",
			3009 => "11111110100100000010111110001001",
			3010 => "00000000000000000010111110001001",
			3011 => "0000000111000000001001001000010000",
			3012 => "0000000011000000001011111000001100",
			3013 => "0000001001000000001010100000001000",
			3014 => "0000001100000000001101111000000100",
			3015 => "00000000000000000010111110001001",
			3016 => "00000001101000110010111110001001",
			3017 => "00000000000000000010111110001001",
			3018 => "00000000000000000010111110001001",
			3019 => "0000000001000000000001111000010000",
			3020 => "0000001110000000000110010000000100",
			3021 => "00000000010010110010111110001001",
			3022 => "0000001001000000000111101100001000",
			3023 => "0000000111000000001000011000000100",
			3024 => "11111110111011110010111110001001",
			3025 => "00000000000000000010111110001001",
			3026 => "00000000000000000010111110001001",
			3027 => "0000001101000000000101001000001100",
			3028 => "0000000010000000001111010100000100",
			3029 => "00000000000000000010111110001001",
			3030 => "0000001110000000001011111000000100",
			3031 => "00000001001001110010111110001001",
			3032 => "00000000000000000010111110001001",
			3033 => "0000001100000000000100011000001100",
			3034 => "0000001001000000000000001000000100",
			3035 => "00000000000000000010111110001001",
			3036 => "0000000110000000000100111100000100",
			3037 => "00000000101011100010111110001001",
			3038 => "00000000000000000010111110001001",
			3039 => "0000001001000000000000001000000100",
			3040 => "00000000000000000010111110001001",
			3041 => "11111111001110010010111110001001",
			3042 => "0000001000000000000001110000111100",
			3043 => "0000000100000000000010010100101000",
			3044 => "0000001110000000000110111100100000",
			3045 => "0000000100000000001100111000010100",
			3046 => "0000001110000000000110010000001100",
			3047 => "0000000110000000001010011000000100",
			3048 => "00000000000000000011000000000101",
			3049 => "0000001101000000000000110100000100",
			3050 => "00000000000000000011000000000101",
			3051 => "00000000101100000011000000000101",
			3052 => "0000001111000000001010000100000100",
			3053 => "11111110111110110011000000000101",
			3054 => "00000000000000000011000000000101",
			3055 => "0000000001000000001110010100000100",
			3056 => "00000000000000000011000000000101",
			3057 => "0000001000000000001010110000000100",
			3058 => "00000000000000000011000000000101",
			3059 => "00000001001001100011000000000101",
			3060 => "0000000001000000001101111100000100",
			3061 => "11111110100110110011000000000101",
			3062 => "00000000000000000011000000000101",
			3063 => "0000001101000000000111111100010000",
			3064 => "0000000001000000000001000100000100",
			3065 => "00000000000000000011000000000101",
			3066 => "0000000110000000000100111100001000",
			3067 => "0000001110000000001011111000000100",
			3068 => "00000001101010100011000000000101",
			3069 => "00000000000000000011000000000101",
			3070 => "00000000000000000011000000000101",
			3071 => "11111111110010010011000000000101",
			3072 => "11111110100100110011000000000101",
			3073 => "0000000001000000000001000100000100",
			3074 => "11111110011010110011000010010001",
			3075 => "0000000111000000001001001000011000",
			3076 => "0000000100000000001101101100001100",
			3077 => "0000000011000000001100010000000100",
			3078 => "00000001011101100011000010010001",
			3079 => "0000000100000000001011101100000100",
			3080 => "11111110011110010011000010010001",
			3081 => "00000000000000000011000010010001",
			3082 => "0000001110000000001011111000001000",
			3083 => "0000000100000000000010110000000100",
			3084 => "00000001100010010011000010010001",
			3085 => "00000011000001100011000010010001",
			3086 => "11111111100101110011000010010001",
			3087 => "0000001110000000000110111100010100",
			3088 => "0000001010000000000011101000001000",
			3089 => "0000000011000000001100010000000100",
			3090 => "00000000010001110011000010010001",
			3091 => "11111110011101110011000010010001",
			3092 => "0000001001000000000100101100000100",
			3093 => "11111111000101110011000010010001",
			3094 => "0000000000000000000110001000000100",
			3095 => "00000000000000110011000010010001",
			3096 => "00000001100100110011000010010001",
			3097 => "0000000011000000000111010100000100",
			3098 => "11111101110010110011000010010001",
			3099 => "0000000101000000001100100100010000",
			3100 => "0000000111000000000110100100001000",
			3101 => "0000000011000000001111100100000100",
			3102 => "00000000100001000011000010010001",
			3103 => "00000000000000000011000010010001",
			3104 => "0000000111000000000001101000000100",
			3105 => "11111111001111110011000010010001",
			3106 => "00000000000000000011000010010001",
			3107 => "11111110100110010011000010010001",
			3108 => "0000000001000000000001000100000100",
			3109 => "11111110011001100011000011101101",
			3110 => "0000001110000000001011111000101000",
			3111 => "0000000011000000001100010000000100",
			3112 => "00000001101101000011000011101101",
			3113 => "0000000100000000001011101100001100",
			3114 => "0000001111000000000110111100001000",
			3115 => "0000001110000000001110110100000100",
			3116 => "00000000000011010011000011101101",
			3117 => "11111110110001000011000011101101",
			3118 => "11111101100100000011000011101101",
			3119 => "0000000001000000000111101000001000",
			3120 => "0000001110000000001111010100000100",
			3121 => "11111111100011010011000011101101",
			3122 => "11111110000111100011000011101101",
			3123 => "0000000100000000000011000000001000",
			3124 => "0000001010000000000111110100000100",
			3125 => "00000000111001010011000011101101",
			3126 => "11111100100110110011000011101101",
			3127 => "0000000010000000001101101100000100",
			3128 => "00000001101010010011000011101101",
			3129 => "00000010101100110011000011101101",
			3130 => "11111110011011010011000011101101",
			3131 => "0000001001000000000101010000000100",
			3132 => "11111110011000100011000101011001",
			3133 => "0000001110000000001011111000110000",
			3134 => "0000001100000000001011000000011100",
			3135 => "0000000010000000001101101100011000",
			3136 => "0000001101000000001111010000010000",
			3137 => "0000001110000000000110111100001000",
			3138 => "0000000100000000001011101100000100",
			3139 => "00000001101010100011000101011001",
			3140 => "00000010000001010011000101011001",
			3141 => "0000000100000000000011000000000100",
			3142 => "11111101100111110011000101011001",
			3143 => "00000001100101100011000101011001",
			3144 => "0000000100000000000011000000000100",
			3145 => "11111110011100110011000101011001",
			3146 => "00000000110001100011000101011001",
			3147 => "00000100010011000011000101011001",
			3148 => "0000001100000000001000000000001000",
			3149 => "0000001001000000000111101100000100",
			3150 => "11111100101010010011000101011001",
			3151 => "00000000011100100011000101011001",
			3152 => "0000001101000000001001010000000100",
			3153 => "00000010001100000011000101011001",
			3154 => "0000000001000000000001111000000100",
			3155 => "11111110011110010011000101011001",
			3156 => "00000000010110010011000101011001",
			3157 => "11111110011001000011000101011001",
			3158 => "0000000001000000000001000100000100",
			3159 => "11111110011010100011000111110101",
			3160 => "0000000111000000001001001000011100",
			3161 => "0000000100000000000011001100010100",
			3162 => "0000000011000000001100010000000100",
			3163 => "00000001100100110011000111110101",
			3164 => "0000000100000000001011101100000100",
			3165 => "11111110011000010011000111110101",
			3166 => "0000001110000000001011111000001000",
			3167 => "0000000100000000001101101100000100",
			3168 => "00000000000000000011000111110101",
			3169 => "00000001011110100011000111110101",
			3170 => "11111111110010000011000111110101",
			3171 => "0000001111000000001110000000000100",
			3172 => "00000011101000010011000111110101",
			3173 => "00000000000000000011000111110101",
			3174 => "0000001110000000000110111100010000",
			3175 => "0000001010000000000011101000001000",
			3176 => "0000000011000000001100010000000100",
			3177 => "00000000010101000011000111110101",
			3178 => "11111110011010110011000111110101",
			3179 => "0000000001000000000111101000000100",
			3180 => "11111111110111010011000111110101",
			3181 => "00000001100000010011000111110101",
			3182 => "0000001100000000000100011000010000",
			3183 => "0000000111000000000110100100001000",
			3184 => "0000000011000000001111100100000100",
			3185 => "00000000101001010011000111110101",
			3186 => "00000000000000000011000111110101",
			3187 => "0000001100000000000100011000000100",
			3188 => "11111110111100000011000111110101",
			3189 => "00000000000000000011000111110101",
			3190 => "0000001011000000000000011100000100",
			3191 => "11111101101010100011000111110101",
			3192 => "0000000011000000001000001100001000",
			3193 => "0000000101000000001100100100000100",
			3194 => "00000000001111000011000111110101",
			3195 => "00000000000000000011000111110101",
			3196 => "11111110100101100011000111110101",
			3197 => "0000001000000000000001110000111100",
			3198 => "0000000110000000001010011000000100",
			3199 => "11111110101001110011001001110001",
			3200 => "0000001110000000001100010000011000",
			3201 => "0000001110000000000110010000001000",
			3202 => "0000001110000000000101001000000100",
			3203 => "00000000000000000011001001110001",
			3204 => "00000001101010110011001001110001",
			3205 => "0000000010000000001010000100001100",
			3206 => "0000000011000000001100010000001000",
			3207 => "0000001010000000000011101000000100",
			3208 => "00000001001010110011001001110001",
			3209 => "00000000000000000011001001110001",
			3210 => "11111110101110100011001001110001",
			3211 => "00000001100101000011001001110001",
			3212 => "0000000100000000000011000000010000",
			3213 => "0000001010000000000111110100001100",
			3214 => "0000001010000000000011101000000100",
			3215 => "11111110010100100011001001110001",
			3216 => "0000001000000000001100011100000100",
			3217 => "00000000100110110011001001110001",
			3218 => "11111111000101110011001001110001",
			3219 => "11111101000011110011001001110001",
			3220 => "0000001110000000001011111000001100",
			3221 => "0000000100000000000010010100001000",
			3222 => "0000000011000000000111010100000100",
			3223 => "00000001010011100011001001110001",
			3224 => "11111110111101010011001001110001",
			3225 => "00000001011111110011001001110001",
			3226 => "11111110100011100011001001110001",
			3227 => "11111110011010010011001001110001",
			3228 => "0000000001000000000001000100000100",
			3229 => "11111110110101010011001011111101",
			3230 => "0000001110000000000110010000001000",
			3231 => "0000001111000000001000001100000100",
			3232 => "00000000111011010011001011111101",
			3233 => "00000000000000000011001011111101",
			3234 => "0000000001000000000111101000001100",
			3235 => "0000001101000000001101000100000100",
			3236 => "00000000000000000011001011111101",
			3237 => "0000001001000000000111101100000100",
			3238 => "11111110111100100011001011111101",
			3239 => "00000000000000000011001011111101",
			3240 => "0000000111000000000110100100011000",
			3241 => "0000001100000000001010111000001100",
			3242 => "0000000011000000000111011000000100",
			3243 => "00000000000000000011001011111101",
			3244 => "0000001101000000001100100100000100",
			3245 => "00000000000000000011001011111101",
			3246 => "11111111101110110011001011111101",
			3247 => "0000000110000000000100111100001000",
			3248 => "0000000011000000001011111000000100",
			3249 => "00000001000000100011001011111101",
			3250 => "00000000000000000011001011111101",
			3251 => "00000000000000000011001011111101",
			3252 => "0000000111000000000001101000001100",
			3253 => "0000001100000000001010111000000100",
			3254 => "00000000000000000011001011111101",
			3255 => "0000001011000000000110110100000100",
			3256 => "11111111000001000011001011111101",
			3257 => "00000000000000000011001011111101",
			3258 => "0000001111000000001100111000001000",
			3259 => "0000000111000000001000011000000100",
			3260 => "00000000001110110011001011111101",
			3261 => "00000000000000000011001011111101",
			3262 => "00000000000000000011001011111101",
			3263 => "0000000001000000000001000100000100",
			3264 => "11111110011100000011001110110011",
			3265 => "0000001110000000000110010000001000",
			3266 => "0000001011000000000000011100000100",
			3267 => "00000001100000110011001110110011",
			3268 => "00000000000000000011001110110011",
			3269 => "0000001100000000001010111000011100",
			3270 => "0000000101000000000010110100001100",
			3271 => "0000000001000000000111101000000100",
			3272 => "11111111100101110011001110110011",
			3273 => "0000001000000000001100000100000100",
			3274 => "00000000110101000011001110110011",
			3275 => "00000000000000000011001110110011",
			3276 => "0000000001000000000001111000001000",
			3277 => "0000001101000000000101001000000100",
			3278 => "11111110010101100011001110110011",
			3279 => "00000000000000000011001110110011",
			3280 => "0000001001000000000000001000000100",
			3281 => "00000000000000000011001110110011",
			3282 => "11111111101100100011001110110011",
			3283 => "0000000111000000000001101000100000",
			3284 => "0000001010000000000011101000010000",
			3285 => "0000001101000000001110000100001000",
			3286 => "0000000111000000001001001000000100",
			3287 => "00000000000000000011001110110011",
			3288 => "00000000110000100011001110110011",
			3289 => "0000001011000000000101100100000100",
			3290 => "11111111010100000011001110110011",
			3291 => "00000000000000000011001110110011",
			3292 => "0000001100000000001011000000001000",
			3293 => "0000001110000000001000001100000100",
			3294 => "00000001100101010011001110110011",
			3295 => "00000000000000000011001110110011",
			3296 => "0000001100000000001000000000000100",
			3297 => "11111111011011100011001110110011",
			3298 => "00000000000000000011001110110011",
			3299 => "0000001100000000000100011000001100",
			3300 => "0000001010000000000011101000000100",
			3301 => "00000000000000000011001110110011",
			3302 => "0000001000000000000001010100000100",
			3303 => "00000001000000000011001110110011",
			3304 => "00000000000000000011001110110011",
			3305 => "0000001000000000001100011100000100",
			3306 => "00000000000000000011001110110011",
			3307 => "11111110011110100011001110110011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1096, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(2190, initial_addr_3'length));
	end generate gen_rom_11;

	gen_rom_12: if SELECT_ROM = 12 generate
		bank <= (
			0 => "00000000000000000000000000000101",
			1 => "00000000000000000000000000001001",
			2 => "00000000000000000000000000001101",
			3 => "00000000000000000000000000010001",
			4 => "00000000000000000000000000010101",
			5 => "00000000000000000000000000011001",
			6 => "00000000000000000000000000011101",
			7 => "00000000000000000000000000100001",
			8 => "00000000000000000000000000100101",
			9 => "00000000000000000000000000101001",
			10 => "00000000000000000000000000101101",
			11 => "00000000000000000000000000110001",
			12 => "00000000000000000000000000110101",
			13 => "00000000000000000000000000111001",
			14 => "00000000000000000000000000111101",
			15 => "00000000000000000000000001000001",
			16 => "00000000000000000000000001000101",
			17 => "00000000000000000000000001001001",
			18 => "00000000000000000000000001001101",
			19 => "00000000000000000000000001010001",
			20 => "00000000000000000000000001010101",
			21 => "00000000000000000000000001011001",
			22 => "00000000000000000000000001011101",
			23 => "00000000000000000000000001100001",
			24 => "00000000000000000000000001100101",
			25 => "00000000000000000000000001101001",
			26 => "00000000000000000000000001101101",
			27 => "00000000000000000000000001110001",
			28 => "00000000000000000000000001110101",
			29 => "0000000100000000000001001100000100",
			30 => "11111111111110100000000010000001",
			31 => "00000000000000000000000010000001",
			32 => "0000000100000000000011011000000100",
			33 => "11111111111110110000000010001101",
			34 => "00000000000000000000000010001101",
			35 => "0000000100000000000100111000000100",
			36 => "11111111111001110000000010011001",
			37 => "00000000000000000000000010011001",
			38 => "0000000100000000000011111000000100",
			39 => "11111111111011000000000010100101",
			40 => "00000000000000000000000010100101",
			41 => "0000000100000000000100111000000100",
			42 => "11111111111000100000000010110001",
			43 => "00000000000000000000000010110001",
			44 => "0000000001000000001111001100000100",
			45 => "11111111111011010000000010111101",
			46 => "00000000000000000000000010111101",
			47 => "0000000100000000000011111000000100",
			48 => "11111111111110000000000011001001",
			49 => "00000000000000000000000011001001",
			50 => "0000000100000000000000010100000100",
			51 => "11111111111100000000000011011101",
			52 => "0000000100000000001010010000000100",
			53 => "00000000000001010000000011011101",
			54 => "00000000000000000000000011011101",
			55 => "0000000100000000000101100000001000",
			56 => "0000001001000000001010011000000100",
			57 => "11111111101011100000000011110001",
			58 => "00000000000000000000000011110001",
			59 => "00000000000000000000000011110001",
			60 => "0000000010000000000110101100000100",
			61 => "11111111111101100000000100000101",
			62 => "0000000010000000001101101100000100",
			63 => "00000000000010110000000100000101",
			64 => "00000000000000000000000100000101",
			65 => "0000000010000000001011111000000100",
			66 => "00000000000000000000000100011001",
			67 => "0000000010000000001101101100000100",
			68 => "00000000001101010000000100011001",
			69 => "00000000000000000000000100011001",
			70 => "0000000010000000000110101100000100",
			71 => "11111111111011110000000100101101",
			72 => "0000000010000000001111101000000100",
			73 => "00000000001101100000000100101101",
			74 => "00000000000000000000000100101101",
			75 => "0000000100000000000100111000001000",
			76 => "0000001001000000001010011000000100",
			77 => "11111111110101100000000101000001",
			78 => "00000000000000000000000101000001",
			79 => "00000000000000000000000101000001",
			80 => "0000000001000000001101011100001000",
			81 => "0000000010000000001011101100000100",
			82 => "11111111110110100000000101010101",
			83 => "00000000000000000000000101010101",
			84 => "00000000000000000000000101010101",
			85 => "0000000010000000001011111000001100",
			86 => "0000000110000000001001100100001000",
			87 => "0000000001000000000000111100000100",
			88 => "11111111101100010000000101110001",
			89 => "00000000000000000000000101110001",
			90 => "00000000000000000000000101110001",
			91 => "00000000000000000000000101110001",
			92 => "0000001110000000000111110000001100",
			93 => "0000000100000000001001000000000100",
			94 => "00000000000000000000000110001101",
			95 => "0000000100000000001010010000000100",
			96 => "00000000000100010000000110001101",
			97 => "00000000000000000000000110001101",
			98 => "11111111111111010000000110001101",
			99 => "0000000100000000000010100100000100",
			100 => "11111111111101100000000110101001",
			101 => "0000000010000000000000010000000100",
			102 => "00000000000000000000000110101001",
			103 => "0000000010000000001111101000000100",
			104 => "00000000000101000000000110101001",
			105 => "00000000000000000000000110101001",
			106 => "0000000001000000001101011100001100",
			107 => "0000000010000000001011101100001000",
			108 => "0000001001000000001101011000000100",
			109 => "11111111110011000000000111000101",
			110 => "00000000000000000000000111000101",
			111 => "00000000000000000000000111000101",
			112 => "00000000000000000000000111000101",
			113 => "0000000001000000001101011100001000",
			114 => "0000000010000000001011101100000100",
			115 => "11111111101100110000000111101001",
			116 => "00000000000000000000000111101001",
			117 => "0000000101000000000111110000001000",
			118 => "0000000100000000001110111000000100",
			119 => "00000000000000000000000111101001",
			120 => "00000000001001110000000111101001",
			121 => "00000000000000000000000111101001",
			122 => "0000000001000000001101101000000100",
			123 => "11111111101100010000001000001101",
			124 => "0000001110000000001110101100001100",
			125 => "0000000110000000001011001100001000",
			126 => "0000000111000000000111001000000100",
			127 => "00000000001011110000001000001101",
			128 => "00000000000000000000001000001101",
			129 => "00000000000000000000001000001101",
			130 => "00000000000000000000001000001101",
			131 => "0000000100000000000011010100000100",
			132 => "11111111111101000000001000110001",
			133 => "0000000010000000000110101100000100",
			134 => "00000000000000000000001000110001",
			135 => "0000000010000000000011000000001000",
			136 => "0000000100000000001010010000000100",
			137 => "00000000010001100000001000110001",
			138 => "00000000000000000000001000110001",
			139 => "00000000000000000000001000110001",
			140 => "0000000100000000000011011000000100",
			141 => "11111111110111100000001001010101",
			142 => "0000001101000000000100010000001100",
			143 => "0000001110000000000110000100000100",
			144 => "00000000000000000000001001010101",
			145 => "0000001101000000001000011000000100",
			146 => "00000000000000000000001001010101",
			147 => "00000000001001010000001001010101",
			148 => "00000000000000000000001001010101",
			149 => "0000000001000000001011101000001000",
			150 => "0000000100000000000011111000000100",
			151 => "11111111100001110000001010000001",
			152 => "00000000000000000000001010000001",
			153 => "0000001110000000001001010100001100",
			154 => "0000000111000000001101111000000100",
			155 => "00000000000000000000001010000001",
			156 => "0000000001000000001111001100000100",
			157 => "00000000000000000000001010000001",
			158 => "00000000011100010000001010000001",
			159 => "00000000000000000000001010000001",
			160 => "0000000001000000001111001100001000",
			161 => "0000000100000000000100111000000100",
			162 => "11111111100110010000001010101101",
			163 => "00000000000000000000001010101101",
			164 => "0000001110000000000111110000001100",
			165 => "0000000111000000001101111000000100",
			166 => "00000000000000000000001010101101",
			167 => "0000000110000000001001100100000100",
			168 => "00000000010011010000001010101101",
			169 => "00000000000000000000001010101101",
			170 => "00000000000000000000001010101101",
			171 => "0000000010000000000110101100001100",
			172 => "0000000000000000000011111100000100",
			173 => "00000000000000000000001011100001",
			174 => "0000001100000000001110001100000100",
			175 => "11111111010111100000001011100001",
			176 => "00000000000000000000001011100001",
			177 => "0000001111000000001100010000001100",
			178 => "0000001010000000000001110000001000",
			179 => "0000001100000000000011011100000100",
			180 => "00000000000000000000001011100001",
			181 => "00000000100110100000001011100001",
			182 => "00000000000000000000001011100001",
			183 => "00000000000000000000001011100001",
			184 => "0000000100000000000011110100000100",
			185 => "11111111010111010000001100010101",
			186 => "0000001011000000000011100000001100",
			187 => "0000000001000000001111001100000100",
			188 => "00000000000000000000001100010101",
			189 => "0000000111000000001101111000000100",
			190 => "00000000000000000000001100010101",
			191 => "00000000101010000000001100010101",
			192 => "0000001000000000001011010100000100",
			193 => "00000000000000000000001100010101",
			194 => "0000001110000000000111110000000100",
			195 => "00000000000000000000001100010101",
			196 => "11111111100011000000001100010101",
			197 => "0000001001000000000001111000001000",
			198 => "0000000010000000001011101100000100",
			199 => "11111111100011110000001101001001",
			200 => "00000000000000000000001101001001",
			201 => "0000001110000000001001010100010000",
			202 => "0000001100000000001100110000000100",
			203 => "00000000000000000000001101001001",
			204 => "0000000010000000000111011000000100",
			205 => "00000000000000000000001101001001",
			206 => "0000000110000000001111000000000100",
			207 => "00000000010110000000001101001001",
			208 => "00000000000000000000001101001001",
			209 => "00000000000000000000001101001001",
			210 => "0000001001000000001011111100000100",
			211 => "11111111101011100000001101110101",
			212 => "0000001110000000001110101100010000",
			213 => "0000000110000000001011001100001100",
			214 => "0000001011000000000001111100000100",
			215 => "00000000000000000000001101110101",
			216 => "0000001111000000000001000000000100",
			217 => "00000000000000000000001101110101",
			218 => "00000000001100100000001101110101",
			219 => "00000000000000000000001101110101",
			220 => "00000000000000000000001101110101",
			221 => "0000000010000000001000001100001100",
			222 => "0000000111000000001100101000001000",
			223 => "0000001100000000001110001100000100",
			224 => "11111110110001110000001110111001",
			225 => "00000000000000000000001110111001",
			226 => "00000000000000000000001110111001",
			227 => "0000001111000000000010000000010000",
			228 => "0000001000000000001010101100001100",
			229 => "0000001110000000000111110000001000",
			230 => "0000000001000000001011101000000100",
			231 => "00000000000000000000001110111001",
			232 => "00000000111111010000001110111001",
			233 => "00000000000000000000001110111001",
			234 => "00000000000000000000001110111001",
			235 => "0000001110000000001110101100000100",
			236 => "00000000000000000000001110111001",
			237 => "11111111100110000000001110111001",
			238 => "0000000100000000000011010100000100",
			239 => "11111111000010000000001111110101",
			240 => "0000000001000000001111001100001000",
			241 => "0000000100000000000101100000000100",
			242 => "11111111100011000000001111110101",
			243 => "00000000000000000000001111110101",
			244 => "0000000110000000001011001100001100",
			245 => "0000000011000000001101000100001000",
			246 => "0000001010000000001010110000000100",
			247 => "00000000010111010000001111110101",
			248 => "00000000000000000000001111110101",
			249 => "11111111111110000000001111110101",
			250 => "0000001110000000001110101000000100",
			251 => "00000000110011010000001111110101",
			252 => "00000000000000000000001111110101",
			253 => "0000000100000000000011010100000100",
			254 => "00000000000000000000010000101001",
			255 => "0000000110000000001001100100010100",
			256 => "0000000001000000000110101000000100",
			257 => "00000000000000000000010000101001",
			258 => "0000000011000000001101000100001100",
			259 => "0000001111000000000010000000001000",
			260 => "0000000111000000000110000100000100",
			261 => "00000000000000000000010000101001",
			262 => "00000000011000000000010000101001",
			263 => "00000000000000000000010000101001",
			264 => "00000000000000000000010000101001",
			265 => "00000000000000000000010000101001",
			266 => "0000000100000000000011010100000100",
			267 => "11111111000101000000010001101101",
			268 => "0000000001000000001111001100001000",
			269 => "0000000100000000000101100000000100",
			270 => "11111111100101110000010001101101",
			271 => "00000000000000000000010001101101",
			272 => "0000000110000000001011001100010000",
			273 => "0000001111000000001100010100001000",
			274 => "0000001010000000001010110000000100",
			275 => "00000000001011110000010001101101",
			276 => "00000000000000000000010001101101",
			277 => "0000001010000000000110011000000100",
			278 => "00000000000000000000010001101101",
			279 => "11111111111010010000010001101101",
			280 => "0000001111000000000111011000000100",
			281 => "00000000101110110000010001101101",
			282 => "00000000000000000000010001101101",
			283 => "0000000010000000000111011000000100",
			284 => "11111110100011100000010010111001",
			285 => "0000000110000000001011001100001100",
			286 => "0000000001000000000110101000000100",
			287 => "00000000000000000000010010111001",
			288 => "0000001111000000001110110100000100",
			289 => "00000001001100000000010010111001",
			290 => "00000000000000000000010010111001",
			291 => "0000000001000000001101011100001100",
			292 => "0000000111000000000011100000001000",
			293 => "0000001010000000000001010000000100",
			294 => "00000000000000000000010010111001",
			295 => "11111110111111000000010010111001",
			296 => "00000000000000000000010010111001",
			297 => "0000001110000000001110101000001000",
			298 => "0000001010000000000001010000000100",
			299 => "00000000000000000000010010111001",
			300 => "00000000111111000000010010111001",
			301 => "11111111011101100000010010111001",
			302 => "0000000100000000000010100100001000",
			303 => "0000000100000000000011110100000100",
			304 => "11111110100101010000010100000101",
			305 => "00000000000000000000010100000101",
			306 => "0000000001000000000110101000000100",
			307 => "11111111000011110000010100000101",
			308 => "0000000101000000000101100100001100",
			309 => "0000000110000000001111000000001000",
			310 => "0000001010000000001100000100000100",
			311 => "00000001010110010000010100000101",
			312 => "00000000000000000000010100000101",
			313 => "00000000000000000000010100000101",
			314 => "0000000001000000001101011100000100",
			315 => "11111111000111100000010100000101",
			316 => "0000001111000000000111011000001000",
			317 => "0000000010000000001011111000000100",
			318 => "00000000000000000000010100000101",
			319 => "00000001000100000000010100000101",
			320 => "00000000000000000000010100000101",
			321 => "0000000010000000000000010000010100",
			322 => "0000000001000000001111001100000100",
			323 => "11111110011110000000010101101001",
			324 => "0000000101000000001011011100001100",
			325 => "0000000010000000000000010000001000",
			326 => "0000001110000000001110101100000100",
			327 => "00000000111010110000010101101001",
			328 => "00000000000000000000010101101001",
			329 => "00000000000000000000010101101001",
			330 => "11111110100111000000010101101001",
			331 => "0000000110000000001011001100001100",
			332 => "0000000001000000000110101000000100",
			333 => "00000000000000000000010101101001",
			334 => "0000000011000000000011001000000100",
			335 => "00000010001010100000010101101001",
			336 => "00000000000000000000010101101001",
			337 => "0000001111000000001100000000010000",
			338 => "0000001001000000001010011000000100",
			339 => "11111111001110000000010101101001",
			340 => "0000000010000000001011111000001000",
			341 => "0000000011000000001101000100000100",
			342 => "00000000000000000000010101101001",
			343 => "11111111110101000000010101101001",
			344 => "00000001010001110000010101101001",
			345 => "11111110110100000000010101101001",
			346 => "0000000010000000000000010000001100",
			347 => "0000001100000000001110001100001000",
			348 => "0000000111000000000001111100000100",
			349 => "11111110111100100000010110110101",
			350 => "00000000000000000000010110110101",
			351 => "00000000000000000000010110110101",
			352 => "0000001100000000000100001000011000",
			353 => "0000001100000000001100110000000100",
			354 => "00000000000000000000010110110101",
			355 => "0000000010000000001101101100010000",
			356 => "0000000010000000001011111000000100",
			357 => "00000000000000000000010110110101",
			358 => "0000000100000000000011110100000100",
			359 => "00000000000000000000010110110101",
			360 => "0000000000000000001100101100000100",
			361 => "00000000111010110000010110110101",
			362 => "00000000000000000000010110110101",
			363 => "00000000000000000000010110110101",
			364 => "00000000000000000000010110110101",
			365 => "0000000010000000000111011000000100",
			366 => "11111110100010100000010111111001",
			367 => "0000001111000000001100000000011100",
			368 => "0000000010000000000110101100010000",
			369 => "0000001010000000000001010000001100",
			370 => "0000001110000000001110101100001000",
			371 => "0000000001000000001111001100000100",
			372 => "00000000000000000000010111111001",
			373 => "00000000111111010000010111111001",
			374 => "00000000000000000000010111111001",
			375 => "11111111001100010000010111111001",
			376 => "0000001010000000001100000100001000",
			377 => "0000001100000000000011011100000100",
			378 => "00000000000000000000010111111001",
			379 => "00000001000010110000010111111001",
			380 => "00000000000000000000010111111001",
			381 => "11111110111111000000010111111001",
			382 => "0000000010000000000000010000011000",
			383 => "0000000001000000001111001100000100",
			384 => "11111110011110100000011001011101",
			385 => "0000001011000000000011100000001100",
			386 => "0000000010000000000000010000001000",
			387 => "0000001110000000001110101000000100",
			388 => "00000000110100110000011001011101",
			389 => "00000000000000000000011001011101",
			390 => "00000000000000000000011001011101",
			391 => "0000001110000000000111110000000100",
			392 => "00000000000000000000011001011101",
			393 => "11111110101011000000011001011101",
			394 => "0000001111000000001100000000011000",
			395 => "0000000110000000001011001100001000",
			396 => "0000000001000000000110101000000100",
			397 => "00000000000000000000011001011101",
			398 => "00000001111110110000011001011101",
			399 => "0000001001000000001010011000000100",
			400 => "11111111010010110000011001011101",
			401 => "0000000010000000001011111000001000",
			402 => "0000001101000000000101110100000100",
			403 => "00000000000000000000011001011101",
			404 => "11111111111010100000011001011101",
			405 => "00000001001111000000011001011101",
			406 => "11111110110110010000011001011101",
			407 => "0000000100000000000000010100000100",
			408 => "11111111111000010000011010011001",
			409 => "0000000001000000000110101000000100",
			410 => "00000000000000000000011010011001",
			411 => "0000000010000000001101101100010100",
			412 => "0000000110000000001111000000010000",
			413 => "0000001100000000000100001000001100",
			414 => "0000000111000000000110000100000100",
			415 => "00000000000000000000011010011001",
			416 => "0000001100000000001100110000000100",
			417 => "00000000000000000000011010011001",
			418 => "00000000011001100000011010011001",
			419 => "00000000000000000000011010011001",
			420 => "00000000000000000000011010011001",
			421 => "00000000000000000000011010011001",
			422 => "0000000001000000000110101000000100",
			423 => "11111111000110010000011011101101",
			424 => "0000000110000000001011001100001100",
			425 => "0000000100000000001110111000000100",
			426 => "00000000000000000000011011101101",
			427 => "0000000110000000001011001100000100",
			428 => "00000000100100000000011011101101",
			429 => "00000000000000000000011011101101",
			430 => "0000001000000000000110001000010100",
			431 => "0000001100000000000100001000010000",
			432 => "0000000110000000001011001100000100",
			433 => "00000000000000000000011011101101",
			434 => "0000000110000000001001100100001000",
			435 => "0000000000000000000010011000000100",
			436 => "00000000000000000000011011101101",
			437 => "00000000001110100000011011101101",
			438 => "00000000000000000000011011101101",
			439 => "00000000000000000000011011101101",
			440 => "0000000001000000001101011100000100",
			441 => "11111111100000110000011011101101",
			442 => "00000000000000000000011011101101",
			443 => "0000000001000000001101101000000100",
			444 => "11111110011011010000011101001001",
			445 => "0000001100000000000100001000100100",
			446 => "0000001110000000001001010100010100",
			447 => "0000001101000000000010001000001100",
			448 => "0000001111000000001001010000000100",
			449 => "00000000000000000000011101001001",
			450 => "0000001011000000000001111100000100",
			451 => "00000000000000000000011101001001",
			452 => "00000001110101000000011101001001",
			453 => "0000001001000000001010011000000100",
			454 => "11111110110011000000011101001001",
			455 => "00000001011010010000011101001001",
			456 => "0000001100000000001110001100001000",
			457 => "0000001010000000000110011000000100",
			458 => "00000000000000000000011101001001",
			459 => "11111110010011000000011101001001",
			460 => "0000001110000000001110101000000100",
			461 => "00000001010000100000011101001001",
			462 => "00000000000000000000011101001001",
			463 => "0000001110000000000111110000000100",
			464 => "00000000000000000000011101001001",
			465 => "11111110100001000000011101001001",
			466 => "0000001001000000001110010100000100",
			467 => "11111110011011100000011110100101",
			468 => "0000000011000000000110100000010100",
			469 => "0000000100000000000000010100000100",
			470 => "11111111110000110000011110100101",
			471 => "0000001000000000001000101100001100",
			472 => "0000001100000000001100110000000100",
			473 => "00000000000000000000011110100101",
			474 => "0000000010000000001111100100000100",
			475 => "00000000111110110000011110100101",
			476 => "00000001111110100000011110100101",
			477 => "00000000000000000000011110100101",
			478 => "0000001101000000000000110100010100",
			479 => "0000000010000000001011111000001100",
			480 => "0000001010000000000110011000001000",
			481 => "0000000100000000001110111000000100",
			482 => "00000000000000000000011110100101",
			483 => "00000000100101000000011110100101",
			484 => "11111110010100010000011110100101",
			485 => "0000001111000000000111011000000100",
			486 => "00000001011011010000011110100101",
			487 => "00000000000000000000011110100101",
			488 => "11111110100000000000011110100101",
			489 => "0000000100000000000010100100001000",
			490 => "0000000100000000000011110100000100",
			491 => "11111110100011010000100000011001",
			492 => "00000000000000000000100000011001",
			493 => "0000000010000000000110101100010100",
			494 => "0000001000000000001011010100001100",
			495 => "0000001111000000001100010100001000",
			496 => "0000000001000000001111001100000100",
			497 => "00000000000000000000100000011001",
			498 => "00000000101110010000100000011001",
			499 => "00000000000000000000100000011001",
			500 => "0000001010000000000110011000000100",
			501 => "00000000000000000000100000011001",
			502 => "11111110111000000000100000011001",
			503 => "0000000011000000000010110100010100",
			504 => "0000001010000000001100000100010000",
			505 => "0000000010000000000110101100000100",
			506 => "00000000000000000000100000011001",
			507 => "0000000010000000001101101100001000",
			508 => "0000000111000000000110000100000100",
			509 => "00000000000000000000100000011001",
			510 => "00000001110110000000100000011001",
			511 => "00000000000000000000100000011001",
			512 => "00000000000000000000100000011001",
			513 => "0000000001000000001101011100000100",
			514 => "11111111001001100000100000011001",
			515 => "0000001101000000001110101100000100",
			516 => "00000000101110110000100000011001",
			517 => "00000000000000000000100000011001",
			518 => "0000000001000000001101101000000100",
			519 => "11111110011010010000100001100101",
			520 => "0000001101000000000000110100100000",
			521 => "0000000100000000001110111000000100",
			522 => "11111110111010110000100001100101",
			523 => "0000000101000000000101100100001100",
			524 => "0000001100000000001100110000000100",
			525 => "00000000001010100000100001100101",
			526 => "0000000000000000001100001000000100",
			527 => "00000001100100000000100001100101",
			528 => "00000010101100100000100001100101",
			529 => "0000001001000000001010011000000100",
			530 => "11111110011011110000100001100101",
			531 => "0000001100000000000110000100000100",
			532 => "00000000000000000000100001100101",
			533 => "0000000001000000001101011100000100",
			534 => "00000000000000000000100001100101",
			535 => "00000001011110110000100001100101",
			536 => "11111110011010000000100001100101",
			537 => "0000000001000000001101101000000100",
			538 => "11111110011010110000100011000001",
			539 => "0000001101000000000000110100101000",
			540 => "0000000010000000001011111000011100",
			541 => "0000001110000000001001010100001100",
			542 => "0000001010000000001010110000001000",
			543 => "0000000010000000000111011000000100",
			544 => "00000000000000000000100011000001",
			545 => "00000001011110100000100011000001",
			546 => "11111111000011010000100011000001",
			547 => "0000001100000000001110001100001000",
			548 => "0000001010000000000110011000000100",
			549 => "00000000000000000000100011000001",
			550 => "11111110000010110000100011000001",
			551 => "0000000011000000000111100000000100",
			552 => "00000000001001100000100011000001",
			553 => "00000000000000000000100011000001",
			554 => "0000000110000000000100111100001000",
			555 => "0000001010000000000001010100000100",
			556 => "00000001101100000000100011000001",
			557 => "00000000000000000000100011000001",
			558 => "00000000000000000000100011000001",
			559 => "11111110011100100000100011000001",
			560 => "0000000010000000001111010100001000",
			561 => "0000000010000000000111011000000100",
			562 => "11111110011100110000100100110101",
			563 => "00000000000000000000100100110101",
			564 => "0000001110000000001010111000010000",
			565 => "0000000001000000000110101000000100",
			566 => "00000000000000000000100100110101",
			567 => "0000001011000000000000001100000100",
			568 => "00000110001010000000100100110101",
			569 => "0000000001000000000111100100000100",
			570 => "00000000000000000000100100110101",
			571 => "00000010000001010000100100110101",
			572 => "0000001110000000001110101000100000",
			573 => "0000001000000000001011010100001100",
			574 => "0000000111000000001101010100000100",
			575 => "00000001011000000000100100110101",
			576 => "0000000111000000000111001000000100",
			577 => "00000000000000000000100100110101",
			578 => "00000000011110010000100100110101",
			579 => "0000000010000000000110101100001100",
			580 => "0000001011000000001010111000001000",
			581 => "0000000001000000001101101000000100",
			582 => "00000000000000000000100100110101",
			583 => "00000000001110100000100100110101",
			584 => "11111110101111010000100100110101",
			585 => "0000001000000000000001110100000100",
			586 => "00000001001100000000100100110101",
			587 => "11111111011010100000100100110101",
			588 => "11111110101010000000100100110101",
			589 => "0000000010000000000111011000000100",
			590 => "11111110100101110000100110010001",
			591 => "0000001111000000001100000000101000",
			592 => "0000001000000000001011010100001100",
			593 => "0000000100000000001110111000000100",
			594 => "00000000000000000000100110010001",
			595 => "0000000001000000001111001100000100",
			596 => "00000000000000000000100110010001",
			597 => "00000001000110010000100110010001",
			598 => "0000000110000000001101011000001000",
			599 => "0000000001000000000110101000000100",
			600 => "00000000000000000000100110010001",
			601 => "00000000111001000000100110010001",
			602 => "0000000010000000001000100000001000",
			603 => "0000000110000000001011001100000100",
			604 => "00000000000000000000100110010001",
			605 => "11111111001111000000100110010001",
			606 => "0000001001000000001010011000001000",
			607 => "0000000110000000001011001100000100",
			608 => "00000000000000000000100110010001",
			609 => "11111111110100100000100110010001",
			610 => "00000000101010000000100110010001",
			611 => "11111111001001000000100110010001",
			612 => "0000000010000000001111010100001000",
			613 => "0000000010000000000111011000000100",
			614 => "11111110011000100000101000010101",
			615 => "11111110110011100000101000010101",
			616 => "0000001100000000000100001000101000",
			617 => "0000000001000000001101101000001100",
			618 => "0000001100000000000110000100000100",
			619 => "11111110011101000000101000010101",
			620 => "0000000000000000001100101100000100",
			621 => "00000110001101110000101000010101",
			622 => "11111110101100110000101000010101",
			623 => "0000000011000000000001011000000100",
			624 => "00010101011000010000101000010101",
			625 => "0000000011000000000111110000001000",
			626 => "0000001010000000000101000100000100",
			627 => "00000101000111110000101000010101",
			628 => "11111111111101010000101000010101",
			629 => "0000001001000000001010011000001000",
			630 => "0000001010000000000001010000000100",
			631 => "00000000010011110000101000010101",
			632 => "11111101001000010000101000010101",
			633 => "0000000011000000001001011100000100",
			634 => "00000001101111000000101000010101",
			635 => "11111110101000010000101000010101",
			636 => "0000000111000000000111001000001100",
			637 => "0000000101000000000101100100000100",
			638 => "11111111000011000000101000010101",
			639 => "0000001100000000000100001000000100",
			640 => "11111111011111110000101000010101",
			641 => "00000001010011110000101000010101",
			642 => "0000001100000000000100001000000100",
			643 => "00000000000000000000101000010101",
			644 => "11111110011001010000101000010101",
			645 => "0000000010000000001111010100001100",
			646 => "0000000010000000000111011000000100",
			647 => "11111110011010000000101010000001",
			648 => "0000000010000000000110111100000100",
			649 => "00000000000000000000101010000001",
			650 => "11111111000100000000101010000001",
			651 => "0000001111000000001100000000101000",
			652 => "0000001001000000001110010100000100",
			653 => "11111110100100010000101010000001",
			654 => "0000000101000000000101100100001100",
			655 => "0000001100000000000011011100000100",
			656 => "00000000000000000000101010000001",
			657 => "0000001010000000000001010100000100",
			658 => "00000001101111010000101010000001",
			659 => "00000000000000000000101010000001",
			660 => "0000000010000000000110101100001100",
			661 => "0000001000000000001011010100001000",
			662 => "0000000011000000000111100000000100",
			663 => "00000001010110100000101010000001",
			664 => "11111111001001110000101010000001",
			665 => "11111110000101000000101010000001",
			666 => "0000001001000000001010011000000100",
			667 => "11111111011011100000101010000001",
			668 => "0000000111000000000100001000000100",
			669 => "00000000000000000000101010000001",
			670 => "00000001101011000000101010000001",
			671 => "11111110011001000000101010000001",
			672 => "0000000001000000001101101000000100",
			673 => "11111110011010000000101011011101",
			674 => "0000001101000000000000110100101000",
			675 => "0000000100000000001110111000000100",
			676 => "11111110110110100000101011011101",
			677 => "0000000101000000000101100100001100",
			678 => "0000000000000000000100000000001000",
			679 => "0000001010000000000110011100000100",
			680 => "00000001100101110000101011011101",
			681 => "00000000000000000000101011011101",
			682 => "00000011011011000000101011011101",
			683 => "0000000001000000001101011100001100",
			684 => "0000001010000000001010110000000100",
			685 => "00000000110100100000101011011101",
			686 => "0000001111000000000010000000000100",
			687 => "11111110010001100000101011011101",
			688 => "00000000000000000000101011011101",
			689 => "0000001100000000001110001100001000",
			690 => "0000000010000000001011111000000100",
			691 => "00000000000000000000101011011101",
			692 => "00000000110111100000101011011101",
			693 => "00000001101010000000101011011101",
			694 => "11111110011001100000101011011101",
			695 => "0000000010000000001111010100000100",
			696 => "11111110011001110000101101011011",
			697 => "0000001100000000000100001000101100",
			698 => "0000000001000000001101101000000100",
			699 => "11111110011110110000101101011011",
			700 => "0000001110000000001001010100010000",
			701 => "0000001000000000001000101100001100",
			702 => "0000000001000000001111001100000100",
			703 => "00000011010011010000101101011011",
			704 => "0000000001000000001101011100000100",
			705 => "00000000001001010000101101011011",
			706 => "00000001101011100000101101011011",
			707 => "11111110101001010000101101011011",
			708 => "0000000001000000001001011000001100",
			709 => "0000000100000000001101110100001000",
			710 => "0000000100000000000000010100000100",
			711 => "11111110111100010000101101011011",
			712 => "00000000000000000000101101011011",
			713 => "11111011111100010000101101011011",
			714 => "0000001110000000001110101000001000",
			715 => "0000000010000000000110101100000100",
			716 => "00000000100111110000101101011011",
			717 => "00000011011000010000101101011011",
			718 => "11111110101111110000101101011011",
			719 => "0000000111000000000111001000001100",
			720 => "0000001110000000000111110000001000",
			721 => "0000001110000000001000110000000100",
			722 => "11111111100100110000101101011011",
			723 => "00000000111100000000101101011011",
			724 => "11111110011110100000101101011011",
			725 => "11111110011001100000101101011011",
			726 => "00000000000000000000101101011101",
			727 => "00000000000000000000101101100001",
			728 => "00000000000000000000101101100101",
			729 => "00000000000000000000101101101001",
			730 => "00000000000000000000101101101101",
			731 => "00000000000000000000101101110001",
			732 => "00000000000000000000101101110101",
			733 => "00000000000000000000101101111001",
			734 => "00000000000000000000101101111101",
			735 => "00000000000000000000101110000001",
			736 => "00000000000000000000101110000101",
			737 => "00000000000000000000101110001001",
			738 => "00000000000000000000101110001101",
			739 => "00000000000000000000101110010001",
			740 => "00000000000000000000101110010101",
			741 => "00000000000000000000101110011001",
			742 => "00000000000000000000101110011101",
			743 => "00000000000000000000101110100001",
			744 => "00000000000000000000101110100101",
			745 => "00000000000000000000101110101001",
			746 => "00000000000000000000101110101101",
			747 => "00000000000000000000101110110001",
			748 => "00000000000000000000101110110101",
			749 => "00000000000000000000101110111001",
			750 => "00000000000000000000101110111101",
			751 => "00000000000000000000101111000001",
			752 => "00000000000000000000101111000101",
			753 => "00000000000000000000101111001001",
			754 => "00000000000000000000101111001101",
			755 => "0000000100000000000100111000000100",
			756 => "11111111111110110000101111011001",
			757 => "00000000000000000000101111011001",
			758 => "0000000100000000000011011000000100",
			759 => "11111111111110010000101111100101",
			760 => "00000000000000000000101111100101",
			761 => "0000000010000000000110101100000100",
			762 => "11111111111010010000101111110001",
			763 => "00000000000000000000101111110001",
			764 => "0000000100000000000011111000000100",
			765 => "11111111111011100000101111111101",
			766 => "00000000000000000000101111111101",
			767 => "0000000001000000001111001100000100",
			768 => "11111111111001110000110000001001",
			769 => "00000000000000000000110000001001",
			770 => "0000000010000000001011101100000100",
			771 => "11111111111111010000110000010101",
			772 => "00000000000000000000110000010101",
			773 => "0000000100000000000011111000000100",
			774 => "11111111111110110000110000100001",
			775 => "00000000000000000000110000100001",
			776 => "0000000100000000000000010100000100",
			777 => "11111111111100100000110000110101",
			778 => "0000000100000000001010010000000100",
			779 => "00000000000001100000110000110101",
			780 => "00000000000000000000110000110101",
			781 => "0000000100000000000011010100000100",
			782 => "00000000000000000000110001001001",
			783 => "0000000100000000001010010000000100",
			784 => "00000000000010110000110001001001",
			785 => "00000000000000000000110001001001",
			786 => "0000000100000000000010100100000100",
			787 => "00000000000000000000110001011101",
			788 => "0000000100000000001010010000000100",
			789 => "00000000000011110000110001011101",
			790 => "00000000000000000000110001011101",
			791 => "0000000010000000001011111000000100",
			792 => "11111111111111110000110001110001",
			793 => "0000000010000000001101101100000100",
			794 => "00000000001100000000110001110001",
			795 => "00000000000000000000110001110001",
			796 => "0000000010000000000110101100000100",
			797 => "11111111111101010000110010000101",
			798 => "0000000010000000001111101000000100",
			799 => "00000000001010010000110010000101",
			800 => "00000000000000000000110010000101",
			801 => "0000000100000000000011011000001000",
			802 => "0000001010000000000110011000000100",
			803 => "00000000000000000000110010011001",
			804 => "11111111110111110000110010011001",
			805 => "00000000000000000000110010011001",
			806 => "0000000001000000001111001100000100",
			807 => "11111111100101100000110010110101",
			808 => "0000001110000000001001010100001000",
			809 => "0000000111000000001101111000000100",
			810 => "00000000000000000000110010110101",
			811 => "00000000100000000000110010110101",
			812 => "00000000000000000000110010110101",
			813 => "0000000100000000000101100000001100",
			814 => "0000000001000000001101011100001000",
			815 => "0000001001000000001101011000000100",
			816 => "11111111100100010000110011010001",
			817 => "00000000000000000000110011010001",
			818 => "00000000000000000000110011010001",
			819 => "00000000000000000000110011010001",
			820 => "0000000100000000000011010100000100",
			821 => "11111111111100100000110011101101",
			822 => "0000000010000000000000010000000100",
			823 => "00000000000000000000110011101101",
			824 => "0000000010000000001111101000000100",
			825 => "00000000000110010000110011101101",
			826 => "00000000000000000000110011101101",
			827 => "0000001001000000001101011000001100",
			828 => "0000000100000000000100111000001000",
			829 => "0000000001000000001101011100000100",
			830 => "11111111101100100000110100001001",
			831 => "00000000000000000000110100001001",
			832 => "00000000000000000000110100001001",
			833 => "00000000000000000000110100001001",
			834 => "0000000001000000001101011100001100",
			835 => "0000000010000000001011101100001000",
			836 => "0000001001000000001101011000000100",
			837 => "11111111110101000000110100100101",
			838 => "00000000000000000000110100100101",
			839 => "00000000000000000000110100100101",
			840 => "00000000000000000000110100100101",
			841 => "0000000001000000001111001100000100",
			842 => "11111111010011010000110101001001",
			843 => "0000001101000000001001010100001100",
			844 => "0000001100000000000000001100001000",
			845 => "0000001110000000001110101000000100",
			846 => "00000000100110010000110101001001",
			847 => "00000000000000000000110101001001",
			848 => "00000000000000000000110101001001",
			849 => "00000000000000000000110101001001",
			850 => "0000000100000000000000010100000100",
			851 => "11111111111000100000110101101101",
			852 => "0000001001000000001011111100000100",
			853 => "00000000000000000000110101101101",
			854 => "0000000010000000001111101000001000",
			855 => "0000000111000000001110001100000100",
			856 => "00000000000000000000110101101101",
			857 => "00000000001000110000110101101101",
			858 => "00000000000000000000110101101101",
			859 => "0000000100000000000011010100000100",
			860 => "11111111111101100000110110010001",
			861 => "0000000010000000000110101100000100",
			862 => "00000000000000000000110110010001",
			863 => "0000000010000000000011000000001000",
			864 => "0000000100000000001010010000000100",
			865 => "00000000001111010000110110010001",
			866 => "00000000000000000000110110010001",
			867 => "00000000000000000000110110010001",
			868 => "0000000100000000000011011000000100",
			869 => "11111111111001010000110110110101",
			870 => "0000001101000000000100010000001100",
			871 => "0000001101000000001000011000000100",
			872 => "00000000000000000000110110110101",
			873 => "0000001011000000001000000000000100",
			874 => "00000000000111010000110110110101",
			875 => "00000000000000000000110110110101",
			876 => "00000000000000000000110110110101",
			877 => "0000000001000000001111001100001000",
			878 => "0000000100000000000100111000000100",
			879 => "11111111100001000000110111100001",
			880 => "00000000000000000000110111100001",
			881 => "0000001110000000000111110000001100",
			882 => "0000000111000000001101111000000100",
			883 => "00000000000000000000110111100001",
			884 => "0000000110000000001001100100000100",
			885 => "00000000010111010000110111100001",
			886 => "00000000000000000000110111100001",
			887 => "00000000000000000000110111100001",
			888 => "0000000001000000001101011100001000",
			889 => "0000000010000000001011101100000100",
			890 => "11111111101010100000111000001101",
			891 => "00000000000000000000111000001101",
			892 => "0000001011000000000001101000001100",
			893 => "0000000111000000001100101000000100",
			894 => "00000000000000000000111000001101",
			895 => "0000000100000000001110111000000100",
			896 => "00000000000000000000111000001101",
			897 => "00000000010000000000111000001101",
			898 => "00000000000000000000111000001101",
			899 => "0000000010000000000110101100001100",
			900 => "0000000000000000000011111100000100",
			901 => "00000000000000000000111001000001",
			902 => "0000000110000000001001100100000100",
			903 => "11111111011111000000111001000001",
			904 => "00000000000000000000111001000001",
			905 => "0000001111000000001100010000001100",
			906 => "0000000001000000001111001100000100",
			907 => "00000000000000000000111001000001",
			908 => "0000000010000000000001011100000100",
			909 => "00000000100111010000111001000001",
			910 => "00000000000000000000111001000001",
			911 => "00000000000000000000111001000001",
			912 => "0000000100000000000011110100000100",
			913 => "11111111011001110000111001110101",
			914 => "0000001011000000000011100000001100",
			915 => "0000000001000000001111001100000100",
			916 => "00000000000000000000111001110101",
			917 => "0000000111000000001101111000000100",
			918 => "00000000000000000000111001110101",
			919 => "00000000100110010000111001110101",
			920 => "0000001000000000001011010100000100",
			921 => "00000000000000000000111001110101",
			922 => "0000001101000000000101110100000100",
			923 => "00000000000000000000111001110101",
			924 => "11111111101010010000111001110101",
			925 => "0000001001000000000100110100000100",
			926 => "11111111011011000000111010100001",
			927 => "0000001101000000001001010100010000",
			928 => "0000001100000000000000001100001100",
			929 => "0000000111000000001110001100000100",
			930 => "00000000000000000000111010100001",
			931 => "0000001110000000001110101000000100",
			932 => "00000000011100010000111010100001",
			933 => "00000000000000000000111010100001",
			934 => "00000000000000000000111010100001",
			935 => "00000000000000000000111010100001",
			936 => "0000000100000000000000010100000100",
			937 => "11111111111010010000111011001101",
			938 => "0000001100000000001100110000000100",
			939 => "00000000000000000000111011001101",
			940 => "0000000010000000001101101100001100",
			941 => "0000000100000000001010010000001000",
			942 => "0000001100000000000100001000000100",
			943 => "00000000010001100000111011001101",
			944 => "00000000000000000000111011001101",
			945 => "00000000000000000000111011001101",
			946 => "00000000000000000000111011001101",
			947 => "0000000111000000000110000100001000",
			948 => "0000000001000000001111001100000100",
			949 => "11111110110111110000111100010001",
			950 => "00000000000000000000111100010001",
			951 => "0000000011000000001101000100010000",
			952 => "0000000001000000001111001100000100",
			953 => "00000000000000000000111100010001",
			954 => "0000000111000000001101111000000100",
			955 => "00000000000000000000111100010001",
			956 => "0000001100000000000000001100000100",
			957 => "00000001000001100000111100010001",
			958 => "00000000000000000000111100010001",
			959 => "0000000101000000000101100100000100",
			960 => "00000000000000000000111100010001",
			961 => "0000001010000000000001010000000100",
			962 => "11111111001111000000111100010001",
			963 => "00000000000000000000111100010001",
			964 => "0000000100000000000011111000011000",
			965 => "0000001001000000001100011000000100",
			966 => "11111110011111110000111101011101",
			967 => "0000001110000000000111110000001000",
			968 => "0000001001000000001010011000000100",
			969 => "00000000000000000000111101011101",
			970 => "00000001001101110000111101011101",
			971 => "0000001011000000000011100000000100",
			972 => "00000000000000000000111101011101",
			973 => "0000001100000000000110000100000100",
			974 => "00000000000000000000111101011101",
			975 => "11111110111000000000111101011101",
			976 => "0000001010000000001100000100001100",
			977 => "0000001101000000000001011000001000",
			978 => "0000000010000000001111100100000100",
			979 => "00000000000000000000111101011101",
			980 => "00000010001101100000111101011101",
			981 => "00000000000000000000111101011101",
			982 => "11111111010000100000111101011101",
			983 => "0000000100000000000000010100000100",
			984 => "11111111010010000000111110011001",
			985 => "0000000010000000000110101100001000",
			986 => "0000001000000000001011010100000100",
			987 => "00000000001000110000111110011001",
			988 => "11111111100101110000111110011001",
			989 => "0000000110000000000100111100010000",
			990 => "0000001100000000000011011100000100",
			991 => "00000000000000000000111110011001",
			992 => "0000001010000000001100000100001000",
			993 => "0000001100000000000100001000000100",
			994 => "00000000101111000000111110011001",
			995 => "00000000000000000000111110011001",
			996 => "00000000000000000000111110011001",
			997 => "00000000000000000000111110011001",
			998 => "0000000010000000001000001100001100",
			999 => "0000001100000000001110001100001000",
			1000 => "0000000111000000001100101000000100",
			1001 => "11111110101000010000111111100101",
			1002 => "00000000000000000000111111100101",
			1003 => "00000000000000000000111111100101",
			1004 => "0000001111000000001100000000011000",
			1005 => "0000000001000000001111001100010000",
			1006 => "0000001111000000001110000100001100",
			1007 => "0000000000000000001100101100001000",
			1008 => "0000000000000000001001110000000100",
			1009 => "00000000000000000000111111100101",
			1010 => "00000000011001000000111111100101",
			1011 => "00000000000000000000111111100101",
			1012 => "11111111101110100000111111100101",
			1013 => "0000000010000000001011111000000100",
			1014 => "00000000000000000000111111100101",
			1015 => "00000000111110100000111111100101",
			1016 => "11111111011001110000111111100101",
			1017 => "0000000001000000001111001100100000",
			1018 => "0000000001000000001111001100011000",
			1019 => "0000000010000000001011111000000100",
			1020 => "10111101000111000001000000111001",
			1021 => "0000000010000000000110101100001000",
			1022 => "0000000001000000000110000000000100",
			1023 => "10111110000000110001000000111001",
			1024 => "11001011100010010001000000111001",
			1025 => "0000000110000000001011001100001000",
			1026 => "0000000001000000000110101000000100",
			1027 => "10111101001100000001000000111001",
			1028 => "11001011100010010001000000111001",
			1029 => "10111101000111100001000000111001",
			1030 => "0000001110000000000100010000000100",
			1031 => "11100101111110010001000000111001",
			1032 => "10111101001001000001000000111001",
			1033 => "0000001110000000001110101100000100",
			1034 => "00011001100100010001000000111001",
			1035 => "0000001110000000001110101000000100",
			1036 => "11011000001111010001000000111001",
			1037 => "10111101000111000001000000111001",
			1038 => "0000000100000000000010100100001000",
			1039 => "0000000100000000000011110100000100",
			1040 => "11111110100110110001000010000101",
			1041 => "00000000000000000001000010000101",
			1042 => "0000000001000000000110101000000100",
			1043 => "11111111000111100001000010000101",
			1044 => "0000001101000000000101110100001100",
			1045 => "0000000110000000001111000000001000",
			1046 => "0000001010000000001100000100000100",
			1047 => "00000001000111010001000010000101",
			1048 => "00000000000000000001000010000101",
			1049 => "00000000000000000001000010000101",
			1050 => "0000000001000000001101011100000100",
			1051 => "11111111001011110001000010000101",
			1052 => "0000000110000000000100111100001000",
			1053 => "0000000010000000001011111000000100",
			1054 => "00000000000000000001000010000101",
			1055 => "00000000111000110001000010000101",
			1056 => "00000000000000000001000010000101",
			1057 => "0000000010000000000000010000001100",
			1058 => "0000001001000000001111000000001000",
			1059 => "0000001100000000001110001100000100",
			1060 => "11111110100111000001000011011001",
			1061 => "00000000000000000001000011011001",
			1062 => "00000000000000000001000011011001",
			1063 => "0000001111000000000010000100011000",
			1064 => "0000000010000000000110101100000100",
			1065 => "00000000000000000001000011011001",
			1066 => "0000001100000000001100110000000100",
			1067 => "00000000000000000001000011011001",
			1068 => "0000001010000000001100000100001100",
			1069 => "0000000010000000000001011100001000",
			1070 => "0000000110000000001111000000000100",
			1071 => "00000001001001110001000011011001",
			1072 => "00000000000000000001000011011001",
			1073 => "00000000000000000001000011011001",
			1074 => "00000000000000000001000011011001",
			1075 => "0000001111000000001100000000000100",
			1076 => "00000000000000000001000011011001",
			1077 => "11111111010011000001000011011001",
			1078 => "0000000010000000001000001100001100",
			1079 => "0000000111000000001100101000001000",
			1080 => "0000001100000000001110001100000100",
			1081 => "11111110111011010001000100100101",
			1082 => "00000000000000000001000100100101",
			1083 => "00000000000000000001000100100101",
			1084 => "0000001100000000000100001000011000",
			1085 => "0000001100000000001100110000000100",
			1086 => "00000000000000000001000100100101",
			1087 => "0000000010000000001011111000000100",
			1088 => "00000000000000000001000100100101",
			1089 => "0000000010000000001101101100001100",
			1090 => "0000000100000000000011110100000100",
			1091 => "00000000000000000001000100100101",
			1092 => "0000000000000000001100101100000100",
			1093 => "00000000110110110001000100100101",
			1094 => "00000000000000000001000100100101",
			1095 => "00000000000000000001000100100101",
			1096 => "00000000000000000001000100100101",
			1097 => "0000000010000000001000001100001000",
			1098 => "0000001100000000001110001100000100",
			1099 => "11111111000001100001000101101001",
			1100 => "00000000000000000001000101101001",
			1101 => "0000001100000000000100001000011000",
			1102 => "0000001100000000001100110000000100",
			1103 => "00000000000000000001000101101001",
			1104 => "0000000010000000001011111000000100",
			1105 => "00000000000000000001000101101001",
			1106 => "0000000010000000001101101100001100",
			1107 => "0000000100000000000011110100000100",
			1108 => "00000000000000000001000101101001",
			1109 => "0000000000000000001100101100000100",
			1110 => "00000000110010110001000101101001",
			1111 => "00000000000000000001000101101001",
			1112 => "00000000000000000001000101101001",
			1113 => "00000000000000000001000101101001",
			1114 => "0000000111000000000110000100000100",
			1115 => "11111111000100010001000110111101",
			1116 => "0000000011000000001101000100010100",
			1117 => "0000001010000000000101000100010000",
			1118 => "0000001001000000001110010100000100",
			1119 => "00000000000000000001000110111101",
			1120 => "0000001100000000001100110000000100",
			1121 => "00000000000000000001000110111101",
			1122 => "0000000100000000000000010100000100",
			1123 => "00000000000000000001000110111101",
			1124 => "00000000101010110001000110111101",
			1125 => "00000000000000000001000110111101",
			1126 => "0000000110000000001001100100001000",
			1127 => "0000001011000000000011100000000100",
			1128 => "00000000000000000001000110111101",
			1129 => "11111111101000000001000110111101",
			1130 => "0000000110000000001001100100001000",
			1131 => "0000001011000000000110100100000100",
			1132 => "00000000001101100001000110111101",
			1133 => "00000000000000000001000110111101",
			1134 => "00000000000000000001000110111101",
			1135 => "0000000100000000000000010100000100",
			1136 => "11111111111001100001000111111001",
			1137 => "0000000001000000000110101000000100",
			1138 => "00000000000000000001000111111001",
			1139 => "0000000010000000001101101100010100",
			1140 => "0000000110000000001111000000010000",
			1141 => "0000001100000000000100001000001100",
			1142 => "0000000111000000000110000100000100",
			1143 => "00000000000000000001000111111001",
			1144 => "0000001100000000001100110000000100",
			1145 => "00000000000000000001000111111001",
			1146 => "00000000010110100001000111111001",
			1147 => "00000000000000000001000111111001",
			1148 => "00000000000000000001000111111001",
			1149 => "00000000000000000001000111111001",
			1150 => "0000000111000000000110000100001000",
			1151 => "0000000001000000001111001100000100",
			1152 => "11111110100100100001001001011101",
			1153 => "00000000000000000001001001011101",
			1154 => "0000001100000000000100001000100100",
			1155 => "0000000001000000001101011100011000",
			1156 => "0000000110000000001011001100001100",
			1157 => "0000001111000000001110101000000100",
			1158 => "00000000000000000001001001011101",
			1159 => "0000000000000000001101010000000100",
			1160 => "00000000000000000001001001011101",
			1161 => "00000001000010100001001001011101",
			1162 => "0000000101000000000110110100001000",
			1163 => "0000001001000000001101011000000100",
			1164 => "11111111000010110001001001011101",
			1165 => "00000000000000000001001001011101",
			1166 => "00000000000000000001001001011101",
			1167 => "0000001110000000001110101000001000",
			1168 => "0000001000000000000110001000000100",
			1169 => "00000001001000000001001001011101",
			1170 => "00000000000000000001001001011101",
			1171 => "00000000000000000001001001011101",
			1172 => "0000000111000000001101010100000100",
			1173 => "00000000000000000001001001011101",
			1174 => "11111111001000010001001001011101",
			1175 => "0000000001000000001101101000000100",
			1176 => "11111110011010010001001010100001",
			1177 => "0000001101000000000000110100011100",
			1178 => "0000000100000000001110111000000100",
			1179 => "11111110111110110001001010100001",
			1180 => "0000000101000000000101100100001000",
			1181 => "0000001100000000001100110000000100",
			1182 => "00000000000111000001001010100001",
			1183 => "00000001110100000001001010100001",
			1184 => "0000001001000000001010011000000100",
			1185 => "11111110100010000001001010100001",
			1186 => "0000001100000000000110000100000100",
			1187 => "00000000000000000001001010100001",
			1188 => "0000000001000000001101011100000100",
			1189 => "00000000000000000001001010100001",
			1190 => "00000001011011110001001010100001",
			1191 => "11111110011010100001001010100001",
			1192 => "0000000001000000001101101000000100",
			1193 => "11111110011011110001001011111101",
			1194 => "0000001110000000000111110000010100",
			1195 => "0000001000000000001000101100010000",
			1196 => "0000000010000000000111011000000100",
			1197 => "00000000000000000001001011111101",
			1198 => "0000000010000000001011101100001000",
			1199 => "0000001111000000000010000000000100",
			1200 => "00000001000010110001001011111101",
			1201 => "00000000000000000001001011111101",
			1202 => "00000001111110010001001011111101",
			1203 => "00000000000000000001001011111101",
			1204 => "0000001101000000000000110100010100",
			1205 => "0000000010000000001011111000001100",
			1206 => "0000001010000000000110011000001000",
			1207 => "0000000100000000001110111000000100",
			1208 => "00000000000000000001001011111101",
			1209 => "00000000100010000001001011111101",
			1210 => "11111110011100000001001011111101",
			1211 => "0000001111000000000111011000000100",
			1212 => "00000001011000010001001011111101",
			1213 => "00000000000000000001001011111101",
			1214 => "11111110100001010001001011111101",
			1215 => "0000000100000000000010100100000100",
			1216 => "11111110101101010001001101100001",
			1217 => "0000001110000000000111110000011100",
			1218 => "0000000001000000000110101000000100",
			1219 => "11111111100010110001001101100001",
			1220 => "0000001101000000000001011000001100",
			1221 => "0000000110000000001001100100001000",
			1222 => "0000001100000000001100110000000100",
			1223 => "00000000000000000001001101100001",
			1224 => "00000001001000110001001101100001",
			1225 => "00000000000000000001001101100001",
			1226 => "0000001010000000001100011100001000",
			1227 => "0000001111000000001001011100000100",
			1228 => "00000000000000000001001101100001",
			1229 => "00000000110100010001001101100001",
			1230 => "11111111101100000001001101100001",
			1231 => "0000001000000000001011010100001000",
			1232 => "0000000111000000001101010100000100",
			1233 => "00000000001111010001001101100001",
			1234 => "00000000000000000001001101100001",
			1235 => "0000001101000000000101110100000100",
			1236 => "00000000000000000001001101100001",
			1237 => "0000001011000000001000000000000100",
			1238 => "11111110111010000001001101100001",
			1239 => "00000000000000000001001101100001",
			1240 => "0000000010000000000111011000000100",
			1241 => "11111110011010100001001110101101",
			1242 => "0000001111000000001100000000100000",
			1243 => "0000001001000000001110010100000100",
			1244 => "11111110100111000001001110101101",
			1245 => "0000000010000000001011111000010100",
			1246 => "0000001000000000001011010100001000",
			1247 => "0000001110000000001110101100000100",
			1248 => "00000001100010000001001110101101",
			1249 => "11111111001101000001001110101101",
			1250 => "0000000101000000000101100100001000",
			1251 => "0000001001000000000100110100000100",
			1252 => "00000000000000000001001110101101",
			1253 => "00000000011000000001001110101101",
			1254 => "11111110000010000001001110101101",
			1255 => "0000001010000000000001010100000100",
			1256 => "00000001101111100001001110101101",
			1257 => "00000000000000000001001110101101",
			1258 => "11111110011011100001001110101101",
			1259 => "0000000001000000001101101000000100",
			1260 => "11111110011100010001010000010001",
			1261 => "0000001101000000000000110100101000",
			1262 => "0000000010000000001011111000011000",
			1263 => "0000001000000000001011010100010000",
			1264 => "0000000000000000001000110000000100",
			1265 => "11111111101101000001010000010001",
			1266 => "0000001111000000000010000000001000",
			1267 => "0000000001000000001111001100000100",
			1268 => "00000000000000000001010000010001",
			1269 => "00000001010011100001010000010001",
			1270 => "00000000000000000001010000010001",
			1271 => "0000000101000000000101100100000100",
			1272 => "00000000000000000001010000010001",
			1273 => "11111110100100110001010000010001",
			1274 => "0000001100000000001100110000000100",
			1275 => "00000000000000000001010000010001",
			1276 => "0000001000000000001000101100001000",
			1277 => "0000001111000000000111011000000100",
			1278 => "00000001100111110001010000010001",
			1279 => "00000000000000000001010000010001",
			1280 => "00000000000000000001010000010001",
			1281 => "0000000101000000001011110100000100",
			1282 => "00000000000000000001010000010001",
			1283 => "11111110100011000001010000010001",
			1284 => "0000000010000000001111010100001000",
			1285 => "0000000010000000000111011000000100",
			1286 => "11111110011101010001010010000101",
			1287 => "00000000000000000001010010000101",
			1288 => "0000000110000000001011001100010000",
			1289 => "0000000111000000001101010100001100",
			1290 => "0000000001000000000110101000000100",
			1291 => "00000000000000000001010010000101",
			1292 => "0000001100000000001100110000000100",
			1293 => "00000000000000000001010010000101",
			1294 => "00000010011011010001010010000101",
			1295 => "00000000000000000001010010000101",
			1296 => "0000001111000000001100000000100000",
			1297 => "0000000001000000001101011100010000",
			1298 => "0000001111000000001100010100001000",
			1299 => "0000001010000000000001010000000100",
			1300 => "00000000000000000001010010000101",
			1301 => "11111110110101010001010010000101",
			1302 => "0000001001000000001010011000000100",
			1303 => "00000000000000000001010010000101",
			1304 => "00000000010101000001010010000101",
			1305 => "0000000010000000001011111000001100",
			1306 => "0000000011000000001101000100000100",
			1307 => "00000000011011010001010010000101",
			1308 => "0000001100000000001110001100000100",
			1309 => "11111111011100000001010010000101",
			1310 => "00000000000000000001010010000101",
			1311 => "00000001010101100001010010000101",
			1312 => "11111110101101000001010010000101",
			1313 => "0000000010000000000111011000000100",
			1314 => "11111110011010100001010011110001",
			1315 => "0000001100000000001010111100101100",
			1316 => "0000000010000000001011111000011100",
			1317 => "0000001000000000001011010100001100",
			1318 => "0000001110000000001110101100001000",
			1319 => "0000000001000000001111001100000100",
			1320 => "00000000000000000001010011110001",
			1321 => "00000001100000010001010011110001",
			1322 => "11111111001001000001010011110001",
			1323 => "0000001100000000001110001100001000",
			1324 => "0000001010000000000110011000000100",
			1325 => "00000000000000000001010011110001",
			1326 => "11111110010010000001010011110001",
			1327 => "0000000011000000000010001000000100",
			1328 => "00000000000000000001010011110001",
			1329 => "00000000000001000001010011110001",
			1330 => "0000001010000000000001010100001100",
			1331 => "0000000100000000000011110100000100",
			1332 => "11111111100001100001010011110001",
			1333 => "0000001100000000000011011100000100",
			1334 => "00000000000000000001010011110001",
			1335 => "00000001101101110001010011110001",
			1336 => "11111111010001000001010011110001",
			1337 => "0000001100000000001010111100000100",
			1338 => "00000000000000000001010011110001",
			1339 => "11111110011100100001010011110001",
			1340 => "0000000100000000000011110100001100",
			1341 => "0000000100000000000011010100000100",
			1342 => "11111110011010100001010101110101",
			1343 => "0000000100000000000011010100000100",
			1344 => "11111111111000000001010101110101",
			1345 => "11111110111000110001010101110101",
			1346 => "0000001000000000000010101000100100",
			1347 => "0000001001000000001110010100000100",
			1348 => "11111110100011110001010101110101",
			1349 => "0000001110000000000111110000001100",
			1350 => "0000000101000000000101100100000100",
			1351 => "00000001110011100001010101110101",
			1352 => "0000000101000000000101100100000100",
			1353 => "11111111110011000001010101110101",
			1354 => "00000001101011010001010101110101",
			1355 => "0000001000000000001011010100001000",
			1356 => "0000000110000000001011001100000100",
			1357 => "00000000101010100001010101110101",
			1358 => "00000010001100110001010101110101",
			1359 => "0000000110000000001001100100000100",
			1360 => "11111101011110000001010101110101",
			1361 => "0000001110000000001110101100000100",
			1362 => "00000001010101110001010101110101",
			1363 => "11111111000100110001010101110101",
			1364 => "0000001010000000000001110000010000",
			1365 => "0000001001000000001011111100000100",
			1366 => "11111110011101100001010101110101",
			1367 => "0000000111000000001101111000000100",
			1368 => "00000100011010010001010101110101",
			1369 => "0000001010000000000101000100000100",
			1370 => "00000000000000000001010101110101",
			1371 => "11111111100000100001010101110101",
			1372 => "11111110011010000001010101110101",
			1373 => "0000000010000000000110111100000100",
			1374 => "11111110011001010001010111101001",
			1375 => "0000001100000000000100001000100100",
			1376 => "0000001100000000000011011100001000",
			1377 => "0000000111000000001101111000000100",
			1378 => "11111110011110010001010111101001",
			1379 => "00000000000000000001010111101001",
			1380 => "0000001010000000001100000100011000",
			1381 => "0000001110000000000001101000001000",
			1382 => "0000000010000000000110101100000100",
			1383 => "00000010101011110001010111101001",
			1384 => "00000111101110010001010111101001",
			1385 => "0000000101000000000101100100001000",
			1386 => "0000000001000000001111001100000100",
			1387 => "11111111001100110001010111101001",
			1388 => "00000001110111100001010111101001",
			1389 => "0000001001000000001010011000000100",
			1390 => "11111101001010110001010111101001",
			1391 => "00000001000111010001010111101001",
			1392 => "11111110100110000001010111101001",
			1393 => "0000000111000000000111001000001100",
			1394 => "0000000101000000000101100100000100",
			1395 => "11111111001000010001010111101001",
			1396 => "0000001100000000000100001000000100",
			1397 => "11111111101000000001010111101001",
			1398 => "00000001001010100001010111101001",
			1399 => "0000001100000000000100001000000100",
			1400 => "00000000000000000001010111101001",
			1401 => "11111110011001100001010111101001",
			1402 => "0000000001000000001101101000000100",
			1403 => "11111110011001100001011001110101",
			1404 => "0000001110000000001001010100100000",
			1405 => "0000000101000000000101100100010000",
			1406 => "0000001110000000001001001000000100",
			1407 => "00000011100001000001011001110101",
			1408 => "0000000100000000000000010100000100",
			1409 => "11111111011001000001011001110101",
			1410 => "0000001010000000000110011100000100",
			1411 => "00000001101110000001011001110101",
			1412 => "00000000000000000001011001110101",
			1413 => "0000000001000000001101011100001100",
			1414 => "0000001111000000001100010100001000",
			1415 => "0000001110000000001011011100000100",
			1416 => "00000000000000000001011001110101",
			1417 => "11111110010101110001011001110101",
			1418 => "00000000011001010001011001110101",
			1419 => "00000001100101010001011001110101",
			1420 => "0000001101000000000000110100100000",
			1421 => "0000001100000000001110001100010100",
			1422 => "0000001000000000001011010100001000",
			1423 => "0000000100000000000110001100000100",
			1424 => "11111111001000110001011001110101",
			1425 => "00000000010010100001011001110101",
			1426 => "0000001101000000000100010000001000",
			1427 => "0000000101000000000100000100000100",
			1428 => "11111111100001000001011001110101",
			1429 => "00000000000000010001011001110101",
			1430 => "11111101010101100001011001110101",
			1431 => "0000000100000000000000010100000100",
			1432 => "11111111001010100001011001110101",
			1433 => "0000001001000000001111000000000100",
			1434 => "00000000010011010001011001110101",
			1435 => "00000010001101100001011001110101",
			1436 => "11111110011000100001011001110101",
			1437 => "0000000010000000001111010100000100",
			1438 => "11111110011010000001011011111011",
			1439 => "0000001100000000000100001000110000",
			1440 => "0000001001000000001110010100000100",
			1441 => "11111110011111110001011011111011",
			1442 => "0000001110000000001001010100010100",
			1443 => "0000001000000000001000101100010000",
			1444 => "0000000001000000001111001100001000",
			1445 => "0000001111000000001110010000000100",
			1446 => "00000011000100110001011011111011",
			1447 => "00000001000101010001011011111011",
			1448 => "0000000001000000001101011100000100",
			1449 => "00000000000111010001011011111011",
			1450 => "00000001101010100001011011111011",
			1451 => "11111110110010000001011011111011",
			1452 => "0000000001000000001001011000001100",
			1453 => "0000001000000000001100000100000100",
			1454 => "00000000000000000001011011111011",
			1455 => "0000001011000000000100011000000100",
			1456 => "11111110111110010001011011111011",
			1457 => "11111100110001110001011011111011",
			1458 => "0000001110000000001110101000001000",
			1459 => "0000001100000000001110001100000100",
			1460 => "00000000011101110001011011111011",
			1461 => "00000010111101110001011011111011",
			1462 => "11111110110011010001011011111011",
			1463 => "0000000111000000000111001000001100",
			1464 => "0000001110000000000111110000001000",
			1465 => "0000001110000000001000110000000100",
			1466 => "11111111101010100001011011111011",
			1467 => "00000000110101000001011011111011",
			1468 => "11111110101111000001011011111011",
			1469 => "11111110011001110001011011111011",
			1470 => "00000000000000000001011011111101",
			1471 => "00000000000000000001011100000001",
			1472 => "00000000000000000001011100000101",
			1473 => "00000000000000000001011100001001",
			1474 => "00000000000000000001011100001101",
			1475 => "00000000000000000001011100010001",
			1476 => "00000000000000000001011100010101",
			1477 => "00000000000000000001011100011001",
			1478 => "00000000000000000001011100011101",
			1479 => "00000000000000000001011100100001",
			1480 => "00000000000000000001011100100101",
			1481 => "00000000000000000001011100101001",
			1482 => "00000000000000000001011100101101",
			1483 => "00000000000000000001011100110001",
			1484 => "00000000000000000001011100110101",
			1485 => "00000000000000000001011100111001",
			1486 => "00000000000000000001011100111101",
			1487 => "00000000000000000001011101000001",
			1488 => "00000000000000000001011101000101",
			1489 => "00000000000000000001011101001001",
			1490 => "00000000000000000001011101001101",
			1491 => "00000000000000000001011101010001",
			1492 => "00000000000000000001011101010101",
			1493 => "00000000000000000001011101011001",
			1494 => "00000000000000000001011101011101",
			1495 => "00000000000000000001011101100001",
			1496 => "00000000000000000001011101100101",
			1497 => "00000000000000000001011101101001",
			1498 => "00000000000000000001011101101101",
			1499 => "0000000100000000000100111000000100",
			1500 => "11111111111111110001011101111001",
			1501 => "00000000000000000001011101111001",
			1502 => "0000000100000000000011011000000100",
			1503 => "11111111111101100001011110000101",
			1504 => "00000000000000000001011110000101",
			1505 => "0000000010000000000110101100000100",
			1506 => "11111111111011110001011110010001",
			1507 => "00000000000000000001011110010001",
			1508 => "0000000000000000001100001000000100",
			1509 => "11111111111111010001011110011101",
			1510 => "00000000000000000001011110011101",
			1511 => "0000000001000000001111001100000100",
			1512 => "11111111111010010001011110101001",
			1513 => "00000000000000000001011110101001",
			1514 => "0000000100000000000011111000000100",
			1515 => "11111111111100010001011110110101",
			1516 => "00000000000000000001011110110101",
			1517 => "0000000010000000001011111000001000",
			1518 => "0000000001000000000000111100000100",
			1519 => "11111111101000100001011111001001",
			1520 => "00000000000000000001011111001001",
			1521 => "00000000000000000001011111001001",
			1522 => "0000000100000000000000010100000100",
			1523 => "11111111111101000001011111011101",
			1524 => "0000000100000000001010010000000100",
			1525 => "00000000000000110001011111011101",
			1526 => "00000000000000000001011111011101",
			1527 => "0000000010000000000110101100000100",
			1528 => "11111111111100010001011111110001",
			1529 => "0000000010000000001101101100000100",
			1530 => "00000000000010100001011111110001",
			1531 => "00000000000000000001011111110001",
			1532 => "0000000100000000000010100100000100",
			1533 => "00000000000000000001100000000101",
			1534 => "0000000100000000001010010000000100",
			1535 => "00000000000011000001100000000101",
			1536 => "00000000000000000001100000000101",
			1537 => "0000000010000000001011111000000100",
			1538 => "11111111111111110001100000011001",
			1539 => "0000000010000000001100111000000100",
			1540 => "00000000001010000001100000011001",
			1541 => "00000000000000000001100000011001",
			1542 => "0000000010000000000110101100000100",
			1543 => "11111111111111000001100000101101",
			1544 => "0000000010000000001111101000000100",
			1545 => "00000000000111010001100000101101",
			1546 => "00000000000000000001100000101101",
			1547 => "0000000001000000001101011100001000",
			1548 => "0000000100000000000100111000000100",
			1549 => "11111111110011000001100001000001",
			1550 => "00000000000000000001100001000001",
			1551 => "00000000000000000001100001000001",
			1552 => "0000000100000000000011111000001100",
			1553 => "0000000001000000001101011100001000",
			1554 => "0000001001000000001101011000000100",
			1555 => "11111111011010110001100001011101",
			1556 => "00000000000000000001100001011101",
			1557 => "00000000000000000001100001011101",
			1558 => "00000000000000000001100001011101",
			1559 => "0000000100000000000101100000001100",
			1560 => "0000000001000000001101011100001000",
			1561 => "0000001001000000001101011000000100",
			1562 => "11111111100111010001100001111001",
			1563 => "00000000000000000001100001111001",
			1564 => "00000000000000000001100001111001",
			1565 => "00000000000000000001100001111001",
			1566 => "0000000100000000000010100100000100",
			1567 => "11111111111101010001100010010101",
			1568 => "0000000010000000000000010000000100",
			1569 => "00000000000000000001100010010101",
			1570 => "0000000010000000001111101000000100",
			1571 => "00000000000110000001100010010101",
			1572 => "00000000000000000001100010010101",
			1573 => "0000001001000000001101011000001100",
			1574 => "0000000100000000000100111000001000",
			1575 => "0000000001000000001101011100000100",
			1576 => "11111111101110010001100010110001",
			1577 => "00000000000000000001100010110001",
			1578 => "00000000000000000001100010110001",
			1579 => "00000000000000000001100010110001",
			1580 => "0000001001000000001010011000001000",
			1581 => "0000000100000000000100111000000100",
			1582 => "11111111000010110001100011010101",
			1583 => "00000000000000000001100011010101",
			1584 => "0000001110000000001001010100001000",
			1585 => "0000000101000000000100010000000100",
			1586 => "00000000100001100001100011010101",
			1587 => "00000000000000000001100011010101",
			1588 => "00000000000000000001100011010101",
			1589 => "0000000001000000001111001100000100",
			1590 => "11111111010101110001100011111001",
			1591 => "0000000111000000001101010100001100",
			1592 => "0000001110000000001110101000001000",
			1593 => "0000001100000000000000001100000100",
			1594 => "00000000100000000001100011111001",
			1595 => "00000000000000000001100011111001",
			1596 => "00000000000000000001100011111001",
			1597 => "00000000000000000001100011111001",
			1598 => "0000000100000000000011010100000100",
			1599 => "11111111111100010001100100011101",
			1600 => "0000000010000000000110101100000100",
			1601 => "00000000000000000001100100011101",
			1602 => "0000000010000000000011000000001000",
			1603 => "0000000100000000001010010000000100",
			1604 => "00000000010011100001100100011101",
			1605 => "00000000000000000001100100011101",
			1606 => "00000000000000000001100100011101",
			1607 => "0000000100000000000010100100000100",
			1608 => "00000000000000000001100101000001",
			1609 => "0000000010000000001100111000001100",
			1610 => "0000000010000000000000010000000100",
			1611 => "00000000000000000001100101000001",
			1612 => "0000000100000000001010010000000100",
			1613 => "00000000001101110001100101000001",
			1614 => "00000000000000000001100101000001",
			1615 => "00000000000000000001100101000001",
			1616 => "0000001001000000001010011000001000",
			1617 => "0000000100000000000100111000000100",
			1618 => "11111111001101010001100101101101",
			1619 => "00000000000000000001100101101101",
			1620 => "0000001110000000001110101000001100",
			1621 => "0000000010000000001011111000000100",
			1622 => "00000000000000000001100101101101",
			1623 => "0000001100000000000100001000000100",
			1624 => "00000000100011000001100101101101",
			1625 => "00000000000000000001100101101101",
			1626 => "00000000000000000001100101101101",
			1627 => "0000000001000000001111001100001000",
			1628 => "0000000100000000000100111000000100",
			1629 => "11111111100011100001100110011001",
			1630 => "00000000000000000001100110011001",
			1631 => "0000001110000000000111110000001100",
			1632 => "0000000111000000001101111000000100",
			1633 => "00000000000000000001100110011001",
			1634 => "0000000110000000001001100100000100",
			1635 => "00000000010101010001100110011001",
			1636 => "00000000000000000001100110011001",
			1637 => "00000000000000000001100110011001",
			1638 => "0000000100000000000011110100000100",
			1639 => "11111111011100000001100111000101",
			1640 => "0000001011000000000011100000001000",
			1641 => "0000000001000000001111001100000100",
			1642 => "00000000000000000001100111000101",
			1643 => "00000000100000100001100111000101",
			1644 => "0000001000000000001011010100000100",
			1645 => "00000000000000000001100111000101",
			1646 => "0000001111000000000011001000000100",
			1647 => "00000000000000000001100111000101",
			1648 => "11111111110010110001100111000101",
			1649 => "0000000010000000000110101100010000",
			1650 => "0000000000000000000011111100000100",
			1651 => "00000000000000000001101000000001",
			1652 => "0000000110000000001001100100001000",
			1653 => "0000001100000000000000001100000100",
			1654 => "11111111010100110001101000000001",
			1655 => "00000000000000000001101000000001",
			1656 => "00000000000000000001101000000001",
			1657 => "0000001111000000001100010000001100",
			1658 => "0000001010000000000001110000001000",
			1659 => "0000000111000000001110001100000100",
			1660 => "00000000000000000001101000000001",
			1661 => "00000000101010000001101000000001",
			1662 => "00000000000000000001101000000001",
			1663 => "00000000000000000001101000000001",
			1664 => "0000000010000000001011111000001000",
			1665 => "0000001000000000001011010100000100",
			1666 => "00000000000000000001101000110101",
			1667 => "11111111011000010001101000110101",
			1668 => "0000001111000000001100000000010000",
			1669 => "0000000111000000000110000100000100",
			1670 => "00000000000000000001101000110101",
			1671 => "0000001010000000001100000100001000",
			1672 => "0000000010000000000110101100000100",
			1673 => "00000000000000000001101000110101",
			1674 => "00000000011100000001101000110101",
			1675 => "00000000000000000001101000110101",
			1676 => "00000000000000000001101000110101",
			1677 => "0000000001000000001101101000000100",
			1678 => "11111111101001010001101001100001",
			1679 => "0000001110000000001110101100010000",
			1680 => "0000001100000000000100001000001100",
			1681 => "0000001111000000001111010000000100",
			1682 => "00000000000000000001101001100001",
			1683 => "0000001100000000000110000100000100",
			1684 => "00000000000000000001101001100001",
			1685 => "00000000001000010001101001100001",
			1686 => "00000000000000000001101001100001",
			1687 => "00000000000000000001101001100001",
			1688 => "0000000010000000001000001100001100",
			1689 => "0000000111000000001100101000001000",
			1690 => "0000001100000000001110001100000100",
			1691 => "11111110110101010001101010100101",
			1692 => "00000000000000000001101010100101",
			1693 => "00000000000000000001101010100101",
			1694 => "0000001111000000000011001000001100",
			1695 => "0000001000000000001010101100001000",
			1696 => "0000000001000000001011101000000100",
			1697 => "00000000000000000001101010100101",
			1698 => "00000000111001100001101010100101",
			1699 => "00000000000000000001101010100101",
			1700 => "0000001110000000001110101100001000",
			1701 => "0000000001000000001101011100000100",
			1702 => "11111111111010100001101010100101",
			1703 => "00000000010011000001101010100101",
			1704 => "11111111101000100001101010100101",
			1705 => "0000000010000000000111011000000100",
			1706 => "11111110110000010001101011100001",
			1707 => "0000000110000000001011001100001100",
			1708 => "0000000001000000000110101000000100",
			1709 => "00000000000000000001101011100001",
			1710 => "0000001110000000001110101100000100",
			1711 => "00000000110110110001101011100001",
			1712 => "00000000000000000001101011100001",
			1713 => "0000001001000000001010011000000100",
			1714 => "11111111000101100001101011100001",
			1715 => "0000001110000000001001010100000100",
			1716 => "00000000011101110001101011100001",
			1717 => "0000000110000000001011001100000100",
			1718 => "00000000000000000001101011100001",
			1719 => "11111111101011110001101011100001",
			1720 => "0000000010000000001011111000001100",
			1721 => "0000001000000000001011010100000100",
			1722 => "00000000000000000001101100100101",
			1723 => "0000001100000000000000001100000100",
			1724 => "11111111010011000001101100100101",
			1725 => "00000000000000000001101100100101",
			1726 => "0000001111000000001100000000010100",
			1727 => "0000001100000000000110000100000100",
			1728 => "00000000000000000001101100100101",
			1729 => "0000001100000000000100001000001100",
			1730 => "0000000110000000001001100100001000",
			1731 => "0000000001000000000110101000000100",
			1732 => "00000000000000000001101100100101",
			1733 => "00000000101010110001101100100101",
			1734 => "00000000000000000001101100100101",
			1735 => "00000000000000000001101100100101",
			1736 => "00000000000000000001101100100101",
			1737 => "0000000100000000001011100000000100",
			1738 => "11111110111010110001101101101001",
			1739 => "0000000010000000000110101100010000",
			1740 => "0000001000000000001011010100001100",
			1741 => "0000001111000000000010000000001000",
			1742 => "0000000001000000001111001100000100",
			1743 => "00000000000000000001101101101001",
			1744 => "00000000001110110001101101101001",
			1745 => "00000000000000000001101101101001",
			1746 => "11111111100010000001101101101001",
			1747 => "0000000110000000000100111100001100",
			1748 => "0000001010000000001100000100001000",
			1749 => "0000000001000000000110101000000100",
			1750 => "00000000000000000001101101101001",
			1751 => "00000000011001010001101101101001",
			1752 => "00000000000000000001101101101001",
			1753 => "00000000000000000001101101101001",
			1754 => "0000000010000000001000001100001100",
			1755 => "0000001100000000001110001100001000",
			1756 => "0000000111000000001100101000000100",
			1757 => "11111110101010100001101110110101",
			1758 => "00000000000000000001101110110101",
			1759 => "00000000000000000001101110110101",
			1760 => "0000001111000000001100000000011000",
			1761 => "0000000001000000001111001100010000",
			1762 => "0000000110000000001101011000001100",
			1763 => "0000000100000000001111101100001000",
			1764 => "0000000100000000000011111000000100",
			1765 => "00000000000000000001101110110101",
			1766 => "00000000011010110001101110110101",
			1767 => "00000000000000000001101110110101",
			1768 => "11111111101001010001101110110101",
			1769 => "0000000010000000001011111000000100",
			1770 => "00000000000000000001101110110101",
			1771 => "00000000111010110001101110110101",
			1772 => "11111111011100100001101110110101",
			1773 => "0000000100000000001001000000001000",
			1774 => "0000001001000000001010011000000100",
			1775 => "11111110101101110001110000010001",
			1776 => "00000000000000000001110000010001",
			1777 => "0000000010000000000110101100010000",
			1778 => "0000001000000000001011010100001100",
			1779 => "0000001111000000000010000000001000",
			1780 => "0000001111000000000101110000000100",
			1781 => "00000000000000000001110000010001",
			1782 => "00000000001010100001110000010001",
			1783 => "00000000000000000001110000010001",
			1784 => "11111111011100110001110000010001",
			1785 => "0000001100000000000110000100001100",
			1786 => "0000000001000000001101011100001000",
			1787 => "0000000001000000001101101000000100",
			1788 => "00000000000000000001110000010001",
			1789 => "11111111110110010001110000010001",
			1790 => "00000000000000000001110000010001",
			1791 => "0000001111000000000111011000001000",
			1792 => "0000001010000000001100000100000100",
			1793 => "00000000101110010001110000010001",
			1794 => "00000000000000000001110000010001",
			1795 => "00000000000000000001110000010001",
			1796 => "0000000001000000000110101000000100",
			1797 => "11111111001101010001110001011101",
			1798 => "0000000011000000001101000100010100",
			1799 => "0000001100000000000100001000010000",
			1800 => "0000000111000000000110000100000100",
			1801 => "00000000000000000001110001011101",
			1802 => "0000000100000000000000010100000100",
			1803 => "00000000000000000001110001011101",
			1804 => "0000001010000000001100000100000100",
			1805 => "00000000110000110001110001011101",
			1806 => "00000000000000000001110001011101",
			1807 => "00000000000000000001110001011101",
			1808 => "0000001001000000001111000000001000",
			1809 => "0000001101000000000101110100000100",
			1810 => "00000000000000000001110001011101",
			1811 => "11111111110001010001110001011101",
			1812 => "0000001011000000000110100100000100",
			1813 => "00000000000000110001110001011101",
			1814 => "00000000000000000001110001011101",
			1815 => "0000000010000000000000010000001100",
			1816 => "0000001001000000001111000000001000",
			1817 => "0000001100000000001110001100000100",
			1818 => "11111110101010010001110010110001",
			1819 => "00000000000000000001110010110001",
			1820 => "00000000000000000001110010110001",
			1821 => "0000001111000000000010000100011000",
			1822 => "0000000010000000000110101100000100",
			1823 => "00000000000000000001110010110001",
			1824 => "0000001100000000001100110000000100",
			1825 => "00000000000000000001110010110001",
			1826 => "0000001010000000001100000100001100",
			1827 => "0000001110000000001001010100001000",
			1828 => "0000000110000000001001100100000100",
			1829 => "00000001001011010001110010110001",
			1830 => "00000000000000000001110010110001",
			1831 => "00000000000000000001110010110001",
			1832 => "00000000000000000001110010110001",
			1833 => "0000001111000000001100000000000100",
			1834 => "00000000000000000001110010110001",
			1835 => "11111111010110100001110010110001",
			1836 => "0000001011000000000011100000011100",
			1837 => "0000001100000000000011011100000100",
			1838 => "00000000000000000001110011111101",
			1839 => "0000001111000000001001100000010100",
			1840 => "0000000010000000000111011000000100",
			1841 => "00000000000000000001110011111101",
			1842 => "0000000100000000001010010000001100",
			1843 => "0000001101000000001000011000000100",
			1844 => "00000000000000000001110011111101",
			1845 => "0000000010000000001000101000000100",
			1846 => "00000000010011110001110011111101",
			1847 => "00000000000000000001110011111101",
			1848 => "00000000000000000001110011111101",
			1849 => "00000000000000000001110011111101",
			1850 => "0000001111000000000011001000000100",
			1851 => "00000000000000000001110011111101",
			1852 => "0000001101000000000101110100000100",
			1853 => "00000000000000000001110011111101",
			1854 => "11111111110000010001110011111101",
			1855 => "0000000001000000000110101000000100",
			1856 => "11111111001011100001110101000001",
			1857 => "0000001111000000001100010000011100",
			1858 => "0000001000000000000110001000001000",
			1859 => "0000000100000000001110111000000100",
			1860 => "00000000000000000001110101000001",
			1861 => "00000000100100010001110101000001",
			1862 => "0000000100000000000100111000001100",
			1863 => "0000001011000000001000000000001000",
			1864 => "0000000010000000001100111000000100",
			1865 => "11111111100111100001110101000001",
			1866 => "00000000000000000001110101000001",
			1867 => "00000000000000000001110101000001",
			1868 => "0000001011000000001010111100000100",
			1869 => "00000000000000100001110101000001",
			1870 => "00000000000000000001110101000001",
			1871 => "11111111111011100001110101000001",
			1872 => "0000000010000000000000010000010100",
			1873 => "0000000001000000001111001100000100",
			1874 => "11111110011101100001110110101101",
			1875 => "0000001011000000000011100000001100",
			1876 => "0000000010000000000000010000001000",
			1877 => "0000001100000000000011011100000100",
			1878 => "00000000000000000001110110101101",
			1879 => "00000000111111000001110110101101",
			1880 => "00000000000000000001110110101101",
			1881 => "11111110100010010001110110101101",
			1882 => "0000000110000000001011001100010000",
			1883 => "0000000001000000000110101000000100",
			1884 => "00000000000000000001110110101101",
			1885 => "0000000011000000000011001000001000",
			1886 => "0000001100000000000110000100000100",
			1887 => "00000000000000000001110110101101",
			1888 => "00000010011000000001110110101101",
			1889 => "00000000000000000001110110101101",
			1890 => "0000000011000000001001011100010000",
			1891 => "0000001001000000001010011000000100",
			1892 => "11111111000101000001110110101101",
			1893 => "0000000010000000001011111000001000",
			1894 => "0000001101000000000101110100000100",
			1895 => "00000000000000000001110110101101",
			1896 => "11111111101101010001110110101101",
			1897 => "00000001010100100001110110101101",
			1898 => "11111110110010010001110110101101",
			1899 => "0000000111000000000110000100001000",
			1900 => "0000001100000000000110000100000100",
			1901 => "11111111001111100001111000001001",
			1902 => "00000000000000000001111000001001",
			1903 => "0000000011000000001101000100011000",
			1904 => "0000001100000000000100001000010100",
			1905 => "0000001001000000001101011100000100",
			1906 => "00000000000000000001111000001001",
			1907 => "0000000100000000000000010100000100",
			1908 => "00000000000000000001111000001001",
			1909 => "0000000000000000001100101100001000",
			1910 => "0000000010000000001000101000000100",
			1911 => "00000000101100100001111000001001",
			1912 => "00000000000000000001111000001001",
			1913 => "00000000000000000001111000001001",
			1914 => "00000000000000000001111000001001",
			1915 => "0000001011000000000011100000000100",
			1916 => "00000000000000000001111000001001",
			1917 => "0000000110000000001001100100001000",
			1918 => "0000001001000000000100111100000100",
			1919 => "11111111110001010001111000001001",
			1920 => "00000000000000000001111000001001",
			1921 => "00000000000000000001111000001001",
			1922 => "0000000100000000000011110100000100",
			1923 => "11111110011011010001111001100101",
			1924 => "0000000001000000001111001100001100",
			1925 => "0000000001000000001101101000000100",
			1926 => "11111110011010110001111001100101",
			1927 => "0000000110000000001011001100000100",
			1928 => "00000010001100000001111001100101",
			1929 => "11111110011111000001111001100101",
			1930 => "0000001110000000001001010100010000",
			1931 => "0000000000000000001110111100000100",
			1932 => "00000001101010110001111001100101",
			1933 => "0000000010000000001011101100000100",
			1934 => "11111111101001010001111001100101",
			1935 => "0000000010000000000001011100000100",
			1936 => "00000010010111000001111001100101",
			1937 => "00000000001010110001111001100101",
			1938 => "0000001000000000001011010100000100",
			1939 => "00000001001010010001111001100101",
			1940 => "0000000001000000000000111100000100",
			1941 => "11111110000111000001111001100101",
			1942 => "0000000001000000000101011100000100",
			1943 => "00000000000101000001111001100101",
			1944 => "11111111000100100001111001100101",
			1945 => "0000000100000000000010100100001000",
			1946 => "0000000100000000000011110100000100",
			1947 => "11111110100100110001111011100001",
			1948 => "00000000000000000001111011100001",
			1949 => "0000000010000000000110101100011100",
			1950 => "0000001000000000001011010100001100",
			1951 => "0000000001000000001111001100000100",
			1952 => "00000000000000000001111011100001",
			1953 => "0000001111000000001100010100000100",
			1954 => "00000000101011110001111011100001",
			1955 => "00000000000000000001111011100001",
			1956 => "0000000110000000001001100100001100",
			1957 => "0000001011000000001000000000001000",
			1958 => "0000001010000000000110011000000100",
			1959 => "00000000000000000001111011100001",
			1960 => "11111110111100100001111011100001",
			1961 => "00000000000000000001111011100001",
			1962 => "00000000000000000001111011100001",
			1963 => "0000001101000000000001011000001100",
			1964 => "0000001010000000001100000100001000",
			1965 => "0000001100000000001100110000000100",
			1966 => "00000000000000000001111011100001",
			1967 => "00000001110010000001111011100001",
			1968 => "00000000000000000001111011100001",
			1969 => "0000000001000000001101011100001000",
			1970 => "0000001110000000000100010000000100",
			1971 => "00000000000000000001111011100001",
			1972 => "11111111010001010001111011100001",
			1973 => "0000001101000000001110101100000100",
			1974 => "00000000111011100001111011100001",
			1975 => "00000000000000000001111011100001",
			1976 => "0000000100000000000010100100000100",
			1977 => "11111110110100010001111100111101",
			1978 => "0000001110000000001001010100011100",
			1979 => "0000000001000000001111001100011000",
			1980 => "0000000100000000000100111000001000",
			1981 => "0000001100000000001110001100000100",
			1982 => "11111111011110100001111100111101",
			1983 => "00000000000000000001111100111101",
			1984 => "0000001010000000001100000100001100",
			1985 => "0000001101000000001010001100001000",
			1986 => "0000001111000000000111110000000100",
			1987 => "00000000000000000001111100111101",
			1988 => "00000000010011000001111100111101",
			1989 => "00000000000000000001111100111101",
			1990 => "00000000000000000001111100111101",
			1991 => "00000000111001010001111100111101",
			1992 => "0000001100000000001110001100001000",
			1993 => "0000001100000000001100110000000100",
			1994 => "00000000000000000001111100111101",
			1995 => "11111111001011000001111100111101",
			1996 => "0000001111000000000111011000000100",
			1997 => "00000000001011010001111100111101",
			1998 => "00000000000000000001111100111101",
			1999 => "0000000010000000001111010100001100",
			2000 => "0000000010000000000111011000000100",
			2001 => "11111110011011010001111111001001",
			2002 => "0000000010000000000110111100000100",
			2003 => "00000000000000000001111111001001",
			2004 => "11111111100110000001111111001001",
			2005 => "0000001100000000000100001000101100",
			2006 => "0000000010000000000110101100011000",
			2007 => "0000001000000000001011010100001100",
			2008 => "0000001110000000001110101100001000",
			2009 => "0000001100000000001100110000000100",
			2010 => "00000000000000000001111111001001",
			2011 => "00000001011000100001111111001001",
			2012 => "11111111010111110001111111001001",
			2013 => "0000001100000000001110001100001000",
			2014 => "0000000010000000001011111000000100",
			2015 => "11111110100011010001111111001001",
			2016 => "00000000000000000001111111001001",
			2017 => "00000000000000000001111111001001",
			2018 => "0000001100000000001100110000001000",
			2019 => "0000001010000000001010110000000100",
			2020 => "00000000000000000001111111001001",
			2021 => "11111111100000010001111111001001",
			2022 => "0000001010000000000001110000001000",
			2023 => "0000000011000000001001011100000100",
			2024 => "00000001101101110001111111001001",
			2025 => "00000000000000000001111111001001",
			2026 => "11111111110110100001111111001001",
			2027 => "0000000111000000001110110000001100",
			2028 => "0000001011000000001000000000000100",
			2029 => "11111111011001100001111111001001",
			2030 => "0000001110000000001001010000000100",
			2031 => "00000000000111000001111111001001",
			2032 => "00000000000000000001111111001001",
			2033 => "11111110100000010001111111001001",
			2034 => "0000001001000000001010011000101000",
			2035 => "0000000001000000001101011100100100",
			2036 => "0000000001000000001111001100011000",
			2037 => "0000000010000000001011111000000100",
			2038 => "11111110011000010010000001000101",
			2039 => "0000000010000000000110101100001000",
			2040 => "0000000001000000000110000000000100",
			2041 => "11111111011010000010000001000101",
			2042 => "00001011001110010010000001000101",
			2043 => "0000001011000000001010111100001000",
			2044 => "0000001100000000000110000100000100",
			2045 => "11111110100100000010000001000101",
			2046 => "00011000011111110010000001000101",
			2047 => "11111110011001000010000001000101",
			2048 => "0000001101000000000101100100001000",
			2049 => "0000000000000000000010011000000100",
			2050 => "11111111001000100010000001000101",
			2051 => "00001000010000110010000001000101",
			2052 => "11111110010101010010000001000101",
			2053 => "11111100010101010010000001000101",
			2054 => "0000001110000000001110101000010100",
			2055 => "0000001001000000000100111100010000",
			2056 => "0000001110000000000111110000001000",
			2057 => "0000000001000000001101011100000100",
			2058 => "00000010110001110010000001000101",
			2059 => "00000001111000100010000001000101",
			2060 => "0000000101000000001011011100000100",
			2061 => "00000001110010010010000001000101",
			2062 => "11111110001100110010000001000101",
			2063 => "00000101100000100010000001000101",
			2064 => "11111110011000100010000001000101",
			2065 => "0000000001000000001101101000000100",
			2066 => "11111110011011000010000010111001",
			2067 => "0000001100000000000100001000101100",
			2068 => "0000001110000000001001010100011100",
			2069 => "0000001101000000000010001000001100",
			2070 => "0000001111000000001001010000000100",
			2071 => "00000000000000000010000010111001",
			2072 => "0000001011000000000001111100000100",
			2073 => "00000000000000000010000010111001",
			2074 => "00000001110111000010000010111001",
			2075 => "0000000100000000000010010000001000",
			2076 => "0000000000000000001000110000000100",
			2077 => "00000000000000000010000010111001",
			2078 => "00000001011010110010000010111001",
			2079 => "0000001111000000000010000000000100",
			2080 => "11111110110111000010000010111001",
			2081 => "00000000000000000010000010111001",
			2082 => "0000001100000000001110001100001000",
			2083 => "0000001010000000000110011000000100",
			2084 => "00000000000000000010000010111001",
			2085 => "11111110001110010010000010111001",
			2086 => "0000001110000000001110101000000100",
			2087 => "00000001010100110010000010111001",
			2088 => "00000000000000000010000010111001",
			2089 => "0000000101000000000100010000000100",
			2090 => "00000000000000000010000010111001",
			2091 => "0000001100000000000100001000000100",
			2092 => "00000000000000000010000010111001",
			2093 => "11111110011111010010000010111001",
			2094 => "0000000010000000001111010100001100",
			2095 => "0000000010000000000111011000000100",
			2096 => "11111110011001110010000100110101",
			2097 => "0000000010000000000110111100000100",
			2098 => "00000000000000000010000100110101",
			2099 => "11111111000000100010000100110101",
			2100 => "0000001100000000001010111100101100",
			2101 => "0000001110000000001001010100010100",
			2102 => "0000001001000000001110010100000100",
			2103 => "11111110101000000010000100110101",
			2104 => "0000001010000000000001010100001100",
			2105 => "0000001100000000000100001000001000",
			2106 => "0000000000000000000100000000000100",
			2107 => "00000001011011100010000100110101",
			2108 => "00000010111001000010000100110101",
			2109 => "00000000000000000010000100110101",
			2110 => "11111111001001100010000100110101",
			2111 => "0000001000000000001011010100001000",
			2112 => "0000000100000000001110111000000100",
			2113 => "11111111000000000010000100110101",
			2114 => "00000001001100000010000100110101",
			2115 => "0000000010000000000110101100000100",
			2116 => "11111101101110100010000100110101",
			2117 => "0000000001000000001001011000000100",
			2118 => "11111110111110100010000100110101",
			2119 => "0000001001000000001000010000000100",
			2120 => "00000000110111010010000100110101",
			2121 => "00000000000000000010000100110101",
			2122 => "0000000111000000000111001000000100",
			2123 => "00000000000000000010000100110101",
			2124 => "11111110011000100010000100110101",
			2125 => "0000000010000000001111010100000100",
			2126 => "11111110011001000010000110101001",
			2127 => "0000001100000000000100001000100100",
			2128 => "0000000001000000001101101000001100",
			2129 => "0000001100000000000110000100000100",
			2130 => "11111110011100010010000110101001",
			2131 => "0000000111000000001101111000000100",
			2132 => "00000101111011100010000110101001",
			2133 => "11111110110011000010000110101001",
			2134 => "0000001110000000001000011000000100",
			2135 => "00001011110111110010000110101001",
			2136 => "0000001000000000000001110100001100",
			2137 => "0000001110000000001110101000001000",
			2138 => "0000001110000000001110101100000100",
			2139 => "00000001101110010010000110101001",
			2140 => "00000110111100110010000110101001",
			2141 => "11111110100100100010000110101001",
			2142 => "0000000110000000001111000000000100",
			2143 => "11111100111010000010000110101001",
			2144 => "11111110110010100010000110101001",
			2145 => "0000000111000000000111001000010000",
			2146 => "0000001011000000001000000000001000",
			2147 => "0000000111000000000111001000000100",
			2148 => "11111110001110010010000110101001",
			2149 => "00000000000000000010000110101001",
			2150 => "0000000011000000000111100000000100",
			2151 => "00000001100101000010000110101001",
			2152 => "11111111001110110010000110101001",
			2153 => "11111110011000010010000110101001",
			2154 => "0000000010000000001111010100001000",
			2155 => "0000000010000000000111011000000100",
			2156 => "11111110011000110010001000010101",
			2157 => "11111110110110010010001000010101",
			2158 => "0000001110000000001110101000101100",
			2159 => "0000000001000000001101101000001100",
			2160 => "0000000001000000000110101000000100",
			2161 => "11111110011011000010001000010101",
			2162 => "0000000001000000000110101000000100",
			2163 => "00000111110001100010001000010101",
			2164 => "11111110100101100010001000010101",
			2165 => "0000001110000000000001101000001000",
			2166 => "0000001000000000001000110000000100",
			2167 => "00001001001011010010001000010101",
			2168 => "00000010101001100010001000010101",
			2169 => "0000001000000000000001110100010000",
			2170 => "0000000001000000001111001100001000",
			2171 => "0000001111000000000010000000000100",
			2172 => "00000100000110110010001000010101",
			2173 => "11111111100000010010001000010101",
			2174 => "0000000001000000001101011100000100",
			2175 => "00000000001000100010001000010101",
			2176 => "00000001101100110010001000010101",
			2177 => "0000000110000000001001100100000100",
			2178 => "00000000000000000010001000010101",
			2179 => "11111101110110100010001000010101",
			2180 => "11111110011001000010001000010101",
			2181 => "0000000010000000001111010100001000",
			2182 => "0000000010000000001111010100000100",
			2183 => "11111110011110000010001010001001",
			2184 => "00000000000000000010001010001001",
			2185 => "0000001110000000001100101100001000",
			2186 => "0000000011000000001011000000000100",
			2187 => "00000000000000000010001010001001",
			2188 => "00010010111101100010001010001001",
			2189 => "0000000110000000001011001100001100",
			2190 => "0000001011000000001001001000001000",
			2191 => "0000000001000000001101101000000100",
			2192 => "00000000000000000010001010001001",
			2193 => "00000001111101100010001010001001",
			2194 => "00000000000000000010001010001001",
			2195 => "0000001110000000001110101000011100",
			2196 => "0000000001000000001101011100010000",
			2197 => "0000000010000000001111100100001000",
			2198 => "0000000000000000000011010000000100",
			2199 => "00000000000000000010001010001001",
			2200 => "11111110101101100010001010001001",
			2201 => "0000001001000000001010011000000100",
			2202 => "11111111100000110010001010001001",
			2203 => "00000000100010000010001010001001",
			2204 => "0000000010000000001011111000001000",
			2205 => "0000000011000000001101000100000100",
			2206 => "00000000100101010010001010001001",
			2207 => "11111111101000000010001010001001",
			2208 => "00000001011001100010001010001001",
			2209 => "11111110101000110010001010001001",
			2210 => "0000000010000000000110111100001100",
			2211 => "0000000010000000000111011000000100",
			2212 => "11111110011001010010001100011101",
			2213 => "0000000010000000000110111100000100",
			2214 => "11111111101111110010001100011101",
			2215 => "11111110110100000010001100011101",
			2216 => "0000001100000000000100001000110000",
			2217 => "0000001001000000001011111100000100",
			2218 => "11111110100000100010001100011101",
			2219 => "0000001110000000001001010100010000",
			2220 => "0000001110000000001011000000000100",
			2221 => "00000101111010110010001100011101",
			2222 => "0000001000000000001010101100001000",
			2223 => "0000000101000000000101100100000100",
			2224 => "00000001110011010010001100011101",
			2225 => "00000000111101110010001100011101",
			2226 => "11111110110000010010001100011101",
			2227 => "0000001000000000001011010100001100",
			2228 => "0000001110000000001110101000001000",
			2229 => "0000001100000000001110001100000100",
			2230 => "00000000110011100010001100011101",
			2231 => "00000010101100010010001100011101",
			2232 => "11111110111011100010001100011101",
			2233 => "0000000010000000001000100000001000",
			2234 => "0000000101000000001010011100000100",
			2235 => "11111111101011010010001100011101",
			2236 => "11111100100000110010001100011101",
			2237 => "0000001111000000001111010100000100",
			2238 => "00000000101010110010001100011101",
			2239 => "11111111000111010010001100011101",
			2240 => "0000000111000000000111001000001100",
			2241 => "0000001011000000001000000000000100",
			2242 => "11111110101111010010001100011101",
			2243 => "0000000011000000000111100000000100",
			2244 => "00000001010000010010001100011101",
			2245 => "00000000000000000010001100011101",
			2246 => "11111110011000000010001100011101",
			2247 => "0000000010000000001111010100000100",
			2248 => "11111110011001100010001110101011",
			2249 => "0000001100000000000100001000110100",
			2250 => "0000000001000000001101101000000100",
			2251 => "11111110011101110010001110101011",
			2252 => "0000001110000000001001010100011000",
			2253 => "0000000001000000001111001100001100",
			2254 => "0000001000000000001000101100001000",
			2255 => "0000001011000000000111001000000100",
			2256 => "00000101010011010010001110101011",
			2257 => "00000011001001000010001110101011",
			2258 => "11111111011100000010001110101011",
			2259 => "0000000001000000001101011100001000",
			2260 => "0000001101000000000010001000000100",
			2261 => "00000001011110000010001110101011",
			2262 => "11111110110000010010001110101011",
			2263 => "00000001101101000010001110101011",
			2264 => "0000000001000000001001011000001100",
			2265 => "0000000100000000001101110100001000",
			2266 => "0000000100000000000000010100000100",
			2267 => "11111110111000110010001110101011",
			2268 => "00000000000000000010001110101011",
			2269 => "11111010001110100010001110101011",
			2270 => "0000001110000000001110101000001000",
			2271 => "0000000010000000000110101100000100",
			2272 => "00000000101110100010001110101011",
			2273 => "00000011101101110010001110101011",
			2274 => "11111110101101000010001110101011",
			2275 => "0000000111000000000111001000001100",
			2276 => "0000001110000000000111110000001000",
			2277 => "0000000101000000000100000100000100",
			2278 => "11111111011101110010001110101011",
			2279 => "00000001000011000010001110101011",
			2280 => "11111110010011000010001110101011",
			2281 => "11111110011001010010001110101011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(726, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(1470, initial_addr_3'length));
	end generate gen_rom_12;

	gen_rom_13: if SELECT_ROM = 13 generate
		bank <= (
			0 => "00000000000000000000000000000101",
			1 => "00000000000000000000000000001001",
			2 => "00000000000000000000000000001101",
			3 => "00000000000000000000000000010001",
			4 => "00000000000000000000000000010101",
			5 => "00000000000000000000000000011001",
			6 => "00000000000000000000000000011101",
			7 => "00000000000000000000000000100001",
			8 => "00000000000000000000000000100101",
			9 => "00000000000000000000000000101001",
			10 => "0000000100000000001110111000000100",
			11 => "11111111111000100000000000110101",
			12 => "00000000000000000000000000110101",
			13 => "0000000001000000001011101000000100",
			14 => "00000000000000000000000001001001",
			15 => "0000000001000000000000111100000100",
			16 => "00000000000010100000000001001001",
			17 => "00000000000000000000000001001001",
			18 => "0000001100000000000110000100001000",
			19 => "0000001100000000000000101000000100",
			20 => "00000000000000000000000001011101",
			21 => "00000000000111100000000001011101",
			22 => "00000000000000000000000001011101",
			23 => "0000001001000000001101101000000100",
			24 => "00000000000000000000000001110001",
			25 => "0000001001000000000100111100000100",
			26 => "00000000000100000000000001110001",
			27 => "00000000000000000000000001110001",
			28 => "0000000011000000000111100000001000",
			29 => "0000000100000000001101000000000100",
			30 => "11111111110001100000000010000101",
			31 => "00000000000000000000000010000101",
			32 => "00000000000000000000000010000101",
			33 => "0000001111000000000110010000001000",
			34 => "0000001111000000000010001000000100",
			35 => "00000000000000000000000010100001",
			36 => "00000000001001110000000010100001",
			37 => "0000001111000000001011110000000100",
			38 => "11111111110110010000000010100001",
			39 => "00000000000000000000000010100001",
			40 => "0000000110000000001011001100001000",
			41 => "0000000000000000000010111100000100",
			42 => "00000000000000000000000010111101",
			43 => "11111111110111110000000010111101",
			44 => "0000000110000000001000010000000100",
			45 => "00000000000010010000000010111101",
			46 => "00000000000000000000000010111101",
			47 => "0000000010000000000100101000000100",
			48 => "00000000000000000000000011011001",
			49 => "0000000100000000000001100100001000",
			50 => "0000001111000000001011110000000100",
			51 => "11111111011010100000000011011001",
			52 => "00000000000000000000000011011001",
			53 => "00000000000000000000000011011001",
			54 => "0000000101000000001011011100001100",
			55 => "0000000000000000000010111100000100",
			56 => "00000000000000000000000011110101",
			57 => "0000000000000000001010111100000100",
			58 => "11111111110101110000000011110101",
			59 => "00000000000000000000000011110101",
			60 => "00000000000000000000000011110101",
			61 => "0000001101000000001011110100001100",
			62 => "0000000000000000000010111100000100",
			63 => "00000000000000000000000100010001",
			64 => "0000000000000000001010111100000100",
			65 => "11111111101111110000000100010001",
			66 => "00000000000000000000000100010001",
			67 => "00000000000000000000000100010001",
			68 => "0000000000000000001110111100000100",
			69 => "00000000000000000000000100101101",
			70 => "0000000001000000001100110100000100",
			71 => "00000000000000000000000100101101",
			72 => "0000000001000000001101011100000100",
			73 => "00000000001011110000000100101101",
			74 => "00000000000000000000000100101101",
			75 => "0000000011000000000010001000001000",
			76 => "0000000110000000001001100100000100",
			77 => "11111111111000010000000101010001",
			78 => "00000000000000000000000101010001",
			79 => "0000001001000000000100111100001000",
			80 => "0000001001000000000001000100000100",
			81 => "00000000000000000000000101010001",
			82 => "00000000000100110000000101010001",
			83 => "00000000000000000000000101010001",
			84 => "0000000110000000001011001100001000",
			85 => "0000000010000000000100101000000100",
			86 => "00000000000000000000000101111101",
			87 => "11111111110000000000000101111101",
			88 => "0000000100000000001100111100001000",
			89 => "0000000100000000001000000100000100",
			90 => "00000000000000000000000101111101",
			91 => "11111111111101000000000101111101",
			92 => "0000000100000000000100100100000100",
			93 => "00000000001001010000000101111101",
			94 => "00000000000000000000000101111101",
			95 => "0000001100000000000011011100001100",
			96 => "0000000111000000001001110000000100",
			97 => "00000000000000000000000110101001",
			98 => "0000001101000000000100011000000100",
			99 => "00000000000000000000000110101001",
			100 => "00000000000100100000000110101001",
			101 => "0000001101000000001001010100001000",
			102 => "0000000111000000000110000100000100",
			103 => "00000000000000000000000110101001",
			104 => "11111111110110000000000110101001",
			105 => "00000000000000000000000110101001",
			106 => "0000000111000000001100101000010000",
			107 => "0000000111000000001001110000000100",
			108 => "00000000000000000000000111001101",
			109 => "0000001100000000001100110000001000",
			110 => "0000001100000000000000101000000100",
			111 => "00000000000000000000000111001101",
			112 => "00000000001100110000000111001101",
			113 => "00000000000000000000000111001101",
			114 => "11111111111110000000000111001101",
			115 => "0000000101000000001011011100010000",
			116 => "0000000100000000001000000100000100",
			117 => "00000000000000000000000111110001",
			118 => "0000000100000000001010010000001000",
			119 => "0000000010000000000100101000000100",
			120 => "00000000000000000000000111110001",
			121 => "11111111101011000000000111110001",
			122 => "00000000000000000000000111110001",
			123 => "00000000000000000000000111110001",
			124 => "0000000101000000001011011100000100",
			125 => "00000000000000000000001000010101",
			126 => "0000001001000000000101010000001100",
			127 => "0000001001000000000001111000000100",
			128 => "00000000000000000000001000010101",
			129 => "0000001101000000000111111100000100",
			130 => "00000000001111000000001000010101",
			131 => "00000000000000000000001000010101",
			132 => "00000000000000000000001000010101",
			133 => "0000000000000000001110111100000100",
			134 => "00000000000000000000001000111001",
			135 => "0000000001000000001100110100000100",
			136 => "00000000000000000000001000111001",
			137 => "0000000001000000001101011100001000",
			138 => "0000001000000000001101010000000100",
			139 => "00000000001111000000001000111001",
			140 => "00000000000000000000001000111001",
			141 => "00000000000000000000001000111001",
			142 => "0000000010000000000100101000000100",
			143 => "00000000000000000000001001100101",
			144 => "0000001101000000001011110100001000",
			145 => "0000000000000000001010111100000100",
			146 => "11111111101010000000001001100101",
			147 => "00000000000000000000001001100101",
			148 => "0000000111000000000100011000000100",
			149 => "00000000000010110000001001100101",
			150 => "0000000111000000000111010000000100",
			151 => "11111111111001010000001001100101",
			152 => "00000000000000000000001001100101",
			153 => "0000000000000000001110111100001100",
			154 => "0000000000000000000010111100000100",
			155 => "00000000000000000000001010011001",
			156 => "0000000100000000000000100000000100",
			157 => "11111111110101100000001010011001",
			158 => "00000000000000000000001010011001",
			159 => "0000001000000000000001110100001100",
			160 => "0000000111000000001001110000000100",
			161 => "00000000000000000000001010011001",
			162 => "0000000111000000001101010100000100",
			163 => "00000000010000010000001010011001",
			164 => "00000000000000000000001010011001",
			165 => "00000000000000000000001010011001",
			166 => "0000000000000000000011111100001100",
			167 => "0000001010000000000110011000000100",
			168 => "00000000000000000000001011001101",
			169 => "0000001010000000000001010000000100",
			170 => "00000000000100010000001011001101",
			171 => "00000000000000000000001011001101",
			172 => "0000001111000000001000101000001100",
			173 => "0000001010000000000110011000000100",
			174 => "00000000000000000000001011001101",
			175 => "0000000000000000001010111100000100",
			176 => "11111111111000010000001011001101",
			177 => "00000000000000000000001011001101",
			178 => "00000000000000000000001011001101",
			179 => "0000001010000000000001010000001100",
			180 => "0000001010000000000110011000000100",
			181 => "00000000000000000000001100000001",
			182 => "0000001100000000001001110000000100",
			183 => "00000000000000000000001100000001",
			184 => "00000000010011010000001100000001",
			185 => "0000001011000000000110100100001100",
			186 => "0000001100000000001000111100000100",
			187 => "00000000000000000000001100000001",
			188 => "0000000100000000001010010000000100",
			189 => "11111111110000110000001100000001",
			190 => "00000000000000000000001100000001",
			191 => "00000000000000000000001100000001",
			192 => "0000000011000000000010001000001000",
			193 => "0000000110000000001001100100000100",
			194 => "11111111110110110000001100110101",
			195 => "00000000000000000000001100110101",
			196 => "0000000110000000000101010000010000",
			197 => "0000000001000000000101011100001100",
			198 => "0000001001000000000001000100000100",
			199 => "00000000000000000000001100110101",
			200 => "0000000110000000001011001100000100",
			201 => "00000000000000000000001100110101",
			202 => "00000000011010110000001100110101",
			203 => "00000000000000000000001100110101",
			204 => "00000000000000000000001100110101",
			205 => "0000000100000000000100001100001100",
			206 => "0000000100000000001000000100000100",
			207 => "00000000000000000000001101110001",
			208 => "0000000110000000001000010000000100",
			209 => "11111111101000100000001101110001",
			210 => "00000000000000000000001101110001",
			211 => "0000000110000000001111000000010000",
			212 => "0000000001000000001100110100000100",
			213 => "00000000000000000000001101110001",
			214 => "0000000001000000001101011100001000",
			215 => "0000000100000000000100111000000100",
			216 => "00000000010110110000001101110001",
			217 => "00000000000000000000001101110001",
			218 => "00000000000000000000001101110001",
			219 => "00000000000000000000001101110001",
			220 => "0000000101000000001011011100001100",
			221 => "0000000100000000001000000100000100",
			222 => "00000000000000000000001110101101",
			223 => "0000000100000000000101001100000100",
			224 => "11111111111010000000001110101101",
			225 => "00000000000000000000001110101101",
			226 => "0000001100000000001010111000010000",
			227 => "0000000001000000000101011100001100",
			228 => "0000001110000000000100010000000100",
			229 => "00000000000000000000001110101101",
			230 => "0000001010000000000110011000000100",
			231 => "00000000000000000000001110101101",
			232 => "00000000011100010000001110101101",
			233 => "00000000000000000000001110101101",
			234 => "00000000000000000000001110101101",
			235 => "0000000111000000000111001000011100",
			236 => "0000001011000000000100011000010000",
			237 => "0000000100000000001000000100000100",
			238 => "00000000000000000000001111111001",
			239 => "0000000100000000001101000000001000",
			240 => "0000000011000000001000000000000100",
			241 => "00000000000000000000001111111001",
			242 => "11111111100110100000001111111001",
			243 => "00000000000000000000001111111001",
			244 => "0000001101000000000100010000000100",
			245 => "00000000000000000000001111111001",
			246 => "0000000100000000001001000000000100",
			247 => "00000000000000000000001111111001",
			248 => "00000000010111100000001111111001",
			249 => "0000000011000000000011000000001000",
			250 => "0000001100000000000000001100000100",
			251 => "00000000000000000000001111111001",
			252 => "11111111100001100000001111111001",
			253 => "00000000000000000000001111111001",
			254 => "0000001111000000000000010000011100",
			255 => "0000001101000000000100010000001000",
			256 => "0000001110000000000010001000000100",
			257 => "11111111111101100000010000111101",
			258 => "00000000000000000000010000111101",
			259 => "0000001011000000000100011000000100",
			260 => "00000000000000000000010000111101",
			261 => "0000001100000000000100001000001100",
			262 => "0000000001000000000101011100001000",
			263 => "0000001110000000000011001000000100",
			264 => "00000000010101000000010000111101",
			265 => "00000000000000000000010000111101",
			266 => "00000000000000000000010000111101",
			267 => "00000000000000000000010000111101",
			268 => "0000000000000000000010011000000100",
			269 => "00000000000000000000010000111101",
			270 => "11111111100010010000010000111101",
			271 => "0000000000000000000010111100010100",
			272 => "0000000000000000000010011000000100",
			273 => "00000000000000000000010010001001",
			274 => "0000000101000000001000000000000100",
			275 => "00000000000000000000010010001001",
			276 => "0000001000000000001011010100001000",
			277 => "0000000100000000000010100100000100",
			278 => "00000000011000010000010010001001",
			279 => "00000000000000000000010010001001",
			280 => "00000000000000000000010010001001",
			281 => "0000001111000000001010010100000100",
			282 => "00000000000000000000010010001001",
			283 => "0000000100000000000001100100001100",
			284 => "0000000010000000001010001000000100",
			285 => "00000000000000000000010010001001",
			286 => "0000001110000000001010000100000100",
			287 => "11111111100010000000010010001001",
			288 => "00000000000000000000010010001001",
			289 => "00000000000000000000010010001001",
			290 => "0000001101000000001001010100011000",
			291 => "0000000010000000001010001000000100",
			292 => "00000000000000000000010010111101",
			293 => "0000000000000000001010111100010000",
			294 => "0000000001000000001001011000001100",
			295 => "0000000000000000001000111100001000",
			296 => "0000000011000000000111100000000100",
			297 => "11111111101000100000010010111101",
			298 => "00000000000000000000010010111101",
			299 => "00000000000000000000010010111101",
			300 => "00000000000000000000010010111101",
			301 => "00000000000000000000010010111101",
			302 => "00000000000000000000010010111101",
			303 => "0000000000000000000010111100011000",
			304 => "0000001000000000001001101000000100",
			305 => "00000000000000000000010100001001",
			306 => "0000001001000000001001111100010000",
			307 => "0000001101000000001001110100000100",
			308 => "00000000000000000000010100001001",
			309 => "0000001000000000001011010100001000",
			310 => "0000000100000000001000000100000100",
			311 => "00000000000000000000010100001001",
			312 => "00000000101010110000010100001001",
			313 => "00000000000000000000010100001001",
			314 => "00000000000000000000010100001001",
			315 => "0000001001000000001110010100001100",
			316 => "0000000100000000001010010000001000",
			317 => "0000001111000000000010110100000100",
			318 => "00000000000000000000010100001001",
			319 => "11111111011110100000010100001001",
			320 => "00000000000000000000010100001001",
			321 => "00000000000000000000010100001001",
			322 => "0000001001000000000100110100100000",
			323 => "0000000010000000001110010000010100",
			324 => "0000000011000000000011100000000100",
			325 => "00000000000000000000010101011101",
			326 => "0000001011000000001110001100001100",
			327 => "0000001011000000000101101100000100",
			328 => "00000000000000000000010101011101",
			329 => "0000000011000000001010011100000100",
			330 => "00000000001010100000010101011101",
			331 => "00000000000000000000010101011101",
			332 => "00000000000000000000010101011101",
			333 => "0000000100000000001010010000001000",
			334 => "0000001111000000000111110000000100",
			335 => "00000000000000000000010101011101",
			336 => "11111111011100000000010101011101",
			337 => "00000000000000000000010101011101",
			338 => "0000000001000000001001011000001000",
			339 => "0000001001000000001010011000000100",
			340 => "00000000000000000000010101011101",
			341 => "00000000001011100000010101011101",
			342 => "00000000000000000000010101011101",
			343 => "0000001100000000000011011100011000",
			344 => "0000001011000000000101101100000100",
			345 => "00000000000000000000010110110001",
			346 => "0000001000000000001001101000000100",
			347 => "00000000000000000000010110110001",
			348 => "0000000010000000000110010000001100",
			349 => "0000000111000000001001110000000100",
			350 => "00000000000000000000010110110001",
			351 => "0000001101000000000100011000000100",
			352 => "00000000000000000000010110110001",
			353 => "00000000011000000000010110110001",
			354 => "00000000000000000000010110110001",
			355 => "0000001111000000000101110000000100",
			356 => "00000000000000000000010110110001",
			357 => "0000000011000000000011000000001100",
			358 => "0000000010000000000110101100000100",
			359 => "00000000000000000000010110110001",
			360 => "0000000111000000001100101000000100",
			361 => "00000000000000000000010110110001",
			362 => "11111111101011010000010110110001",
			363 => "00000000000000000000010110110001",
			364 => "0000001100000000001100110000011100",
			365 => "0000001100000000000100000000000100",
			366 => "00000000000000000000010111111101",
			367 => "0000000000000000000010111100000100",
			368 => "00000000000000000000010111111101",
			369 => "0000001110000000000101101100000100",
			370 => "00000000000000000000010111111101",
			371 => "0000000110000000000100110100000100",
			372 => "00000000000000000000010111111101",
			373 => "0000000010000000000010010100001000",
			374 => "0000000011000000001001011100000100",
			375 => "00000000010111100000010111111101",
			376 => "00000000000000000000010111111101",
			377 => "00000000000000000000010111111101",
			378 => "0000000010000000000011000000001000",
			379 => "0000000010000000000110101100000100",
			380 => "00000000000000000000010111111101",
			381 => "11111111110010010000010111111101",
			382 => "00000000000000000000010111111101",
			383 => "0000001111000000000110010000011100",
			384 => "0000000111000000001001110000000100",
			385 => "00000000000000000000011001000001",
			386 => "0000001100000000001110001100010100",
			387 => "0000000010000000001011101100010000",
			388 => "0000000110000000001001100100001100",
			389 => "0000000110000000000100110100000100",
			390 => "00000000000000000000011001000001",
			391 => "0000001111000000001011011100000100",
			392 => "00000000000000000000011001000001",
			393 => "00000000011010000000011001000001",
			394 => "00000000000000000000011001000001",
			395 => "00000000000000000000011001000001",
			396 => "00000000000000000000011001000001",
			397 => "0000001100000000000011011100000100",
			398 => "00000000000000000000011001000001",
			399 => "11111111110010010000011001000001",
			400 => "0000001001000000000111101000001000",
			401 => "0000000000000000001010111100000100",
			402 => "11111111101111110000011010000101",
			403 => "00000000000000000000011010000101",
			404 => "0000000111000000000100011000011000",
			405 => "0000001101000000000101110100000100",
			406 => "00000000000000000000011010000101",
			407 => "0000001001000000000100111100010000",
			408 => "0000000001000000001011101000000100",
			409 => "00000000000000000000011010000101",
			410 => "0000001111000000000011001000000100",
			411 => "00000000000000000000011010000101",
			412 => "0000001010000000000110011000000100",
			413 => "00000000000000000000011010000101",
			414 => "00000000011011100000011010000101",
			415 => "00000000000000000000011010000101",
			416 => "00000000000000000000011010000101",
			417 => "0000001001000000000001000100001000",
			418 => "0000000100000000000011111000000100",
			419 => "11111111100111010000011011011001",
			420 => "00000000000000000000011011011001",
			421 => "0000000001000000001111001100011000",
			422 => "0000000110000000001011001100000100",
			423 => "00000000000000000000011011011001",
			424 => "0000000011000000001001011100010000",
			425 => "0000001100000000000011011100000100",
			426 => "00000000000000000000011011011001",
			427 => "0000000000000000000010111100000100",
			428 => "00000000000000000000011011011001",
			429 => "0000001000000000001111000100000100",
			430 => "00000000110111010000011011011001",
			431 => "00000000000000000000011011011001",
			432 => "00000000000000000000011011011001",
			433 => "0000001111000000000010000000000100",
			434 => "00000000000000000000011011011001",
			435 => "0000000110000000000100111100000100",
			436 => "11111111111000010000011011011001",
			437 => "00000000000000000000011011011001",
			438 => "0000001100000000001100110000011100",
			439 => "0000001101000000000100011000000100",
			440 => "00000000000000000000011100101101",
			441 => "0000001000000000001001101000000100",
			442 => "00000000000000000000011100101101",
			443 => "0000001111000000000110010000010000",
			444 => "0000000110000000001111000000001100",
			445 => "0000000000000000000010111100000100",
			446 => "00000000000000000000011100101101",
			447 => "0000001100000000000000101000000100",
			448 => "00000000000000000000011100101101",
			449 => "00000000011100010000011100101101",
			450 => "00000000000000000000011100101101",
			451 => "00000000000000000000011100101101",
			452 => "0000000010000000001011111000000100",
			453 => "00000000000000000000011100101101",
			454 => "0000000000000000000010111100000100",
			455 => "00000000000000000000011100101101",
			456 => "0000000000000000001010111100000100",
			457 => "11111111101111000000011100101101",
			458 => "00000000000000000000011100101101",
			459 => "0000001100000000000011011100011100",
			460 => "0000001100000000000100000000000100",
			461 => "00000000000000000000011110000001",
			462 => "0000001000000000001001101000000100",
			463 => "00000000000000000000011110000001",
			464 => "0000000010000000000110010000010000",
			465 => "0000001001000000001101101000000100",
			466 => "00000000000000000000011110000001",
			467 => "0000001101000000000100011000000100",
			468 => "00000000000000000000011110000001",
			469 => "0000000111000000001001110000000100",
			470 => "00000000000000000000011110000001",
			471 => "00000000011011000000011110000001",
			472 => "00000000000000000000011110000001",
			473 => "0000001111000000000101110000000100",
			474 => "00000000000000000000011110000001",
			475 => "0000000000000000000010111100000100",
			476 => "00000000000000000000011110000001",
			477 => "0000000111000000000110000100000100",
			478 => "00000000000000000000011110000001",
			479 => "11111111101101110000011110000001",
			480 => "0000001001000000001101101000000100",
			481 => "00000000000000000000011110111101",
			482 => "0000000001000000000101011100011000",
			483 => "0000001011000000000101101100000100",
			484 => "00000000000000000000011110111101",
			485 => "0000001000000000001001101000000100",
			486 => "00000000000000000000011110111101",
			487 => "0000000110000000001000010000001100",
			488 => "0000000111000000001110110000001000",
			489 => "0000000000000000000010011000000100",
			490 => "00000000000000000000011110111101",
			491 => "00000000010110110000011110111101",
			492 => "00000000000000000000011110111101",
			493 => "00000000000000000000011110111101",
			494 => "00000000000000000000011110111101",
			495 => "0000001110000000001100101100000100",
			496 => "00000000000000000000011111111001",
			497 => "0000001100000000001110001100011000",
			498 => "0000001010000000000110011000000100",
			499 => "00000000000000000000011111111001",
			500 => "0000001001000000001101101000000100",
			501 => "00000000000000000000011111111001",
			502 => "0000001100000000000100000000000100",
			503 => "00000000000000000000011111111001",
			504 => "0000001001000000000100111100001000",
			505 => "0000001110000000001001011100000100",
			506 => "00000000010010000000011111111001",
			507 => "00000000000000000000011111111001",
			508 => "00000000000000000000011111111001",
			509 => "00000000000000000000011111111001",
			510 => "0000000101000000000000011100011000",
			511 => "0000000010000000001110010000010000",
			512 => "0000000011000000001010111100000100",
			513 => "00000000000000000000100001011101",
			514 => "0000000010000000000101001000000100",
			515 => "00000000000000000000100001011101",
			516 => "0000001111000000000010110100000100",
			517 => "00000000010110000000100001011101",
			518 => "00000000000000000000100001011101",
			519 => "0000000000000000001000111100000100",
			520 => "11111111001010110000100001011101",
			521 => "00000000000000000000100001011101",
			522 => "0000000001000000000000111100011000",
			523 => "0000001100000000001100110000000100",
			524 => "00000000000000000000100001011101",
			525 => "0000000010000000001100001100010000",
			526 => "0000000000000000001111000100000100",
			527 => "00000000000000000000100001011101",
			528 => "0000001001000000001011111100000100",
			529 => "00000000000000000000100001011101",
			530 => "0000001101000000000010001000000100",
			531 => "00000000000000000000100001011101",
			532 => "00000000101001000000100001011101",
			533 => "00000000000000000000100001011101",
			534 => "00000000000000000000100001011101",
			535 => "0000000001000000001011101000011100",
			536 => "0000001111000000000100101000011000",
			537 => "0000001110000000001100101100000100",
			538 => "00000000000000000000100010111001",
			539 => "0000000111000000001001110000000100",
			540 => "00000000000000000000100010111001",
			541 => "0000001100000000000110000100001100",
			542 => "0000001011000000000101101100000100",
			543 => "00000000000000000000100010111001",
			544 => "0000001100000000000100000000000100",
			545 => "00000000000000000000100010111001",
			546 => "00000000010111010000100010111001",
			547 => "00000000000000000000100010111001",
			548 => "11111111101110100000100010111001",
			549 => "0000000001000000001101011100010000",
			550 => "0000000000000000000000110000000100",
			551 => "00000000000000000000100010111001",
			552 => "0000000111000000000001101000001000",
			553 => "0000001010000000001010110000000100",
			554 => "00000000000000000000100010111001",
			555 => "00000000100111100000100010111001",
			556 => "00000000000000000000100010111001",
			557 => "00000000000000000000100010111001",
			558 => "0000000010000000000110101100011100",
			559 => "0000001011000000000101101100000100",
			560 => "00000000000000000000100100010101",
			561 => "0000001100000000001110001100010100",
			562 => "0000000000000000000010111100000100",
			563 => "00000000000000000000100100010101",
			564 => "0000001000000000001001101000000100",
			565 => "00000000000000000000100100010101",
			566 => "0000001100000000000100000000000100",
			567 => "00000000000000000000100100010101",
			568 => "0000000111000000001001110000000100",
			569 => "00000000000000000000100100010101",
			570 => "00000000010101000000100100010101",
			571 => "00000000000000000000100100010101",
			572 => "0000000000000000000010111100000100",
			573 => "00000000000000000000100100010101",
			574 => "0000001100000000001100110000000100",
			575 => "00000000000000000000100100010101",
			576 => "0000000111000000000110000100000100",
			577 => "00000000000000000000100100010101",
			578 => "0000000000000000001010111100000100",
			579 => "11111111101101000000100100010101",
			580 => "00000000000000000000100100010101",
			581 => "0000000111000000001100101000101100",
			582 => "0000000001000000000110101000010100",
			583 => "0000000100000000000011101100000100",
			584 => "11111111100001100000100110001001",
			585 => "0000001110000000000000001100001100",
			586 => "0000000111000000001001110000000100",
			587 => "00000000000000000000100110001001",
			588 => "0000000011000000001110001100000100",
			589 => "00000000000000000000100110001001",
			590 => "00000000010110010000100110001001",
			591 => "00000000000000000000100110001001",
			592 => "0000000110000000001000010000010100",
			593 => "0000000110000000001101011000000100",
			594 => "00000000000000000000100110001001",
			595 => "0000001100000000000011011100000100",
			596 => "00000000000000000000100110001001",
			597 => "0000000000000000000010111100000100",
			598 => "00000000000000000000100110001001",
			599 => "0000001010000000000110011000000100",
			600 => "00000000000000000000100110001001",
			601 => "00000000110011100000100110001001",
			602 => "00000000000000000000100110001001",
			603 => "0000000011000000000111100000001100",
			604 => "0000001011000000001110110000000100",
			605 => "00000000000000000000100110001001",
			606 => "0000000010000000000000010000000100",
			607 => "00000000000000000000100110001001",
			608 => "11111111011111010000100110001001",
			609 => "00000000000000000000100110001001",
			610 => "0000000100000000000011010100011000",
			611 => "0000001111000000000000110100010000",
			612 => "0000001110000000001101111000000100",
			613 => "00000000000000000000101000011101",
			614 => "0000001011000000000101101100000100",
			615 => "00000000000000000000101000011101",
			616 => "0000001011000000001100101100000100",
			617 => "00000000010001100000101000011101",
			618 => "00000000000000000000101000011101",
			619 => "0000000101000000000101110000000100",
			620 => "11111111001011000000101000011101",
			621 => "00000000000000000000101000011101",
			622 => "0000001000000000000111000100010100",
			623 => "0000001001000000000100111100010000",
			624 => "0000001010000000000110011000000100",
			625 => "00000000000000000000101000011101",
			626 => "0000000000000000000111111000001000",
			627 => "0000000001000000001100110100000100",
			628 => "00000000000000000000101000011101",
			629 => "00000000110100100000101000011101",
			630 => "00000000000000000000101000011101",
			631 => "00000000000000000000101000011101",
			632 => "0000000110000000000100111100011000",
			633 => "0000001101000000000001011000001100",
			634 => "0000000100000000000101001100001000",
			635 => "0000000011000000001110110000000100",
			636 => "00000000000000000000101000011101",
			637 => "11111111110000000000101000011101",
			638 => "00000000000000000000101000011101",
			639 => "0000000100000000000110110000000100",
			640 => "00000000000000000000101000011101",
			641 => "0000000001000000000110101000000100",
			642 => "00000000000000000000101000011101",
			643 => "00000000011010000000101000011101",
			644 => "0000001101000000001100100100000100",
			645 => "11111111100101110000101000011101",
			646 => "00000000000000000000101000011101",
			647 => "0000001101000000000100011000000100",
			648 => "11111111110011010000101001111001",
			649 => "0000000111000000001100101000011000",
			650 => "0000000000000000000010111100000100",
			651 => "00000000000000000000101001111001",
			652 => "0000000011000000001001011100010000",
			653 => "0000001001000000001101101000000100",
			654 => "00000000000000000000101001111001",
			655 => "0000001011000000000101101100000100",
			656 => "00000000000000000000101001111001",
			657 => "0000001100000000001110001100000100",
			658 => "00000000101100000000101001111001",
			659 => "00000000000000000000101001111001",
			660 => "00000000000000000000101001111001",
			661 => "0000000010000000000110101100000100",
			662 => "00000000000000000000101001111001",
			663 => "0000000001000000001111001100000100",
			664 => "00000000000000000000101001111001",
			665 => "0000000000000000000010111100000100",
			666 => "00000000000000000000101001111001",
			667 => "0000000000000000001000111000000100",
			668 => "11111111100100010000101001111001",
			669 => "00000000000000000000101001111001",
			670 => "0000001101000000001011000000001000",
			671 => "0000000100000000001101000000000100",
			672 => "11111110111110010000101011110101",
			673 => "00000000000000000000101011110101",
			674 => "0000000010000000000110010000010100",
			675 => "0000000111000000001101100000010000",
			676 => "0000001100000000001000111000000100",
			677 => "00000000000000000000101011110101",
			678 => "0000001011000000001110001100001000",
			679 => "0000000000000000000010111100000100",
			680 => "00000000000000000000101011110101",
			681 => "00000001011100010000101011110101",
			682 => "00000000000000000000101011110101",
			683 => "00000000000000000000101011110101",
			684 => "0000000001000000001011101000010000",
			685 => "0000000100000000000011111000001000",
			686 => "0000001110000000000011100000000100",
			687 => "00000000000000000000101011110101",
			688 => "11111111001010010000101011110101",
			689 => "0000000110000000001011001100000100",
			690 => "00000000000000000000101011110101",
			691 => "00000000010000000000101011110101",
			692 => "0000001010000000000110011000000100",
			693 => "11111111110000010000101011110101",
			694 => "0000000011000000001111101000001100",
			695 => "0000001011000000001110110000000100",
			696 => "00000000000000000000101011110101",
			697 => "0000000001000000000101011100000100",
			698 => "00000000110101010000101011110101",
			699 => "00000000000000000000101011110101",
			700 => "00000000000000000000101011110101",
			701 => "0000001101000000000100011000000100",
			702 => "11111110011010100000101101010001",
			703 => "0000001100000000000100001000011100",
			704 => "0000001010000000000111000100011000",
			705 => "0000000000000000000010011000000100",
			706 => "11111110101000110000101101010001",
			707 => "0000000010000000001001011100000100",
			708 => "00000100100000110000101101010001",
			709 => "0000000101000000000011100000001000",
			710 => "0000000011000000000011100000000100",
			711 => "00000000011101000000101101010001",
			712 => "11111110100110100000101101010001",
			713 => "0000000110000000001101011000000100",
			714 => "11111111101101110000101101010001",
			715 => "00000001000111110000101101010001",
			716 => "11111110100010110000101101010001",
			717 => "0000000010000000000101000000000100",
			718 => "11111110011001010000101101010001",
			719 => "0000001111000000000101000000001000",
			720 => "0000000100000000000011101100000100",
			721 => "00000001011101000000101101010001",
			722 => "11111111011110000000101101010001",
			723 => "11111110100000110000101101010001",
			724 => "0000000100000000001001000000100100",
			725 => "0000000100000000000011010100001100",
			726 => "0000000010000000000101000000000100",
			727 => "11111110011011010000101111110101",
			728 => "0000000010000000000101000000000100",
			729 => "00000000111011100000101111110101",
			730 => "11111110011100000000101111110101",
			731 => "0000001000000000000110001000010100",
			732 => "0000001000000000001001101000001100",
			733 => "0000000100000000000011110100001000",
			734 => "0000000100000000001111100000000100",
			735 => "00000000000000000000101111110101",
			736 => "00000001011100110000101111110101",
			737 => "11111110110100000000101111110101",
			738 => "0000001010000000001010110000000100",
			739 => "00000100011001110000101111110101",
			740 => "11111111011100000000101111110101",
			741 => "11111110011010000000101111110101",
			742 => "0000000001000000000010001100001100",
			743 => "0000000010000000001000101000001000",
			744 => "0000000010000000000001011100000100",
			745 => "11111110011010100000101111110101",
			746 => "11111100101000100000101111110101",
			747 => "00000000010100010000101111110101",
			748 => "0000000010000000001011110000011000",
			749 => "0000000010000000001110110100000100",
			750 => "00000101000010100000101111110101",
			751 => "0000001110000000001001010100001100",
			752 => "0000000001000000001101011100001000",
			753 => "0000000101000000000100011000000100",
			754 => "11111110010100100000101111110101",
			755 => "00000001101011100000101111110101",
			756 => "11111110100101010000101111110101",
			757 => "0000000001000000001001011000000100",
			758 => "00000110000111000000101111110101",
			759 => "00000001000101000000101111110101",
			760 => "0000001000000000000001110100001000",
			761 => "0000001010000000000110011100000100",
			762 => "11111111011010100000101111110101",
			763 => "00000000101101110000101111110101",
			764 => "11111110011000100000101111110101",
			765 => "0000001111000000000110010000110100",
			766 => "0000000111000000001001110000001000",
			767 => "0000001010000000000110001000000100",
			768 => "11111111011001110000110001101001",
			769 => "00000000000000000000110001101001",
			770 => "0000000111000000001101100000010100",
			771 => "0000000010000000000110010000010000",
			772 => "0000001110000000001001110000000100",
			773 => "00000000000000000000110001101001",
			774 => "0000001010000000000110011000000100",
			775 => "00000000000000000000110001101001",
			776 => "0000001101000000000100011000000100",
			777 => "00000000000000000000110001101001",
			778 => "00000001000000100000110001101001",
			779 => "00000000000000000000110001101001",
			780 => "0000000100000000001011001000001000",
			781 => "0000000010000000001010001000000100",
			782 => "00000000000000000000110001101001",
			783 => "11111111101001110000110001101001",
			784 => "0000001110000000001010111000000100",
			785 => "00000000000000000000110001101001",
			786 => "0000000111000000000111001000001000",
			787 => "0000001000000000001011010100000100",
			788 => "00000000000000000000110001101001",
			789 => "00000000100101100000110001101001",
			790 => "00000000000000000000110001101001",
			791 => "0000001110000000000111111100000100",
			792 => "11111111001101100000110001101001",
			793 => "00000000000000000000110001101001",
			794 => "0000000100000000001001000000011000",
			795 => "0000000100000000000100001100000100",
			796 => "11111110011100010000110011011101",
			797 => "0000001000000000000111000100010000",
			798 => "0000000100000000000100001100000100",
			799 => "00000110011110010000110011011101",
			800 => "0000000011000000001001011100000100",
			801 => "11111110101010100000110011011101",
			802 => "0000000111000000000111010000000100",
			803 => "00000010011000010000110011011101",
			804 => "11111110111111110000110011011101",
			805 => "11111110011010110000110011011101",
			806 => "0000000001000000001100110100000100",
			807 => "11111110011010000000110011011101",
			808 => "0000000110000000001000010000011100",
			809 => "0000000010000000000110010000000100",
			810 => "00000100111000110000110011011101",
			811 => "0000000110000000001101011000001000",
			812 => "0000001111000000001100100100000100",
			813 => "00000001011011100000110011011101",
			814 => "11111100101001110000110011011101",
			815 => "0000001101000000001011000000001000",
			816 => "0000000011000000001010111000000100",
			817 => "00000000000000000000110011011101",
			818 => "11111110010111010000110011011101",
			819 => "0000001000000000001011010100000100",
			820 => "11111111101110000000110011011101",
			821 => "00000001101110000000110011011101",
			822 => "11111110010111010000110011011101",
			823 => "0000000010000000000100101000010000",
			824 => "0000001110000000001001110000000100",
			825 => "00000000000000000000110101111001",
			826 => "0000000100000000000010111000000100",
			827 => "00000000000000000000110101111001",
			828 => "0000001011000000001101100000000100",
			829 => "00000000000000000000110101111001",
			830 => "00000000111001100000110101111001",
			831 => "0000000000000000000010111100011000",
			832 => "0000001010000000000110011000000100",
			833 => "00000000000000000000110101111001",
			834 => "0000000001000000000101011100010000",
			835 => "0000001001000000000001000100000100",
			836 => "00000000000000000000110101111001",
			837 => "0000001000000000001011010100001000",
			838 => "0000000100000000001011110000000100",
			839 => "00000000000000000000110101111001",
			840 => "00000000100111100000110101111001",
			841 => "00000000000000000000110101111001",
			842 => "00000000000000000000110101111001",
			843 => "0000000100000000001101110100001100",
			844 => "0000001001000000001111000000001000",
			845 => "0000000010000000000111111100000100",
			846 => "00000000000000000000110101111001",
			847 => "11111111000101110000110101111001",
			848 => "00000000000000000000110101111001",
			849 => "0000000110000000001111000000010000",
			850 => "0000001110000000001011000100000100",
			851 => "00000000000000000000110101111001",
			852 => "0000001011000000001110110000001000",
			853 => "0000000110000000001111000000000100",
			854 => "00000000010110110000110101111001",
			855 => "00000000000000000000110101111001",
			856 => "00000000000000000000110101111001",
			857 => "0000001110000000001001100000001000",
			858 => "0000000011000000000110100000000100",
			859 => "00000000000000000000110101111001",
			860 => "11111111011010000000110101111001",
			861 => "00000000000000000000110101111001",
			862 => "0000000100000000001001000000011100",
			863 => "0000000100000000000000010100000100",
			864 => "11111110011100000000110111101101",
			865 => "0000001011000000000101101100000100",
			866 => "11111110011011000000110111101101",
			867 => "0000001010000000001010110000010000",
			868 => "0000000001000000000101011100001100",
			869 => "0000001010000000000110011000001000",
			870 => "0000000100000000000011110100000100",
			871 => "00000000100011100000110111101101",
			872 => "11111111101001110000110111101101",
			873 => "00000010101010010000110111101101",
			874 => "11111110111010110000110111101101",
			875 => "11111110101011010000110111101101",
			876 => "0000000001000000001100110100000100",
			877 => "11111110011010100000110111101101",
			878 => "0000000110000000001000010000011000",
			879 => "0000000111000000000011100000010100",
			880 => "0000001001000000001101101000000100",
			881 => "00001000100011110000110111101101",
			882 => "0000000101000000000100011000001000",
			883 => "0000000011000000000111001000000100",
			884 => "00000000000000000000110111101101",
			885 => "11111110100001000000110111101101",
			886 => "0000001000000000001011010100000100",
			887 => "11111111100110110000110111101101",
			888 => "00000001100001110000110111101101",
			889 => "11111101110110000000110111101101",
			890 => "11111110011000000000110111101101",
			891 => "0000000110000000001000010000110000",
			892 => "0000001101000000000100011000000100",
			893 => "11111111011110100000111001010001",
			894 => "0000000010000000000110010000010100",
			895 => "0000000101000000001001110100010000",
			896 => "0000001010000000000110011000000100",
			897 => "00000000000000000000111001010001",
			898 => "0000001110000000001001110000000100",
			899 => "00000000000000000000111001010001",
			900 => "0000000000000000000010111100000100",
			901 => "00000000000000000000111001010001",
			902 => "00000000111000000000111001010001",
			903 => "00000000000000000000111001010001",
			904 => "0000000100000000001011001000001000",
			905 => "0000001101000000000110100000000100",
			906 => "11111111011101010000111001010001",
			907 => "00000000000000000000111001010001",
			908 => "0000000001000000000110101000000100",
			909 => "00000000000000000000111001010001",
			910 => "0000001011000000001001110100001000",
			911 => "0000001011000000001010111100000100",
			912 => "00000000000000000000111001010001",
			913 => "00000000011101010000111001010001",
			914 => "00000000000000000000111001010001",
			915 => "11111111010100100000111001010001",
			916 => "0000000100000000001001000000100100",
			917 => "0000000100000000000000010100000100",
			918 => "11111110011001110000111011111101",
			919 => "0000000000000000000010111100001100",
			920 => "0000000001000000000101011100001000",
			921 => "0000001010000000000110011000000100",
			922 => "11111110111011110000111011111101",
			923 => "00001011010010110000111011111101",
			924 => "11111110100110010000111011111101",
			925 => "0000001011000000000101101100000100",
			926 => "11111110011000010000111011111101",
			927 => "0000000110000000001010011000000100",
			928 => "00000100101001100000111011111101",
			929 => "0000001010000000001010110000001000",
			930 => "0000000001000000001001011000000100",
			931 => "00000111101011110000111011111101",
			932 => "11111110110100110000111011111101",
			933 => "11111110011101100000111011111101",
			934 => "0000001001000000001011101000001000",
			935 => "0000000001000000000010001100000100",
			936 => "11111110011000010000111011111101",
			937 => "11111111101011000000111011111101",
			938 => "0000000110000000000100111100100000",
			939 => "0000001110000000000111110000010000",
			940 => "0000001001000000001010011000001100",
			941 => "0000000000000000000100010100000100",
			942 => "00000110100111010000111011111101",
			943 => "0000001111000000001100010100000100",
			944 => "00000010000000100000111011111101",
			945 => "00000100001000100000111011111101",
			946 => "11111110100101110000111011111101",
			947 => "0000000101000000001011011100001000",
			948 => "0000001100000000001110001100000100",
			949 => "00000010110110100000111011111101",
			950 => "00000000000000000000111011111101",
			951 => "0000000111000000001010111100000100",
			952 => "00100000100001100000111011111101",
			953 => "00001010000100110000111011111101",
			954 => "0000001010000000000101000100000100",
			955 => "00000000101110000000111011111101",
			956 => "0000001101000000001001110100000100",
			957 => "11111011111110110000111011111101",
			958 => "11111110010111110000111011111101",
			959 => "0000001001000000001101101000000100",
			960 => "11111111001000110000111101110001",
			961 => "0000001100000000000011011100011000",
			962 => "0000001011000000000101101100000100",
			963 => "00000000000000000000111101110001",
			964 => "0000000000000000000010111100000100",
			965 => "00000000000000000000111101110001",
			966 => "0000000110000000001000010000001100",
			967 => "0000001100000000000100000000000100",
			968 => "00000000000000000000111101110001",
			969 => "0000000111000000001001110000000100",
			970 => "00000000000000000000111101110001",
			971 => "00000001000010000000111101110001",
			972 => "00000000000000000000111101110001",
			973 => "0000000010000000000011110000011100",
			974 => "0000001011000000000100011000001100",
			975 => "0000000100000000001101000000001000",
			976 => "0000001110000000000000001100000100",
			977 => "00000000000000000000111101110001",
			978 => "11111111011101100000111101110001",
			979 => "00000000000000000000111101110001",
			980 => "0000000001000000000000111100001100",
			981 => "0000000001000000001011101000000100",
			982 => "00000000000000000000111101110001",
			983 => "0000000100000000000000010100000100",
			984 => "00000000000000000000111101110001",
			985 => "00000000110100100000111101110001",
			986 => "00000000000000000000111101110001",
			987 => "11111111001111010000111101110001",
			988 => "0000001101000000000100011000000100",
			989 => "11111110011011010000111111010101",
			990 => "0000001000000000001001101000000100",
			991 => "11111110011111110000111111010101",
			992 => "0000000010000000001110010000001000",
			993 => "0000001011000000001110001100000100",
			994 => "00000010101100110000111111010101",
			995 => "11111111010001110000111111010101",
			996 => "0000000110000000001000010000011000",
			997 => "0000001011000000001110001100001000",
			998 => "0000000011000000000100011000000100",
			999 => "00000000110100100000111111010101",
			1000 => "11111110100101010000111111010101",
			1001 => "0000000110000000001011001100001000",
			1002 => "0000000100000000000101100000000100",
			1003 => "00000000100010110000111111010101",
			1004 => "11111110101101010000111111010101",
			1005 => "0000000001000000001001011000000100",
			1006 => "00000001001011110000111111010101",
			1007 => "11111111111011110000111111010101",
			1008 => "0000001010000000000001010000001000",
			1009 => "0000000001000000001110010100000100",
			1010 => "00000000110001000000111111010101",
			1011 => "11111111101101010000111111010101",
			1012 => "11111110100000010000111111010101",
			1013 => "0000001101000000000100011000000100",
			1014 => "11111110100111000001000001011001",
			1015 => "0000001111000000001101000100010000",
			1016 => "0000001111000000001011011100000100",
			1017 => "00000000000000000001000001011001",
			1018 => "0000000100000000000010111000000100",
			1019 => "00000000000000000001000001011001",
			1020 => "0000001100000000000110000100000100",
			1021 => "00000001011100100001000001011001",
			1022 => "00000000000000000001000001011001",
			1023 => "0000001001000000000100110100010100",
			1024 => "0000000100000000001101000000001000",
			1025 => "0000001100000000000110000100000100",
			1026 => "11111110100110100001000001011001",
			1027 => "00000000000000000001000001011001",
			1028 => "0000001100000000000110000100000100",
			1029 => "00000000100101010001000001011001",
			1030 => "0000000100000000000100111000000100",
			1031 => "00000000000000000001000001011001",
			1032 => "11111110110011010001000001011001",
			1033 => "0000000100000000000011010100000100",
			1034 => "11111111000111000001000001011001",
			1035 => "0000001010000000000110011100010000",
			1036 => "0000001110000000000100010000001000",
			1037 => "0000001001000000001010011000000100",
			1038 => "00000000000000000001000001011001",
			1039 => "11111111110110010001000001011001",
			1040 => "0000000111000000001010111100000100",
			1041 => "00000001010110010001000001011001",
			1042 => "00000000000110010001000001011001",
			1043 => "0000001101000000001001010100000100",
			1044 => "00000000000000000001000001011001",
			1045 => "11111111111100110001000001011001",
			1046 => "0000001010000000000110011000000100",
			1047 => "11111111000101100001000011001101",
			1048 => "0000001000000000001011010100010000",
			1049 => "0000000001000000000101011100001100",
			1050 => "0000001100000000000011011100000100",
			1051 => "00000000000000000001000011001101",
			1052 => "0000000100000000000111011100000100",
			1053 => "00000001010111000001000011001101",
			1054 => "00000000000000000001000011001101",
			1055 => "00000000000000000001000011001101",
			1056 => "0000000100000000000100001100000100",
			1057 => "11111111000110010001000011001101",
			1058 => "0000000010000000001110010000001000",
			1059 => "0000000011000000001010111100000100",
			1060 => "00000000000000000001000011001101",
			1061 => "00000001001011110001000011001101",
			1062 => "0000000001000000000110101000001100",
			1063 => "0000001000000000000010111100001000",
			1064 => "0000001111000000000111110000000100",
			1065 => "00000000000000000001000011001101",
			1066 => "11111111010011110001000011001101",
			1067 => "00000000000000000001000011001101",
			1068 => "0000000110000000001011001100001000",
			1069 => "0000001011000000001010111100000100",
			1070 => "00000000000000000001000011001101",
			1071 => "00000000100101100001000011001101",
			1072 => "0000000100000000001101000000000100",
			1073 => "11111111110001000001000011001101",
			1074 => "00000000000000000001000011001101",
			1075 => "0000000100000000001001000000101100",
			1076 => "0000001011000000000101101100000100",
			1077 => "11111110011001110001000101110001",
			1078 => "0000001101000000000110100100010100",
			1079 => "0000000101000000001000000000001000",
			1080 => "0000000001000000000010001100000100",
			1081 => "00000010110001000001000101110001",
			1082 => "11111110100011000001000101110001",
			1083 => "0000000010000000000110010000001000",
			1084 => "0000000000000000000010111100000100",
			1085 => "11111111110100010001000101110001",
			1086 => "00001000101100010001000101110001",
			1087 => "11111111011000000001000101110001",
			1088 => "0000000100000000000000010100000100",
			1089 => "11111110011010100001000101110001",
			1090 => "0000000000000000000010011000001100",
			1091 => "0000001010000000000110011000000100",
			1092 => "11111111111110100001000101110001",
			1093 => "0000000001000000000111101000000100",
			1094 => "00000001111000010001000101110001",
			1095 => "00000000000000000001000101110001",
			1096 => "11111110101000110001000101110001",
			1097 => "0000000001000000001100110100000100",
			1098 => "11111110011011010001000101110001",
			1099 => "0000000111000000000111001000011100",
			1100 => "0000001111000000000111110000000100",
			1101 => "00000011010101110001000101110001",
			1102 => "0000001011000000001110001100001000",
			1103 => "0000000000000000000100001000000100",
			1104 => "11111110011011110001000101110001",
			1105 => "00000001001110000001000101110001",
			1106 => "0000001100000000001100110000001000",
			1107 => "0000000000000000000100010100000100",
			1108 => "00000100101000010001000101110001",
			1109 => "00000001100101100001000101110001",
			1110 => "0000000110000000001101011000000100",
			1111 => "11111101110100110001000101110001",
			1112 => "00000001001010110001000101110001",
			1113 => "0000001100000000000100001000000100",
			1114 => "00000000000000000001000101110001",
			1115 => "11111110010101100001000101110001",
			1116 => "0000001001000000001111001100000100",
			1117 => "11111110100010010001000111110101",
			1118 => "0000001010000000000110011100100000",
			1119 => "0000000000000000001111000100000100",
			1120 => "11111110110100010001000111110101",
			1121 => "0000001100000000001000111000000100",
			1122 => "11111111000111010001000111110101",
			1123 => "0000001100000000000011011100001100",
			1124 => "0000001010000000000001010000000100",
			1125 => "00000001111010110001000111110101",
			1126 => "0000000000000000001010000000000100",
			1127 => "11111111110001000001000111110101",
			1128 => "00000001000110010001000111110101",
			1129 => "0000001101000000000010001000000100",
			1130 => "11111111001110000001000111110101",
			1131 => "0000001001000000000101010000000100",
			1132 => "00000000110111110001000111110101",
			1133 => "11111111111010000001000111110101",
			1134 => "0000000000000000001100101100011000",
			1135 => "0000001100000000001110001100010000",
			1136 => "0000001100000000001100110000001100",
			1137 => "0000000111000000000101101100000100",
			1138 => "11111111101000110001000111110101",
			1139 => "0000001111000000001100010000000100",
			1140 => "00000000001100100001000111110101",
			1141 => "00000000000000000001000111110101",
			1142 => "11111110011101110001000111110101",
			1143 => "0000001100000000000100001000000100",
			1144 => "00000000011111110001000111110101",
			1145 => "11111111101111100001000111110101",
			1146 => "0000000011000000001010110100000100",
			1147 => "00000000111001110001000111110101",
			1148 => "00000000000000000001000111110101",
			1149 => "0000001010000000000110011000000100",
			1150 => "11111111000001000001001001110001",
			1151 => "0000001000000000001011010100010000",
			1152 => "0000000001000000000101011100001100",
			1153 => "0000001100000000000011011100000100",
			1154 => "00000000000000000001001001110001",
			1155 => "0000000100000000000111011100000100",
			1156 => "00000001011110100001001001110001",
			1157 => "00000000000000000001001001110001",
			1158 => "00000000000000000001001001110001",
			1159 => "0000000100000000000100001100000100",
			1160 => "11111111000010100001001001110001",
			1161 => "0000000010000000001110010000001000",
			1162 => "0000000011000000001010111100000100",
			1163 => "00000000000000000001001001110001",
			1164 => "00000001010011010001001001110001",
			1165 => "0000000110000000001011001100010000",
			1166 => "0000001110000000000100011000001000",
			1167 => "0000001100000000001100110000000100",
			1168 => "00000000000000000001001001110001",
			1169 => "11111111110000110001001001110001",
			1170 => "0000001011000000001010111100000100",
			1171 => "00000000000000000001001001110001",
			1172 => "00000000101000110001001001110001",
			1173 => "0000000100000000001101000000001000",
			1174 => "0000000100000000000011101100000100",
			1175 => "00000000000000000001001001110001",
			1176 => "11111111001010110001001001110001",
			1177 => "0000001010000000001111001000000100",
			1178 => "00000000000111010001001001110001",
			1179 => "00000000000000000001001001110001",
			1180 => "0000001011000000000101101100000100",
			1181 => "11111110011110010001001011100101",
			1182 => "0000000100000000000010111000000100",
			1183 => "11111110101000000001001011100101",
			1184 => "0000001000000000000111000100010100",
			1185 => "0000000001000000000101011100010000",
			1186 => "0000000010000000000011001000000100",
			1187 => "00000001111010010001001011100101",
			1188 => "0000000101000000000101100100000100",
			1189 => "11111111000111100001001011100101",
			1190 => "0000001010000000000110011000000100",
			1191 => "00000000000000000001001011100101",
			1192 => "00000001001100110001001011100101",
			1193 => "11111111011010110001001011100101",
			1194 => "0000001100000000000110000100010000",
			1195 => "0000000100000000000001100100000100",
			1196 => "11111110110111110001001011100101",
			1197 => "0000000010000000000010010100001000",
			1198 => "0000001100000000001100110000000100",
			1199 => "00000001010110100001001011100101",
			1200 => "00000000000000000001001011100101",
			1201 => "11111111100100000001001011100101",
			1202 => "0000000110000000001011001100000100",
			1203 => "11111110001010100001001011100101",
			1204 => "0000000100000000000110110000000100",
			1205 => "11111111001111010001001011100101",
			1206 => "0000001100000000000100001000000100",
			1207 => "00000000110110010001001011100101",
			1208 => "11111111100011100001001011100101",
			1209 => "0000001101000000000100011000000100",
			1210 => "11111110111101110001001110000001",
			1211 => "0000000110000000001100011000010000",
			1212 => "0000001101000000000110100100001100",
			1213 => "0000000100000000000010111000000100",
			1214 => "00000000000000000001001110000001",
			1215 => "0000001111000000000001011000000100",
			1216 => "00000000000000000001001110000001",
			1217 => "00000001000001000001001110000001",
			1218 => "00000000000000000001001110000001",
			1219 => "0000000101000000000000011100010100",
			1220 => "0000000100000000001101000000001000",
			1221 => "0000001111000000001110101100000100",
			1222 => "00000000000000000001001110000001",
			1223 => "11111110111001000001001110000001",
			1224 => "0000001100000000000110000100001000",
			1225 => "0000001110000000000000101000000100",
			1226 => "00000000000000000001001110000001",
			1227 => "00000000001101000001001110000001",
			1228 => "00000000000000000001001110000001",
			1229 => "0000000111000000000001111100010000",
			1230 => "0000000001000000001111001100000100",
			1231 => "00000000000000000001001110000001",
			1232 => "0000001000000000001011010100000100",
			1233 => "00000000000000000001001110000001",
			1234 => "0000000011000000000110010000000100",
			1235 => "00000000111011110001001110000001",
			1236 => "00000000000000000001001110000001",
			1237 => "0000000001000000001001011000001100",
			1238 => "0000000110000000001001100100000100",
			1239 => "00000000000000000001001110000001",
			1240 => "0000001010000000001100000100000100",
			1241 => "00000000100010010001001110000001",
			1242 => "00000000000000000001001110000001",
			1243 => "0000001111000000001110100100001000",
			1244 => "0000000110000000001011001100000100",
			1245 => "00000000000000000001001110000001",
			1246 => "11111111010101100001001110000001",
			1247 => "00000000000000000001001110000001",
			1248 => "0000000111000000001001110000001000",
			1249 => "0000000010000000001000100000000100",
			1250 => "11111110101100010001010000100101",
			1251 => "00000000000000000001010000100101",
			1252 => "0000000111000000001001110000001100",
			1253 => "0000000010000000000110010000001000",
			1254 => "0000001101000000000100011000000100",
			1255 => "00000000000000000001010000100101",
			1256 => "00000001100100000001010000100101",
			1257 => "00000000000000000001010000100101",
			1258 => "0000001000000000000111000100010100",
			1259 => "0000000100000000000010111000000100",
			1260 => "11111111000100010001010000100101",
			1261 => "0000000001000000000101011100001100",
			1262 => "0000000001000000001001111000000100",
			1263 => "00000000000000000001010000100101",
			1264 => "0000001101000000001011000000000100",
			1265 => "00000000000000000001010000100101",
			1266 => "00000000110010110001010000100101",
			1267 => "00000000000000000001010000100101",
			1268 => "0000001111000000000101110000010100",
			1269 => "0000000110000000001101011000001100",
			1270 => "0000000100000000000100111000000100",
			1271 => "00000000000000000001010000100101",
			1272 => "0000000101000000001000000000000100",
			1273 => "00000000000000000001010000100101",
			1274 => "11111111100101100001010000100101",
			1275 => "0000000010000000001111010100000100",
			1276 => "00000000000000000001010000100101",
			1277 => "00000000101010010001010000100101",
			1278 => "0000000001000000001011101000001000",
			1279 => "0000000011000000000100000100000100",
			1280 => "00000000000000000001010000100101",
			1281 => "11111110111000010001010000100101",
			1282 => "0000000001000000001111001100001000",
			1283 => "0000000010000000001011110000000100",
			1284 => "00000000011011000001010000100101",
			1285 => "00000000000000000001010000100101",
			1286 => "0000000001000000001111001100000100",
			1287 => "11111111001110110001010000100101",
			1288 => "00000000000000000001010000100101",
			1289 => "0000000100000000001001000000110000",
			1290 => "0000001011000000000101101100000100",
			1291 => "11111110011010000001010011100001",
			1292 => "0000001101000000000110100100011000",
			1293 => "0000001101000000001001110100001000",
			1294 => "0000001001000000001011101000000100",
			1295 => "00000010000000010001010011100001",
			1296 => "11111110100101000001010011100001",
			1297 => "0000001100000000001000111000000100",
			1298 => "11111111001100000001010011100001",
			1299 => "0000001011000000001110001100001000",
			1300 => "0000000110000000001011001100000100",
			1301 => "00000110100110010001010011100001",
			1302 => "00000000000000000001010011100001",
			1303 => "00000000000000000001010011100001",
			1304 => "0000000100000000000000010100000100",
			1305 => "11111110011010110001010011100001",
			1306 => "0000000000000000000010011000001100",
			1307 => "0000001010000000000110011000000100",
			1308 => "00000000000000000001010011100001",
			1309 => "0000001001000000000100101100000100",
			1310 => "00000001110000010001010011100001",
			1311 => "00000000000000000001010011100001",
			1312 => "11111110101011000001010011100001",
			1313 => "0000000001000000001100110100000100",
			1314 => "11111110011011110001010011100001",
			1315 => "0000000111000000000111001000100000",
			1316 => "0000000110000000001010011000000100",
			1317 => "00000011010100100001010011100001",
			1318 => "0000001011000000001110001100001100",
			1319 => "0000000011000000001000000000001000",
			1320 => "0000001101000000000100011000000100",
			1321 => "11111111010110000001010011100001",
			1322 => "00000001010101110001010011100001",
			1323 => "11111110100000100001010011100001",
			1324 => "0000001100000000001100110000001000",
			1325 => "0000000000000000000100010100000100",
			1326 => "00000011110111010001010011100001",
			1327 => "00000001100011100001010011100001",
			1328 => "0000000110000000001101011000000100",
			1329 => "11111110000111110001010011100001",
			1330 => "00000001000101110001010011100001",
			1331 => "0000001010000000000001110000001000",
			1332 => "0000000100000000000110110000000100",
			1333 => "11111110111100010001010011100001",
			1334 => "00000000100110000001010011100001",
			1335 => "11111110010001100001010011100001",
			1336 => "0000001101000000000100011000000100",
			1337 => "11111110100011000001010110011101",
			1338 => "0000000010000000000110010000100100",
			1339 => "0000000111000000001101100000010000",
			1340 => "0000000000000000000010111100000100",
			1341 => "00000000000000000001010110011101",
			1342 => "0000001010000000001010110000001000",
			1343 => "0000000111000000001001110000000100",
			1344 => "00000000000000000001010110011101",
			1345 => "00000010010000000001010110011101",
			1346 => "00000000000000000001010110011101",
			1347 => "0000000100000000000011010100000100",
			1348 => "11111111011111000001010110011101",
			1349 => "0000000101000000000011100000000100",
			1350 => "00000000000000000001010110011101",
			1351 => "0000000101000000001001110100001000",
			1352 => "0000000111000000001101111000000100",
			1353 => "00000000101011100001010110011101",
			1354 => "00000000000000000001010110011101",
			1355 => "00000000000000000001010110011101",
			1356 => "0000001111000000000110010000100000",
			1357 => "0000000110000000001011001100001100",
			1358 => "0000000010000000001100111000001000",
			1359 => "0000001111000000001101000100000100",
			1360 => "00000000000000000001010110011101",
			1361 => "11111111000101010001010110011101",
			1362 => "00000000000000000001010110011101",
			1363 => "0000000100000000001101110100001000",
			1364 => "0000000100000000000001101100000100",
			1365 => "11111111100100000001010110011101",
			1366 => "00000000000000000001010110011101",
			1367 => "0000001011000000001000000000001000",
			1368 => "0000001011000000000110000100000100",
			1369 => "00000000000000000001010110011101",
			1370 => "00000001010100010001010110011101",
			1371 => "00000000000000000001010110011101",
			1372 => "0000001101000000001110101100001000",
			1373 => "0000001111000000001001100000000100",
			1374 => "00000000000000000001010110011101",
			1375 => "11111110100001100001010110011101",
			1376 => "0000000001000000000101011100001100",
			1377 => "0000000010000000000010110000001000",
			1378 => "0000001000000000001001101000000100",
			1379 => "00000000000000000001010110011101",
			1380 => "00000001000110100001010110011101",
			1381 => "11111111101101010001010110011101",
			1382 => "11111111001001100001010110011101",
			1383 => "0000001101000000000100011000000100",
			1384 => "11111110011011000001011000111001",
			1385 => "0000001100000000000100001000111100",
			1386 => "0000001110000000001010111000011100",
			1387 => "0000001111000000001011011100000100",
			1388 => "11111110110111100001011000111001",
			1389 => "0000000110000000001100011000001000",
			1390 => "0000001011000000001100101100000100",
			1391 => "00000011011110000001011000111001",
			1392 => "00000000000000000001011000111001",
			1393 => "0000000100000000000001100100001000",
			1394 => "0000000011000000001000000000000100",
			1395 => "00000000000000000001011000111001",
			1396 => "11111111011111110001011000111001",
			1397 => "0000000111000000001101100000000100",
			1398 => "00000000000000000001011000111001",
			1399 => "00000001100110100001011000111001",
			1400 => "0000000001000000000110101000000100",
			1401 => "11111110100000010001011000111001",
			1402 => "0000000101000000000000011100010000",
			1403 => "0000001001000000001011111100001000",
			1404 => "0000001100000000001001110000000100",
			1405 => "11111111010011000001011000111001",
			1406 => "00000001101101010001011000111001",
			1407 => "0000001101000000000001011000000100",
			1408 => "11111110100001010001011000111001",
			1409 => "00000000000000000001011000111001",
			1410 => "0000001001000000000100111100001000",
			1411 => "0000000110000000001000010000000100",
			1412 => "00000001011011110001011000111001",
			1413 => "11111111010001010001011000111001",
			1414 => "11111111000100010001011000111001",
			1415 => "0000000110000000001000010000000100",
			1416 => "11111110011111010001011000111001",
			1417 => "0000001111000000000101000000001000",
			1418 => "0000000001000000001011111100000100",
			1419 => "00000001001110100001011000111001",
			1420 => "11111111000011100001011000111001",
			1421 => "11111110101001000001011000111001",
			1422 => "0000000100000000001110111000000100",
			1423 => "11111110100001000001011011110101",
			1424 => "0000001000000000000111000100111000",
			1425 => "0000001000000000000111000100100000",
			1426 => "0000001000000000000110001000011000",
			1427 => "0000000100000000000011101100001100",
			1428 => "0000001110000000001101101100001000",
			1429 => "0000001010000000000110011000000100",
			1430 => "00000000000000000001011011110101",
			1431 => "00000001001100010001011011110101",
			1432 => "00000000000000000001011011110101",
			1433 => "0000001000000000001011010100001000",
			1434 => "0000000111000000001101010100000100",
			1435 => "11111111010110110001011011110101",
			1436 => "00000000000000000001011011110101",
			1437 => "00000000000000000001011011110101",
			1438 => "0000000100000000000000101100000100",
			1439 => "11111111011101110001011011110101",
			1440 => "00000000000000000001011011110101",
			1441 => "0000001111000000000101110100001000",
			1442 => "0000001011000000001100001000000100",
			1443 => "00000000000000000001011011110101",
			1444 => "00000100111100010001011011110101",
			1445 => "0000000100000000000100001100000100",
			1446 => "00000000000000000001011011110101",
			1447 => "0000000001000000001101011100001000",
			1448 => "0000000101000000000111001000000100",
			1449 => "00000000000000000001011011110101",
			1450 => "00000001011111000001011011110101",
			1451 => "00000000000000000001011011110101",
			1452 => "0000000110000000000100111100011100",
			1453 => "0000000100000000000001100100000100",
			1454 => "11111110101101010001011011110101",
			1455 => "0000001100000000001100110000001000",
			1456 => "0000001011000000001110001100000100",
			1457 => "00000000000000000001011011110101",
			1458 => "00000001000101010001011011110101",
			1459 => "0000000110000000001001100100001000",
			1460 => "0000000100000000000011111000000100",
			1461 => "00000000000000000001011011110101",
			1462 => "11111110111010000001011011110101",
			1463 => "0000000001000000001101011100000100",
			1464 => "00000000100100000001011011110101",
			1465 => "00000000000000000001011011110101",
			1466 => "0000001001000000001001100100000100",
			1467 => "11111110011011110001011011110101",
			1468 => "00000000000000000001011011110101",
			1469 => "0000001101000000000100011000000100",
			1470 => "11111110011100110001011111001011",
			1471 => "0000001100000000000011011100011100",
			1472 => "0000001110000000000100001000001100",
			1473 => "0000000100000000001110111000000100",
			1474 => "00000000000000000001011111001011",
			1475 => "0000000110000000001111000000000100",
			1476 => "00000001101111000001011111001011",
			1477 => "00000000000000000001011111001011",
			1478 => "0000001100000000000011011100001000",
			1479 => "0000000100000000001101000000000100",
			1480 => "11111110101001000001011111001011",
			1481 => "00000000001010000001011111001011",
			1482 => "0000000011000000000101110100000100",
			1483 => "00000000000000000001011111001011",
			1484 => "00000001111001100001011111001011",
			1485 => "0000000110000000001011001100011100",
			1486 => "0000001100000000001100110000001000",
			1487 => "0000000000000000001100001000000100",
			1488 => "00000000000000000001011111001011",
			1489 => "00000000001010110001011111001011",
			1490 => "0000001011000000000000001100001100",
			1491 => "0000001011000000000000001100000100",
			1492 => "11111111100110100001011111001011",
			1493 => "0000001101000000000001101000000100",
			1494 => "00000000000000000001011111001011",
			1495 => "11111010101101000001011111001011",
			1496 => "0000000111000000001110001100000100",
			1497 => "00000000000000000001011111001011",
			1498 => "11111110010000110001011111001011",
			1499 => "0000000110000000001111000000011100",
			1500 => "0000000100000000001101110100001100",
			1501 => "0000001101000000001001010100000100",
			1502 => "11111110111101110001011111001011",
			1503 => "0000001100000000000100001000000100",
			1504 => "00000000110110010001011111001011",
			1505 => "11111111011110000001011111001011",
			1506 => "0000000000000000000100010100001000",
			1507 => "0000000010000000000110101100000100",
			1508 => "00000001011000010001011111001011",
			1509 => "11111111010110110001011111001011",
			1510 => "0000000011000000001101010100000100",
			1511 => "00000000000000000001011111001011",
			1512 => "00000001011101010001011111001011",
			1513 => "0000000010000000001000011100001000",
			1514 => "0000000011000000000010110100000100",
			1515 => "00000000000000000001011111001011",
			1516 => "11111110011101110001011111001011",
			1517 => "0000000011000000001111101000001000",
			1518 => "0000001010000000000101000100000100",
			1519 => "00000001000111110001011111001011",
			1520 => "00000000000000000001011111001011",
			1521 => "11111110111010000001011111001011",
			1522 => "00000000000000000001011111001101",
			1523 => "00000000000000000001011111010001",
			1524 => "00000000000000000001011111010101",
			1525 => "00000000000000000001011111011001",
			1526 => "00000000000000000001011111011101",
			1527 => "00000000000000000001011111100001",
			1528 => "00000000000000000001011111100101",
			1529 => "00000000000000000001011111101001",
			1530 => "00000000000000000001011111101101",
			1531 => "00000000000000000001011111110001",
			1532 => "0000000010000000000110010000000100",
			1533 => "00000000000000000001011111111101",
			1534 => "00000000000000000001011111111101",
			1535 => "0000000001000000001011101000000100",
			1536 => "11111111111111110001100000010001",
			1537 => "0000000001000000000000111100000100",
			1538 => "00000000000010000001100000010001",
			1539 => "00000000000000000001100000010001",
			1540 => "0000001100000000000110000100001000",
			1541 => "0000001100000000000000101000000100",
			1542 => "00000000000000000001100000100101",
			1543 => "00000000000111000001100000100101",
			1544 => "00000000000000000001100000100101",
			1545 => "0000000110000000001000010000001000",
			1546 => "0000000110000000000100110100000100",
			1547 => "00000000000000000001100000111001",
			1548 => "00000000000110000001100000111001",
			1549 => "00000000000000000001100000111001",
			1550 => "0000001110000000001110101100001000",
			1551 => "0000000100000000001101000000000100",
			1552 => "11111111110011100001100001001101",
			1553 => "00000000000000000001100001001101",
			1554 => "00000000000000000001100001001101",
			1555 => "0000001111000000000110010000001000",
			1556 => "0000001111000000000010001000000100",
			1557 => "00000000000000000001100001101001",
			1558 => "00000000001000100001100001101001",
			1559 => "0000001111000000001011110000000100",
			1560 => "11111111110111010001100001101001",
			1561 => "00000000000000000001100001101001",
			1562 => "0000001111000000000010000000001000",
			1563 => "0000001111000000000010001000000100",
			1564 => "00000000000000000001100010000101",
			1565 => "00000000000000100001100010000101",
			1566 => "0000001111000000001000110100000100",
			1567 => "11111111110111010001100010000101",
			1568 => "00000000000000000001100010000101",
			1569 => "0000000010000000000100101000000100",
			1570 => "00000000000000000001100010100001",
			1571 => "0000000100000000001101110100001000",
			1572 => "0000001110000000001010000100000100",
			1573 => "11111111011010110001100010100001",
			1574 => "00000000000000000001100010100001",
			1575 => "00000000000000000001100010100001",
			1576 => "0000000000000000001000111100001100",
			1577 => "0000000000000000000011111100000100",
			1578 => "00000000000000000001100010111101",
			1579 => "0000001111000000000101110100000100",
			1580 => "00000000000000000001100010111101",
			1581 => "11111111110010100001100010111101",
			1582 => "00000000000000000001100010111101",
			1583 => "0000001000000000000110001000000100",
			1584 => "00000000000000000001100011011001",
			1585 => "0000001100000000001000111100000100",
			1586 => "00000000000000000001100011011001",
			1587 => "0000000000000000000000111000000100",
			1588 => "00000000000000000001100011011001",
			1589 => "11111111110111000001100011011001",
			1590 => "0000001110000000001100101100000100",
			1591 => "00000000000000000001100011110101",
			1592 => "0000001010000000000110011000000100",
			1593 => "00000000000000000001100011110101",
			1594 => "0000001110000000001101101100000100",
			1595 => "00000000001001010001100011110101",
			1596 => "00000000000000000001100011110101",
			1597 => "0000001111000000000010000000001000",
			1598 => "0000001111000000000010001000000100",
			1599 => "00000000000000000001100100011001",
			1600 => "00000000000000110001100100011001",
			1601 => "0000001111000000001000110100001000",
			1602 => "0000001111000000000110010000000100",
			1603 => "00000000000000000001100100011001",
			1604 => "11111111110100010001100100011001",
			1605 => "00000000000000000001100100011001",
			1606 => "0000001100000000000011011100001100",
			1607 => "0000000111000000001001110000000100",
			1608 => "00000000000000000001100101000101",
			1609 => "0000001101000000000100011000000100",
			1610 => "00000000000000000001100101000101",
			1611 => "00000000000101000001100101000101",
			1612 => "0000001101000000001001010100001000",
			1613 => "0000000111000000000110000100000100",
			1614 => "00000000000000000001100101000101",
			1615 => "11111111110100000001100101000101",
			1616 => "00000000000000000001100101000101",
			1617 => "0000000100000000001100111100001100",
			1618 => "0000000010000000000100101000000100",
			1619 => "00000000000000000001100101110001",
			1620 => "0000000010000000001110100100000100",
			1621 => "11111111100001000001100101110001",
			1622 => "00000000000000000001100101110001",
			1623 => "0000001101000000000001011000000100",
			1624 => "00000000000000000001100101110001",
			1625 => "0000001101000000001001010000000100",
			1626 => "00000000001000000001100101110001",
			1627 => "00000000000000000001100101110001",
			1628 => "0000000111000000001100101000010000",
			1629 => "0000000111000000001001110000000100",
			1630 => "00000000000000000001100110010101",
			1631 => "0000001100000000001100110000001000",
			1632 => "0000001100000000000000101000000100",
			1633 => "00000000000000000001100110010101",
			1634 => "00000000001001110001100110010101",
			1635 => "00000000000000000001100110010101",
			1636 => "11111111111111110001100110010101",
			1637 => "0000001100000000001100110000010000",
			1638 => "0000000001000000001100110100000100",
			1639 => "00000000000000000001100110111001",
			1640 => "0000000001000000001111001100001000",
			1641 => "0000001100000000000000101000000100",
			1642 => "00000000000000000001100110111001",
			1643 => "00000000010010100001100110111001",
			1644 => "00000000000000000001100110111001",
			1645 => "11111111111111110001100110111001",
			1646 => "0000001110000000001100101100000100",
			1647 => "00000000000000000001100111011101",
			1648 => "0000001010000000000110011000000100",
			1649 => "00000000000000000001100111011101",
			1650 => "0000001110000000001101101100001000",
			1651 => "0000001010000000001100000100000100",
			1652 => "00000000001001000001100111011101",
			1653 => "00000000000000000001100111011101",
			1654 => "00000000000000000001100111011101",
			1655 => "0000001001000000001101101000000100",
			1656 => "00000000000000000001101000000001",
			1657 => "0000001001000000001101011000001100",
			1658 => "0000001011000000000101101100000100",
			1659 => "00000000000000000001101000000001",
			1660 => "0000001011000000001011110100000100",
			1661 => "00000000001000010001101000000001",
			1662 => "00000000000000000001101000000001",
			1663 => "00000000000000000001101000000001",
			1664 => "0000001100000000001100110000010000",
			1665 => "0000000111000000001001110000000100",
			1666 => "00000000000000000001101000110101",
			1667 => "0000000111000000001100101000001000",
			1668 => "0000001100000000000000101000000100",
			1669 => "00000000000000000001101000110101",
			1670 => "00000000001011010001101000110101",
			1671 => "00000000000000000001101000110101",
			1672 => "0000001010000000000001010000000100",
			1673 => "00000000000000000001101000110101",
			1674 => "0000001010000000001100000100000100",
			1675 => "11111111111000110001101000110101",
			1676 => "00000000000000000001101000110101",
			1677 => "0000000000000000000011111100001100",
			1678 => "0000001010000000000110011000000100",
			1679 => "00000000000000000001101001101001",
			1680 => "0000001010000000000001010000000100",
			1681 => "00000000000101110001101001101001",
			1682 => "00000000000000000001101001101001",
			1683 => "0000000100000000000001100100001100",
			1684 => "0000001111000000000101110100000100",
			1685 => "00000000000000000001101001101001",
			1686 => "0000001100000000000000001100000100",
			1687 => "11111111100110010001101001101001",
			1688 => "00000000000000000001101001101001",
			1689 => "00000000000000000001101001101001",
			1690 => "0000000100000000001100111100001100",
			1691 => "0000000010000000000100101000000100",
			1692 => "00000000000000000001101010011101",
			1693 => "0000001111000000001011110000000100",
			1694 => "11111111011110100001101010011101",
			1695 => "00000000000000000001101010011101",
			1696 => "0000000110000000001101011000000100",
			1697 => "00000000000000000001101010011101",
			1698 => "0000000110000000001000010000001000",
			1699 => "0000001101000000000101100100000100",
			1700 => "00000000000000000001101010011101",
			1701 => "00000000001111100001101010011101",
			1702 => "00000000000000000001101010011101",
			1703 => "0000000100000000000001100100010000",
			1704 => "0000001010000000000001010000000100",
			1705 => "00000000000000000001101011011001",
			1706 => "0000001111000000000101110100000100",
			1707 => "00000000000000000001101011011001",
			1708 => "0000000000000000000010011000000100",
			1709 => "00000000000000000001101011011001",
			1710 => "11111111100101100001101011011001",
			1711 => "0000000001000000001111001100001100",
			1712 => "0000000001000000000010001100000100",
			1713 => "00000000000000000001101011011001",
			1714 => "0000001111000000001000001100000100",
			1715 => "00000000001100010001101011011001",
			1716 => "00000000000000000001101011011001",
			1717 => "00000000000000000001101011011001",
			1718 => "0000001110000000000111110000001000",
			1719 => "0000000101000000000100010000000100",
			1720 => "11111111111100110001101100001101",
			1721 => "00000000000000000001101100001101",
			1722 => "0000000001000000000101011100010000",
			1723 => "0000000001000000001011101000000100",
			1724 => "00000000000000000001101100001101",
			1725 => "0000000101000000000101100100000100",
			1726 => "00000000000000000001101100001101",
			1727 => "0000000101000000000111111100000100",
			1728 => "00000000010101100001101100001101",
			1729 => "00000000000000000001101100001101",
			1730 => "00000000000000000001101100001101",
			1731 => "0000000110000000001101011000001000",
			1732 => "0000000100000000001110111000000100",
			1733 => "11111111110101110001101101001001",
			1734 => "00000000000000000001101101001001",
			1735 => "0000000110000000001001100100010000",
			1736 => "0000000001000000000111100100000100",
			1737 => "00000000000000000001101101001001",
			1738 => "0000000001000000000000111100001000",
			1739 => "0000000100000000001000000100000100",
			1740 => "00000000000000000001101101001001",
			1741 => "00000000010111100001101101001001",
			1742 => "00000000000000000001101101001001",
			1743 => "0000000100000000000011111000000100",
			1744 => "11111111111011000001101101001001",
			1745 => "00000000000000000001101101001001",
			1746 => "0000001001000000000100110100010000",
			1747 => "0000001111000000001110101000000100",
			1748 => "00000000000000000001101110001101",
			1749 => "0000000100000000001010010000001000",
			1750 => "0000000101000000000100010000000100",
			1751 => "11111111101101110001101110001101",
			1752 => "00000000000000000001101110001101",
			1753 => "00000000000000000001101110001101",
			1754 => "0000000001000000000000111100010000",
			1755 => "0000001001000000000100111100001100",
			1756 => "0000000001000000000000111100001000",
			1757 => "0000000001000000001011101000000100",
			1758 => "00000000000000000001101110001101",
			1759 => "00000000000010010001101110001101",
			1760 => "00000000000000000001101110001101",
			1761 => "00000000000000000001101110001101",
			1762 => "00000000000000000001101110001101",
			1763 => "0000000011000000000101110100001000",
			1764 => "0000000011000000000010001000000100",
			1765 => "11111111111011110001101111001001",
			1766 => "00000000000000000001101111001001",
			1767 => "0000000001000000000101011100010100",
			1768 => "0000000001000000001011101000000100",
			1769 => "00000000000000000001101111001001",
			1770 => "0000001110000000000100010000000100",
			1771 => "00000000000000000001101111001001",
			1772 => "0000000011000000001110101100000100",
			1773 => "00000000000000000001101111001001",
			1774 => "0000000011000000000010010100000100",
			1775 => "00000000010100100001101111001001",
			1776 => "00000000000000000001101111001001",
			1777 => "00000000000000000001101111001001",
			1778 => "0000000100000000000011101100001100",
			1779 => "0000000110000000001000010000001000",
			1780 => "0000001010000000001010110000000100",
			1781 => "11111111100010110001110000001101",
			1782 => "00000000000000000001110000001101",
			1783 => "00000000000000000001110000001101",
			1784 => "0000000110000000001000010000010100",
			1785 => "0000000111000000000100011000010000",
			1786 => "0000000110000000001101011000000100",
			1787 => "00000000000000000001110000001101",
			1788 => "0000001001000000001001011000000100",
			1789 => "00000000000000000001110000001101",
			1790 => "0000001010000000000110011000000100",
			1791 => "00000000000000000001110000001101",
			1792 => "00000000010100010001110000001101",
			1793 => "00000000000000000001110000001101",
			1794 => "00000000000000000001110000001101",
			1795 => "0000000000000000000010111100010100",
			1796 => "0000000000000000000010011000000100",
			1797 => "00000000000000000001110001100001",
			1798 => "0000000101000000001000000000000100",
			1799 => "00000000000000000001110001100001",
			1800 => "0000000001000000000101011100001000",
			1801 => "0000001000000000001011010100000100",
			1802 => "00000000011011010001110001100001",
			1803 => "00000000000000000001110001100001",
			1804 => "00000000000000000001110001100001",
			1805 => "0000001111000000001010010100001000",
			1806 => "0000001110000000001001110000000100",
			1807 => "00000000000000000001110001100001",
			1808 => "00000000000001100001110001100001",
			1809 => "0000000100000000000001100100001100",
			1810 => "0000000010000000001010001000000100",
			1811 => "00000000000000000001110001100001",
			1812 => "0000001110000000001010000100000100",
			1813 => "11111111011111110001110001100001",
			1814 => "00000000000000000001110001100001",
			1815 => "00000000000000000001110001100001",
			1816 => "0000001110000000001100101100000100",
			1817 => "00000000000000000001110010010101",
			1818 => "0000001010000000000110011000000100",
			1819 => "00000000000000000001110010010101",
			1820 => "0000000111000000000110100100010000",
			1821 => "0000001001000000001101101000000100",
			1822 => "00000000000000000001110010010101",
			1823 => "0000000001000000000101011100001000",
			1824 => "0000000111000000001001110000000100",
			1825 => "00000000000000000001110010010101",
			1826 => "00000000001110100001110010010101",
			1827 => "00000000000000000001110010010101",
			1828 => "00000000000000000001110010010101",
			1829 => "0000001100000000001100110000011000",
			1830 => "0000001101000000000100011000000100",
			1831 => "00000000000000000001110011100001",
			1832 => "0000001000000000001001101000000100",
			1833 => "00000000000000000001110011100001",
			1834 => "0000000010000000000110111000001100",
			1835 => "0000000000000000000010111100000100",
			1836 => "00000000000000000001110011100001",
			1837 => "0000000111000000001001110000000100",
			1838 => "00000000000000000001110011100001",
			1839 => "00000000011100000001110011100001",
			1840 => "00000000000000000001110011100001",
			1841 => "0000000010000000001011111000000100",
			1842 => "00000000000000000001110011100001",
			1843 => "0000000000000000000010111100000100",
			1844 => "00000000000000000001110011100001",
			1845 => "0000000000000000001010111100000100",
			1846 => "11111111101100110001110011100001",
			1847 => "00000000000000000001110011100001",
			1848 => "0000000000000000000010111100010100",
			1849 => "0000000000000000000010011000000100",
			1850 => "00000000000000000001110100111101",
			1851 => "0000000101000000001000000000000100",
			1852 => "00000000000000000001110100111101",
			1853 => "0000001000000000001011010100001000",
			1854 => "0000000100000000000010100100000100",
			1855 => "00000000011100100001110100111101",
			1856 => "00000000000000000001110100111101",
			1857 => "00000000000000000001110100111101",
			1858 => "0000001111000000001010010100001100",
			1859 => "0000001110000000001001110000000100",
			1860 => "00000000000000000001110100111101",
			1861 => "0000000011000000001010111100000100",
			1862 => "00000000000000000001110100111101",
			1863 => "00000000000100100001110100111101",
			1864 => "0000000000000000001010111100001100",
			1865 => "0000001110000000001001100000001000",
			1866 => "0000000010000000001010001000000100",
			1867 => "00000000000000000001110100111101",
			1868 => "11111111101001110001110100111101",
			1869 => "00000000000000000001110100111101",
			1870 => "00000000000000000001110100111101",
			1871 => "0000001001000000000001000100001000",
			1872 => "0000000100000000000011111000000100",
			1873 => "11111111101001000001110110001001",
			1874 => "00000000000000000001110110001001",
			1875 => "0000000001000000001111001100011000",
			1876 => "0000000110000000001011001100000100",
			1877 => "00000000000000000001110110001001",
			1878 => "0000000011000000001001011100010000",
			1879 => "0000000000000000000010111100000100",
			1880 => "00000000000000000001110110001001",
			1881 => "0000001011000000001110001100000100",
			1882 => "00000000000000000001110110001001",
			1883 => "0000000110000000001000010000000100",
			1884 => "00000000110001110001110110001001",
			1885 => "00000000000000000001110110001001",
			1886 => "00000000000000000001110110001001",
			1887 => "0000001111000000000010000000000100",
			1888 => "00000000000000000001110110001001",
			1889 => "11111111111110100001110110001001",
			1890 => "0000000100000000000011101100001100",
			1891 => "0000000110000000001000010000001000",
			1892 => "0000001010000000001010110000000100",
			1893 => "11111111100000000001110111010101",
			1894 => "00000000000000000001110111010101",
			1895 => "00000000000000000001110111010101",
			1896 => "0000000110000000001000010000011000",
			1897 => "0000000111000000000100011000010100",
			1898 => "0000000110000000001101011000000100",
			1899 => "00000000000000000001110111010101",
			1900 => "0000000001000000001001111000000100",
			1901 => "00000000000000000001110111010101",
			1902 => "0000001010000000000110011000000100",
			1903 => "00000000000000000001110111010101",
			1904 => "0000000111000000001101100000000100",
			1905 => "00000000000000000001110111010101",
			1906 => "00000000010111000001110111010101",
			1907 => "00000000000000000001110111010101",
			1908 => "00000000000000000001110111010101",
			1909 => "0000001111000000000110010000011100",
			1910 => "0000001100000000000000101000000100",
			1911 => "00000000000000000001111000011001",
			1912 => "0000001010000000001001000100000100",
			1913 => "00000000000000000001111000011001",
			1914 => "0000001111000000001011011100000100",
			1915 => "00000000000000000001111000011001",
			1916 => "0000000010000000001011101100001100",
			1917 => "0000001010000000000001110000001000",
			1918 => "0000001100000000001110001100000100",
			1919 => "00000000011000110001111000011001",
			1920 => "00000000000000000001111000011001",
			1921 => "00000000000000000001111000011001",
			1922 => "00000000000000000001111000011001",
			1923 => "0000001100000000000011011100000100",
			1924 => "00000000000000000001111000011001",
			1925 => "11111111110011110001111000011001",
			1926 => "0000000100000000000011010100011000",
			1927 => "0000000010000000000100101000010000",
			1928 => "0000001011000000000101101100000100",
			1929 => "00000000000000000001111010001101",
			1930 => "0000001011000000000110000100001000",
			1931 => "0000000110000000000100110100000100",
			1932 => "00000000000000000001111010001101",
			1933 => "00000000001111000001111010001101",
			1934 => "00000000000000000001111010001101",
			1935 => "0000000111000000000111010000000100",
			1936 => "11111111001001000001111010001101",
			1937 => "00000000000000000001111010001101",
			1938 => "0000001010000000000101000100010000",
			1939 => "0000000001000000000101011100001100",
			1940 => "0000001010000000000110011000000100",
			1941 => "00000000000000000001111010001101",
			1942 => "0000001101000000000100011000000100",
			1943 => "00000000000000000001111010001101",
			1944 => "00000000101010110001111010001101",
			1945 => "00000000000000000001111010001101",
			1946 => "0000001111000000000001000000000100",
			1947 => "00000000000000000001111010001101",
			1948 => "0000000010000000001011101100000100",
			1949 => "00000000000000000001111010001101",
			1950 => "0000000011000000001111011100000100",
			1951 => "00000000000000000001111010001101",
			1952 => "0000001101000000001011110100000100",
			1953 => "11111111010111100001111010001101",
			1954 => "00000000000000000001111010001101",
			1955 => "0000000110000000001011001100010000",
			1956 => "0000001001000000001001100100001100",
			1957 => "0000001111000000001010010100000100",
			1958 => "00000000000000000001111011100001",
			1959 => "0000001010000000001100000100000100",
			1960 => "11111111100100110001111011100001",
			1961 => "00000000000000000001111011100001",
			1962 => "00000000000000000001111011100001",
			1963 => "0000001001000000001101011000011000",
			1964 => "0000001001000000000001000100000100",
			1965 => "00000000000000000001111011100001",
			1966 => "0000000011000000001001011100010000",
			1967 => "0000001100000000000011011100000100",
			1968 => "00000000000000000001111011100001",
			1969 => "0000000100000000001000000100000100",
			1970 => "00000000000000000001111011100001",
			1971 => "0000001010000000001100000100000100",
			1972 => "00000000101111110001111011100001",
			1973 => "00000000000000000001111011100001",
			1974 => "00000000000000000001111011100001",
			1975 => "00000000000000000001111011100001",
			1976 => "0000001111000000000000010000100100",
			1977 => "0000000011000000000101110100001100",
			1978 => "0000000100000000001101000000001000",
			1979 => "0000001111000000001010010100000100",
			1980 => "00000000000000000001111100110101",
			1981 => "11111111110001110001111100110101",
			1982 => "00000000000000000001111100110101",
			1983 => "0000000001000000000111100100000100",
			1984 => "00000000000000000001111100110101",
			1985 => "0000001100000000000100001000010000",
			1986 => "0000000110000000001011001100000100",
			1987 => "00000000000000000001111100110101",
			1988 => "0000001100000000000011011100000100",
			1989 => "00000000000000000001111100110101",
			1990 => "0000000100000000001000000100000100",
			1991 => "00000000000000000001111100110101",
			1992 => "00000000010110010001111100110101",
			1993 => "00000000000000000001111100110101",
			1994 => "0000000000000000000010011000000100",
			1995 => "00000000000000000001111100110101",
			1996 => "11111111011110010001111100110101",
			1997 => "0000001101000000000100011000000100",
			1998 => "11111111110101100001111101110001",
			1999 => "0000000111000000001100101000011000",
			2000 => "0000000000000000000010111100000100",
			2001 => "00000000000000000001111101110001",
			2002 => "0000000011000000001001011100010000",
			2003 => "0000001000000000000111000100001100",
			2004 => "0000001100000000001110001100001000",
			2005 => "0000000111000000001001110000000100",
			2006 => "00000000000000000001111101110001",
			2007 => "00000000101010000001111101110001",
			2008 => "00000000000000000001111101110001",
			2009 => "00000000000000000001111101110001",
			2010 => "00000000000000000001111101110001",
			2011 => "00000000000000000001111101110001",
			2012 => "0000000001000000000110101000000100",
			2013 => "00000000000000000001111110101101",
			2014 => "0000000001000000000101011100011000",
			2015 => "0000001010000000001001000100000100",
			2016 => "00000000000000000001111110101101",
			2017 => "0000000111000000001001110000000100",
			2018 => "00000000000000000001111110101101",
			2019 => "0000001101000000001001110100000100",
			2020 => "00000000000000000001111110101101",
			2021 => "0000000110000000000101010000001000",
			2022 => "0000001100000000001000111000000100",
			2023 => "00000000000000000001111110101101",
			2024 => "00000000010100000001111110101101",
			2025 => "00000000000000000001111110101101",
			2026 => "00000000000000000001111110101101",
			2027 => "0000001110000000001100101100000100",
			2028 => "00000000000000000001111111101001",
			2029 => "0000000111000000001100101000011000",
			2030 => "0000001000000000001001101000000100",
			2031 => "00000000000000000001111111101001",
			2032 => "0000001001000000001101101000000100",
			2033 => "00000000000000000001111111101001",
			2034 => "0000000111000000001001110000000100",
			2035 => "00000000000000000001111111101001",
			2036 => "0000000110000000001000010000001000",
			2037 => "0000000100000000001000000100000100",
			2038 => "00000000000000000001111111101001",
			2039 => "00000000010111100001111111101001",
			2040 => "00000000000000000001111111101001",
			2041 => "00000000000000000001111111101001",
			2042 => "0000000001000000000110101000010100",
			2043 => "0000001111000000001010010100001100",
			2044 => "0000001110000000001001110000000100",
			2045 => "00000000000000000010000001011101",
			2046 => "0000000100000000001110111000000100",
			2047 => "00000000000000000010000001011101",
			2048 => "00000000011001010010000001011101",
			2049 => "0000001000000000000010111100000100",
			2050 => "11111111011100000010000001011101",
			2051 => "00000000000000000010000001011101",
			2052 => "0000000001000000001111001100011000",
			2053 => "0000000000000000000010111100000100",
			2054 => "00000000000000000010000001011101",
			2055 => "0000000111000000001001110000000100",
			2056 => "00000000000000000010000001011101",
			2057 => "0000000011000000001001011100001100",
			2058 => "0000000101000000001000000000000100",
			2059 => "00000000000000000010000001011101",
			2060 => "0000001100000000001000111000000100",
			2061 => "00000000000000000010000001011101",
			2062 => "00000000110100000010000001011101",
			2063 => "00000000000000000010000001011101",
			2064 => "0000000010000000000110101100000100",
			2065 => "00000000000000000010000001011101",
			2066 => "0000000111000000001101111000000100",
			2067 => "00000000000000000010000001011101",
			2068 => "0000000111000000000111010000000100",
			2069 => "11111111110000010010000001011101",
			2070 => "00000000000000000010000001011101",
			2071 => "0000000010000000000110101100011100",
			2072 => "0000001001000000001101101000000100",
			2073 => "00000000000000000010000010111001",
			2074 => "0000000000000000000010111100000100",
			2075 => "00000000000000000010000010111001",
			2076 => "0000001011000000000101101100000100",
			2077 => "00000000000000000010000010111001",
			2078 => "0000000110000000001001100100001100",
			2079 => "0000001000000000001001101000000100",
			2080 => "00000000000000000010000010111001",
			2081 => "0000000111000000001001110000000100",
			2082 => "00000000000000000010000010111001",
			2083 => "00000000011010100010000010111001",
			2084 => "00000000000000000010000010111001",
			2085 => "0000001100000000001100110000000100",
			2086 => "00000000000000000010000010111001",
			2087 => "0000001110000000001010000100001100",
			2088 => "0000000000000000000010111100000100",
			2089 => "00000000000000000010000010111001",
			2090 => "0000000000000000001010111100000100",
			2091 => "11111111011010110010000010111001",
			2092 => "00000000000000000010000010111001",
			2093 => "00000000000000000010000010111001",
			2094 => "0000000111000000001100101000100100",
			2095 => "0000001101000000000100011000000100",
			2096 => "11111111101001110010000100010101",
			2097 => "0000000110000000001000010000011100",
			2098 => "0000000100000000000011010100010000",
			2099 => "0000001000000000001011010100001100",
			2100 => "0000000111000000001101100000001000",
			2101 => "0000001000000000001001101000000100",
			2102 => "00000000000000000010000100010101",
			2103 => "00000000011000000010000100010101",
			2104 => "00000000000000000010000100010101",
			2105 => "11111111111111110010000100010101",
			2106 => "0000000001000000001100110100000100",
			2107 => "00000000000000000010000100010101",
			2108 => "0000001000000000001011010100000100",
			2109 => "00000000000000000010000100010101",
			2110 => "00000000101001000010000100010101",
			2111 => "00000000000000000010000100010101",
			2112 => "0000001101000000001001010100001000",
			2113 => "0000000010000000000000010000000100",
			2114 => "00000000000000000010000100010101",
			2115 => "11111111011110010010000100010101",
			2116 => "00000000000000000010000100010101",
			2117 => "0000001101000000000100011000000100",
			2118 => "11111110110011010010000101111001",
			2119 => "0000000111000000001100101000100100",
			2120 => "0000001000000000000111000100010000",
			2121 => "0000000000000000000010111100000100",
			2122 => "00000000000000000010000101111001",
			2123 => "0000000111000000001001110000000100",
			2124 => "00000000000000000010000101111001",
			2125 => "0000000110000000001000010000000100",
			2126 => "00000001011100000010000101111001",
			2127 => "00000000000000000010000101111001",
			2128 => "0000000100000000001101000000001000",
			2129 => "0000001011000000000000001100000100",
			2130 => "11111111010110110010000101111001",
			2131 => "00000000000000000010000101111001",
			2132 => "0000000110000000001101011000000100",
			2133 => "00000000000000000010000101111001",
			2134 => "0000000000000000000001001000000100",
			2135 => "00000000101011010010000101111001",
			2136 => "00000000000000000010000101111001",
			2137 => "0000000010000000001000100000001000",
			2138 => "0000001010000000000110011000000100",
			2139 => "11111111111111000010000101111001",
			2140 => "00000000000000000010000101111001",
			2141 => "11111111001001010010000101111001",
			2142 => "0000000111000000001001110000001000",
			2143 => "0000000010000000001000100000000100",
			2144 => "11111110011010110010000111011101",
			2145 => "00000000000000000010000111011101",
			2146 => "0000001100000000000100001000011100",
			2147 => "0000001010000000000111000100011000",
			2148 => "0000000000000000000010011000000100",
			2149 => "11111110101110100010000111011101",
			2150 => "0000000010000000000100101000000100",
			2151 => "00000011010101010010000111011101",
			2152 => "0000001011000000001100101100001000",
			2153 => "0000000100000000000010010000000100",
			2154 => "11111110101000010010000111011101",
			2155 => "00000000000101100010000111011101",
			2156 => "0000000110000000001000010000000100",
			2157 => "00000000111101110010000111011101",
			2158 => "11111110101111000010000111011101",
			2159 => "11111110101000000010000111011101",
			2160 => "0000000010000000000101000000000100",
			2161 => "11111110011011000010000111011101",
			2162 => "0000000011000000001111101000001000",
			2163 => "0000000011000000001101101100000100",
			2164 => "11111111110101000010000111011101",
			2165 => "00000001011011000010000111011101",
			2166 => "11111110100011100010000111011101",
			2167 => "0000000000000000000010111100011000",
			2168 => "0000001000000000001001101000000100",
			2169 => "11111111110111100010001001100001",
			2170 => "0000001100000000001000111000000100",
			2171 => "00000000000000000010001001100001",
			2172 => "0000000001000000000101011100001100",
			2173 => "0000001000000000001011010100001000",
			2174 => "0000000100000000001000000100000100",
			2175 => "00000000000000000010001001100001",
			2176 => "00000001001011110010001001100001",
			2177 => "00000000000000000010001001100001",
			2178 => "00000000000000000010001001100001",
			2179 => "0000000110000000001100011000010000",
			2180 => "0000000011000000000100011000000100",
			2181 => "11111111100111110010001001100001",
			2182 => "0000000001000000000010001100000100",
			2183 => "00000000000000000010001001100001",
			2184 => "0000000100000000000011001100000100",
			2185 => "00000000000000000010001001100001",
			2186 => "00000000110110010010001001100001",
			2187 => "0000000100000000001011001000000100",
			2188 => "11111111000111110010001001100001",
			2189 => "0000000110000000001111000000010000",
			2190 => "0000001110000000001001010100001100",
			2191 => "0000000001000000001111001100001000",
			2192 => "0000001001000000001001011000000100",
			2193 => "00000000000000000010001001100001",
			2194 => "00000000001001000010001001100001",
			2195 => "11111111110000100010001001100001",
			2196 => "00000000011010100010001001100001",
			2197 => "0000000100000000000101001100000100",
			2198 => "11111111010100010010001001100001",
			2199 => "00000000000000000010001001100001",
			2200 => "0000001111000000000110010000110100",
			2201 => "0000000111000000001001110000001000",
			2202 => "0000001010000000000110001000000100",
			2203 => "11111111011101110010001011011101",
			2204 => "00000000000000000010001011011101",
			2205 => "0000000111000000001101100000010100",
			2206 => "0000000010000000000110010000010000",
			2207 => "0000001110000000001001110000000100",
			2208 => "00000000000000000010001011011101",
			2209 => "0000000000000000000010111100000100",
			2210 => "00000000000000000010001011011101",
			2211 => "0000001000000000000111000100000100",
			2212 => "00000001000011000010001011011101",
			2213 => "00000000000000000010001011011101",
			2214 => "00000000000000000010001011011101",
			2215 => "0000001000000000001010101100001100",
			2216 => "0000001111000000000011001000001000",
			2217 => "0000000011000000001010111000000100",
			2218 => "00000000000000000010001011011101",
			2219 => "11111111011111110010001011011101",
			2220 => "00000000000000000010001011011101",
			2221 => "0000000110000000001101011000000100",
			2222 => "00000000000000000010001011011101",
			2223 => "0000000000000000000101100100000100",
			2224 => "00000000010110100010001011011101",
			2225 => "00000000000000000010001011011101",
			2226 => "0000001011000000000110100100000100",
			2227 => "11111111001010010010001011011101",
			2228 => "0000001100000000000100001000000100",
			2229 => "00000000000000110010001011011101",
			2230 => "00000000000000000010001011011101",
			2231 => "0000000100000000001110111000000100",
			2232 => "11111111001101000010001101000001",
			2233 => "0000001000000000000111000100011000",
			2234 => "0000000001000000000101011100010100",
			2235 => "0000000001000000001100110100000100",
			2236 => "00000000000000000010001101000001",
			2237 => "0000001010000000001100011100001100",
			2238 => "0000001010000000000110011000000100",
			2239 => "00000000000000000010001101000001",
			2240 => "0000001101000000000100011000000100",
			2241 => "00000000000000000010001101000001",
			2242 => "00000000011111010010001101000001",
			2243 => "00000000000000000010001101000001",
			2244 => "00000000000000000010001101000001",
			2245 => "0000000110000000000100111100010100",
			2246 => "0000000100000000000110110000001000",
			2247 => "0000000001000000001101011100000100",
			2248 => "11111111111101110010001101000001",
			2249 => "00000000000000000010001101000001",
			2250 => "0000000110000000001011001100000100",
			2251 => "00000000000000000010001101000001",
			2252 => "0000000001000000000010001100000100",
			2253 => "00000000000000000010001101000001",
			2254 => "00000000011101100010001101000001",
			2255 => "11111111100010100010001101000001",
			2256 => "0000000100000000001001000000100100",
			2257 => "0000000100000000000011010100001100",
			2258 => "0000000010000000000101000000000100",
			2259 => "11111110011100010010001111000101",
			2260 => "0000000010000000000101000000000100",
			2261 => "00000000110110100010001111000101",
			2262 => "11111110011101010010001111000101",
			2263 => "0000001000000000000110001000010100",
			2264 => "0000001010000000000110011000001100",
			2265 => "0000000100000000000011110100001000",
			2266 => "0000000110000000001101011000000100",
			2267 => "00000000000000000010001111000101",
			2268 => "00000001001101000010001111000101",
			2269 => "11111110111100010010001111000101",
			2270 => "0000001100000000001000011000000100",
			2271 => "00000011000011100010001111000101",
			2272 => "11111111100111010010001111000101",
			2273 => "11111110011010110010001111000101",
			2274 => "0000000011000000001110001100000100",
			2275 => "11111110011010000010001111000101",
			2276 => "0000000110000000001000010000011000",
			2277 => "0000001100000000000100001000010100",
			2278 => "0000000101000000000100011000000100",
			2279 => "11111110101001010010001111000101",
			2280 => "0000000010000000001011111000001000",
			2281 => "0000001010000000000110011000000100",
			2282 => "11111111000000110010001111000101",
			2283 => "00000010110101010010001111000101",
			2284 => "0000000100000000001100111100000100",
			2285 => "11111110011111110010001111000101",
			2286 => "00000001101000110010001111000101",
			2287 => "11111101100110010010001111000101",
			2288 => "11111110010111000010001111000101",
			2289 => "0000000100000000000001100100111000",
			2290 => "0000000100000000000011101100011100",
			2291 => "0000000100000000001110111000000100",
			2292 => "10111111100110110010010001110001",
			2293 => "0000001000000000001011010100001100",
			2294 => "0000000011000000000010010100001000",
			2295 => "0000001010000000000110011000000100",
			2296 => "10111111110010110010010001110001",
			2297 => "11100001010010100010010001110001",
			2298 => "10111111101011100010010001110001",
			2299 => "0000001011000000000101101100000100",
			2300 => "10111111100110010010010001110001",
			2301 => "0000001101000000000011100000000100",
			2302 => "11000011001110100010010001110001",
			2303 => "10111111101001110010010001110001",
			2304 => "0000000101000000001011011100001100",
			2305 => "0000000101000000000011100000000100",
			2306 => "10111111100110110010010001110001",
			2307 => "0000000011000000000111110000000100",
			2308 => "11001100011001010010010001110001",
			2309 => "10111111101001010010010001110001",
			2310 => "0000001010000000000001010000000100",
			2311 => "11011111001000010010010001110001",
			2312 => "0000001000000000000110001000001000",
			2313 => "0000000001000000001001011000000100",
			2314 => "11010010111101010010010001110001",
			2315 => "11000000011100100010010001110001",
			2316 => "10111111101111000010010001110001",
			2317 => "0000000001000000000010001100000100",
			2318 => "10111111100110000010010001110001",
			2319 => "0000001111000000001100010100001100",
			2320 => "0000000100000000001011100100001000",
			2321 => "0000001101000000001011011100000100",
			2322 => "11000000001110100010010001110001",
			2323 => "11111011000110110010010001110001",
			2324 => "00010000000000010010010001110001",
			2325 => "0000001100000000000100001000001100",
			2326 => "0000000100000000000110110000001000",
			2327 => "0000001011000000000011100000000100",
			2328 => "11000000001100100010010001110001",
			2329 => "11001100011001010010010001110001",
			2330 => "11110011000001100010010001110001",
			2331 => "10111111100110010010010001110001",
			2332 => "0000001101000000000100011000000100",
			2333 => "11111111100110110010010011100101",
			2334 => "0000000010000000001110010000001100",
			2335 => "0000000000000000000010111100000100",
			2336 => "00000000000000000010010011100101",
			2337 => "0000001100000000000011011100000100",
			2338 => "00000000110101010010010011100101",
			2339 => "00000000000000000010010011100101",
			2340 => "0000000001000000001011101000001100",
			2341 => "0000001110000000000000001100000100",
			2342 => "00000000000000000010010011100101",
			2343 => "0000000000000000001010111100000100",
			2344 => "11111111011000100010010011100101",
			2345 => "00000000000000000010010011100101",
			2346 => "0000000001000000001111001100001100",
			2347 => "0000001010000000001100011100000100",
			2348 => "00000000000000000010010011100101",
			2349 => "0000001111000000001111100100000100",
			2350 => "00000000100100000010010011100101",
			2351 => "00000000000000000010010011100101",
			2352 => "0000000010000000000110101100001100",
			2353 => "0000000101000000000101100100000100",
			2354 => "00000000000000000010010011100101",
			2355 => "0000001110000000001110101000000100",
			2356 => "00000000010011110010010011100101",
			2357 => "00000000000000000010010011100101",
			2358 => "0000000010000000001000011100000100",
			2359 => "11111111100101000010010011100101",
			2360 => "00000000000000000010010011100101",
			2361 => "0000000100000000000000010100000100",
			2362 => "11111110101001010010010101110001",
			2363 => "0000001000000000000111000100101000",
			2364 => "0000000000000000001110111100011000",
			2365 => "0000000010000000001011111000001100",
			2366 => "0000001010000000000110011000000100",
			2367 => "00000000000000000010010101110001",
			2368 => "0000001100000000001001110000000100",
			2369 => "00000000000000000010010101110001",
			2370 => "00000000011011110010010101110001",
			2371 => "0000001110000000001011111000000100",
			2372 => "11111111110001100010010101110001",
			2373 => "0000000010000000000011110000000100",
			2374 => "00000000000000010010010101110001",
			2375 => "00000000000000000010010101110001",
			2376 => "0000001000000000001111001000000100",
			2377 => "00000000000000000010010101110001",
			2378 => "0000000000000000000111111000001000",
			2379 => "0000000011000000001010111100000100",
			2380 => "00000000000000000010010101110001",
			2381 => "00000001111100100010010101110001",
			2382 => "00000000000000000010010101110001",
			2383 => "0000001111000000001001100000010100",
			2384 => "0000001001000000001001011000001000",
			2385 => "0000000010000000001011101100000100",
			2386 => "11111111000000000010010101110001",
			2387 => "00000000000000000010010101110001",
			2388 => "0000001001000000001010011000001000",
			2389 => "0000001011000000001010111100000100",
			2390 => "00000000000000000010010101110001",
			2391 => "00000001000101010010010101110001",
			2392 => "00000000000000000010010101110001",
			2393 => "0000000001000000001011101000000100",
			2394 => "11111110101111100010010101110001",
			2395 => "00000000000000000010010101110001",
			2396 => "0000000100000000000000010100000100",
			2397 => "11111110101100010010010111110101",
			2398 => "0000001000000000000111000100100100",
			2399 => "0000000000000000001110111100010100",
			2400 => "0000000110000000001011001100001000",
			2401 => "0000000110000000001101011000000100",
			2402 => "00000000000000000010010111110101",
			2403 => "11111111110110100010010111110101",
			2404 => "0000001100000000001110001100000100",
			2405 => "00000000000000000010010111110101",
			2406 => "0000001100000000001001110100000100",
			2407 => "00000000010110000010010111110101",
			2408 => "00000000000000000010010111110101",
			2409 => "0000001000000000001111001000000100",
			2410 => "00000000000000000010010111110101",
			2411 => "0000000000000000000111111000001000",
			2412 => "0000000011000000001010111100000100",
			2413 => "00000000000000000010010111110101",
			2414 => "00000001101110010010010111110101",
			2415 => "00000000000000000010010111110101",
			2416 => "0000000110000000000100111100011000",
			2417 => "0000000101000000001001110100001000",
			2418 => "0000000000000000001110001100000100",
			2419 => "11111111000101100010010111110101",
			2420 => "00000000000000000010010111110101",
			2421 => "0000000110000000001011001100000100",
			2422 => "00000000000000000010010111110101",
			2423 => "0000001001000000001010011000001000",
			2424 => "0000000100000000000010010000000100",
			2425 => "00000000000000000010010111110101",
			2426 => "00000001000101010010010111110101",
			2427 => "00000000000000000010010111110101",
			2428 => "11111110110010110010010111110101",
			2429 => "0000000100000000000011010100001100",
			2430 => "0000000010000000000101000000000100",
			2431 => "11111110011110100010011010001001",
			2432 => "0000001111000000000101000000000100",
			2433 => "00000001001010010010011010001001",
			2434 => "11111110101000000010011010001001",
			2435 => "0000000001000000001001111000011000",
			2436 => "0000001000000000000111000100001000",
			2437 => "0000001000000000001111001000000100",
			2438 => "11111111010100010010011010001001",
			2439 => "00000110110101100010011010001001",
			2440 => "0000000010000000001000101000001100",
			2441 => "0000000001000000000010001100000100",
			2442 => "11111110011100010010011010001001",
			2443 => "0000000001000000000010001100000100",
			2444 => "00000000001110000010011010001001",
			2445 => "11111110110000010010011010001001",
			2446 => "00000000000000000010011010001001",
			2447 => "0000000010000000000011110000100100",
			2448 => "0000000011000000001010011100001000",
			2449 => "0000000101000000000011100000000100",
			2450 => "00000000000000000010011010001001",
			2451 => "00000001110000000010011010001001",
			2452 => "0000000110000000001011001100001100",
			2453 => "0000001100000000001100110000000100",
			2454 => "00000000000000000010011010001001",
			2455 => "0000000010000000000000010000000100",
			2456 => "00000000000000000010011010001001",
			2457 => "11111101101101100010011010001001",
			2458 => "0000000100000000000000101100001000",
			2459 => "0000001011000000001000000000000100",
			2460 => "11111110100111110010011010001001",
			2461 => "00000001010010100010011010001001",
			2462 => "0000000001000000001101011100000100",
			2463 => "00000001100001000010011010001001",
			2464 => "11111110111010110010011010001001",
			2465 => "11111110011100110010011010001001",
			2466 => "0000000100000000001001000000011100",
			2467 => "0000000100000000000100001100000100",
			2468 => "11111110011100110010011100000101",
			2469 => "0000000000000000001110111100010100",
			2470 => "0000000010000000000100101000000100",
			2471 => "00000101011111010010011100000101",
			2472 => "0000001010000000001010110000001100",
			2473 => "0000000010000000001111100100000100",
			2474 => "11111110111010100010011100000101",
			2475 => "0000000101000000000110010000000100",
			2476 => "00000010001101010010011100000101",
			2477 => "00000000000000000010011100000101",
			2478 => "11111110110010010010011100000101",
			2479 => "11111110011011010010011100000101",
			2480 => "0000000001000000001100110100000100",
			2481 => "11111110011010010010011100000101",
			2482 => "0000000110000000001000010000011100",
			2483 => "0000001100000000000000101000000100",
			2484 => "00001010100001100010011100000101",
			2485 => "0000000001000000001001111000001000",
			2486 => "0000001110000000000101101100000100",
			2487 => "00000001010110100010011100000101",
			2488 => "11111101110111100010011100000101",
			2489 => "0000000010000000001011111000001000",
			2490 => "0000000110000000001001100100000100",
			2491 => "00000010100111110010011100000101",
			2492 => "00000000000000000010011100000101",
			2493 => "0000000001000000001101011100000100",
			2494 => "00000001011110000010011100000101",
			2495 => "11111110100000000010011100000101",
			2496 => "11111110010111110010011100000101",
			2497 => "0000001001000000001101101000000100",
			2498 => "11111111001110000010011101111001",
			2499 => "0000001100000000000011011100011000",
			2500 => "0000001101000000001011000000000100",
			2501 => "00000000000000000010011101111001",
			2502 => "0000001100000000001000111000000100",
			2503 => "00000000000000000010011101111001",
			2504 => "0000001000000000001001101000000100",
			2505 => "00000000000000000010011101111001",
			2506 => "0000000110000000001000010000001000",
			2507 => "0000000111000000001001110000000100",
			2508 => "00000000000000000010011101111001",
			2509 => "00000000111111100010011101111001",
			2510 => "00000000000000000010011101111001",
			2511 => "0000000010000000000011110000011100",
			2512 => "0000001011000000000100011000001100",
			2513 => "0000000100000000001101000000001000",
			2514 => "0000001110000000000000001100000100",
			2515 => "00000000000000000010011101111001",
			2516 => "11111111100001100010011101111001",
			2517 => "00000000000000000010011101111001",
			2518 => "0000001010000000000110011000000100",
			2519 => "00000000000000000010011101111001",
			2520 => "0000000001000000001011101000000100",
			2521 => "00000000000000000010011101111001",
			2522 => "0000000001000000000101011100000100",
			2523 => "00000000101010110010011101111001",
			2524 => "00000000000000000010011101111001",
			2525 => "11111111010011100010011101111001",
			2526 => "0000000001000000001001111000011000",
			2527 => "0000001101000000000100011000000100",
			2528 => "11111110011010000010011111111101",
			2529 => "0000000101000000000111001000000100",
			2530 => "00001000101101010010011111111101",
			2531 => "0000000111000000000110000100001100",
			2532 => "0000001101000000000011100000000100",
			2533 => "11111111001010000010011111111101",
			2534 => "0000001101000000001011000000000100",
			2535 => "00000000010110010010011111111101",
			2536 => "11111111111111110010011111111101",
			2537 => "11111110010110110010011111111101",
			2538 => "0000001010000000000110011000000100",
			2539 => "11111110011010110010011111111101",
			2540 => "0000000110000000000101010000100100",
			2541 => "0000000101000000000011100000001000",
			2542 => "0000001110000000000101101100000100",
			2543 => "00000000000000000010011111111101",
			2544 => "11111110100110000010011111111101",
			2545 => "0000000010000000000110010000001100",
			2546 => "0000001110000000000001101000001000",
			2547 => "0000000000000000000000111000000100",
			2548 => "11111111101100100010011111111101",
			2549 => "00000010001000100010011111111101",
			2550 => "00000110010010000010011111111101",
			2551 => "0000000110000000001011001100001000",
			2552 => "0000000001000000001101101000000100",
			2553 => "00000001000010010010011111111101",
			2554 => "11111101100000010010011111111101",
			2555 => "0000000010000000001000001100000100",
			2556 => "11111111000000000010011111111101",
			2557 => "00000001010011000010011111111101",
			2558 => "11111110011011010010011111111101",
			2559 => "0000000111000000001001110000001000",
			2560 => "0000001010000000000110001000000100",
			2561 => "11111110111000010010100010010001",
			2562 => "00000000000000000010100010010001",
			2563 => "0000000010000000000111111100010000",
			2564 => "0000000010000000001001010000000100",
			2565 => "00000000000000000010100010010001",
			2566 => "0000000100000000000010111000000100",
			2567 => "00000000000000000010100010010001",
			2568 => "0000000111000000001110001100000100",
			2569 => "00000001001001010010100010010001",
			2570 => "00000000000000000010100010010001",
			2571 => "0000000100000000001011001000001100",
			2572 => "0000000010000000001110100100000100",
			2573 => "11111110111101100010100010010001",
			2574 => "0000000011000000001111101000000100",
			2575 => "00000000011100110010100010010001",
			2576 => "00000000000000000010100010010001",
			2577 => "0000000000000000001100001000010000",
			2578 => "0000000011000000001001011100001100",
			2579 => "0000000111000000001010111100001000",
			2580 => "0000001100000000001101111000000100",
			2581 => "00000001000000110010100010010001",
			2582 => "00000000000000000010100010010001",
			2583 => "00000000000000000010100010010001",
			2584 => "00000000000000000010100010010001",
			2585 => "0000000100000000001101000000001000",
			2586 => "0000001001000000000100110100000100",
			2587 => "11111111000011100010100010010001",
			2588 => "00000000000000000010100010010001",
			2589 => "0000001110000000001110110000001000",
			2590 => "0000001100000000000110000100000100",
			2591 => "00000000000000000010100010010001",
			2592 => "11111111100100010010100010010001",
			2593 => "0000000011000000001100010000000100",
			2594 => "00000000011001110010100010010001",
			2595 => "00000000000000000010100010010001",
			2596 => "0000000100000000000000010100000100",
			2597 => "11111110101010110010100100011101",
			2598 => "0000001000000000000111000100101000",
			2599 => "0000000000000000001110111100011000",
			2600 => "0000000110000000001011001100001000",
			2601 => "0000001011000000000000001100000100",
			2602 => "00000000000000000010100100011101",
			2603 => "11111111101011110010100100011101",
			2604 => "0000001011000000000011100000000100",
			2605 => "00000000000000000010100100011101",
			2606 => "0000001010000000001010110000001000",
			2607 => "0000001110000000001101101100000100",
			2608 => "00000000011110110010100100011101",
			2609 => "00000000000000000010100100011101",
			2610 => "00000000000000000010100100011101",
			2611 => "0000001000000000001111001000000100",
			2612 => "00000000000000000010100100011101",
			2613 => "0000000000000000000111111000001000",
			2614 => "0000000011000000001010111100000100",
			2615 => "00000000000000000010100100011101",
			2616 => "00000001110011010010100100011101",
			2617 => "00000000000000000010100100011101",
			2618 => "0000000110000000000100111100011000",
			2619 => "0000000101000000001001110100001000",
			2620 => "0000000000000000001110001100000100",
			2621 => "11111111000010000010100100011101",
			2622 => "00000000000000000010100100011101",
			2623 => "0000000110000000001011001100000100",
			2624 => "00000000000000000010100100011101",
			2625 => "0000001010000000001100011100000100",
			2626 => "00000000000000000010100100011101",
			2627 => "0000000100000000000001100100000100",
			2628 => "00000000000000000010100100011101",
			2629 => "00000001000111010010100100011101",
			2630 => "11111110110000010010100100011101",
			2631 => "0000000100000000000011010100011100",
			2632 => "0000000110000000001011001100000100",
			2633 => "11111110011010010010100111011001",
			2634 => "0000000110000000001011001100001100",
			2635 => "0000001001000000000001000100000100",
			2636 => "11111111011110100010100111011001",
			2637 => "0000001101000000000000110100000100",
			2638 => "00000101011100010010100111011001",
			2639 => "00000000000000000010100111011001",
			2640 => "0000001001000000001101011000001000",
			2641 => "0000000001000000001111001100000100",
			2642 => "11111110101011100010100111011001",
			2643 => "00000001001011010010100111011001",
			2644 => "11111110011101000010100111011001",
			2645 => "0000000001000000001001111000011100",
			2646 => "0000000000000000000111111000001000",
			2647 => "0000000000000000000111111000000100",
			2648 => "11111111010000000010100111011001",
			2649 => "00000101000000000010100111011001",
			2650 => "0000001001000000001101101000000100",
			2651 => "11111110011001000010100111011001",
			2652 => "0000000001000000000010001100001100",
			2653 => "0000000001000000000010001100001000",
			2654 => "0000001001000000001101101000000100",
			2655 => "00000000000000000010100111011001",
			2656 => "11111111011010100010100111011001",
			2657 => "00000000011001110010100111011001",
			2658 => "11111110101111010010100111011001",
			2659 => "0000000110000000000101010000100100",
			2660 => "0000000011000000001010011100001000",
			2661 => "0000000101000000000011100000000100",
			2662 => "00000000000000000010100111011001",
			2663 => "00000001101111110010100111011001",
			2664 => "0000000110000000001011001100001100",
			2665 => "0000001100000000001100110000000100",
			2666 => "00000000000000000010100111011001",
			2667 => "0000001100000000001110001100000100",
			2668 => "11111101111100110010100111011001",
			2669 => "00000000000000000010100111011001",
			2670 => "0000000001000000000111100100001000",
			2671 => "0000000100000000000000000000000100",
			2672 => "11111110110011000010100111011001",
			2673 => "00000000101011000010100111011001",
			2674 => "0000000001000000001101011100000100",
			2675 => "00000001011011010010100111011001",
			2676 => "00000000010101100010100111011001",
			2677 => "11111110011110000010100111011001",
			2678 => "0000001011000000000101101100000100",
			2679 => "11111110100010000010101001100101",
			2680 => "0000001111000000001010010100001100",
			2681 => "0000001111000000000010001000000100",
			2682 => "00000000000000000010101001100101",
			2683 => "0000000100000000001110111000000100",
			2684 => "00000000000000000010101001100101",
			2685 => "00000010100111110010101001100101",
			2686 => "0000001001000000000100110100011000",
			2687 => "0000000100000000001010010000010000",
			2688 => "0000001111000000001110101100000100",
			2689 => "00000000000000000010101001100101",
			2690 => "0000001001000000001110010100000100",
			2691 => "11111110101100010010101001100101",
			2692 => "0000001001000000000100110100000100",
			2693 => "00000000000000000010101001100101",
			2694 => "11111111000011110010101001100101",
			2695 => "0000000101000000001011011100000100",
			2696 => "00000000101011010010101001100101",
			2697 => "00000000000000000010101001100101",
			2698 => "0000000001000000001001011000010000",
			2699 => "0000000110000000001011001100000100",
			2700 => "11111111111011000010101001100101",
			2701 => "0000000000000000001011000100001000",
			2702 => "0000000101000000000101100100000100",
			2703 => "00000000000000000010101001100101",
			2704 => "00000001001011010010101001100101",
			2705 => "00000000000000000010101001100101",
			2706 => "0000000001000000000101011100001100",
			2707 => "0000001101000000001001010100000100",
			2708 => "11111111000110010010101001100101",
			2709 => "0000000100000000000011010100000100",
			2710 => "00000000000000000010101001100101",
			2711 => "00000000110011000010101001100101",
			2712 => "11111111000000000010101001100101",
			2713 => "0000000001000000001001111000000100",
			2714 => "11111110100000110010101100000001",
			2715 => "0000001100000000001100110000100000",
			2716 => "0000001100000000001000111000001000",
			2717 => "0000000100000000001101000000000100",
			2718 => "11111110111001100010101100000001",
			2719 => "00000000000000000010101100000001",
			2720 => "0000001100000000000011011100010000",
			2721 => "0000000000000000000010111100000100",
			2722 => "00000000000000000010101100000001",
			2723 => "0000001010000000000001010000000100",
			2724 => "00000010000101010010101100000001",
			2725 => "0000001010000000001100011100000100",
			2726 => "00000000000000000010101100000001",
			2727 => "00000001000011100010101100000001",
			2728 => "0000000100000000000010010000000100",
			2729 => "11111111010010000010101100000001",
			2730 => "00000001000001100010101100000001",
			2731 => "0000000101000000000000011100010000",
			2732 => "0000001000000000001111000100001100",
			2733 => "0000001100000000000110000100001000",
			2734 => "0000000010000000001111100100000100",
			2735 => "00000000000000000010101100000001",
			2736 => "11111110000100100010101100000001",
			2737 => "00000000000000000010101100000001",
			2738 => "00000000000001100010101100000001",
			2739 => "0000000100000000000000010100000100",
			2740 => "11111110110101010010101100000001",
			2741 => "0000001010000000001100011100001100",
			2742 => "0000000001000000000101011100001000",
			2743 => "0000001011000000000011100000000100",
			2744 => "00000000000000000010101100000001",
			2745 => "00000001001101000010101100000001",
			2746 => "00000000000000000010101100000001",
			2747 => "0000000000000000000100010100000100",
			2748 => "11111111001100010010101100000001",
			2749 => "0000001100000000000100001000000100",
			2750 => "00000000111010000010101100000001",
			2751 => "11111111011111110010101100000001",
			2752 => "0000001101000000000100011000000100",
			2753 => "11111110011100010010101110100101",
			2754 => "0000001100000000000011011100011100",
			2755 => "0000001110000000000100001000001100",
			2756 => "0000000100000000001110111000000100",
			2757 => "00000000000000000010101110100101",
			2758 => "0000000011000000001001110100000100",
			2759 => "00000001110011010010101110100101",
			2760 => "00000000000000000010101110100101",
			2761 => "0000001100000000000011011100001000",
			2762 => "0000000100000000001101000000000100",
			2763 => "11111110100111010010101110100101",
			2764 => "00000000001111100010101110100101",
			2765 => "0000001001000000000001000100000100",
			2766 => "00000000000000000010101110100101",
			2767 => "00000010000101000010101110100101",
			2768 => "0000001011000000000000001100010000",
			2769 => "0000001011000000000000001100001000",
			2770 => "0000000000000000000011011100000100",
			2771 => "11111111010000000010101110100101",
			2772 => "00000000000000000010101110100101",
			2773 => "0000000001000000000110101000000100",
			2774 => "00000000000000000010101110100101",
			2775 => "11110000111000100010101110100101",
			2776 => "0000001100000000001010111000100000",
			2777 => "0000000001000000001011101000010000",
			2778 => "0000001000000000001101010000001000",
			2779 => "0000000010000000001011101100000100",
			2780 => "00000000000000000010101110100101",
			2781 => "11111110000110110010101110100101",
			2782 => "0000000001000000001001111000000100",
			2783 => "11111111000110110010101110100101",
			2784 => "00000001001001000010101110100101",
			2785 => "0000001010000000000110011000001000",
			2786 => "0000000010000000001111100100000100",
			2787 => "11111111000101100010101110100101",
			2788 => "00000000000000000010101110100101",
			2789 => "0000000010000000000110101100000100",
			2790 => "00000001010000100010101110100101",
			2791 => "00000000001111110010101110100101",
			2792 => "11111110101100010010101110100101",
			2793 => "0000000100000000001110111000000100",
			2794 => "11111110100000010010110001010001",
			2795 => "0000001000000000000111000100111000",
			2796 => "0000001000000000000111000100100000",
			2797 => "0000001000000000000110001000011000",
			2798 => "0000000100000000000011101100001100",
			2799 => "0000001110000000001101101100001000",
			2800 => "0000001010000000000110011000000100",
			2801 => "00000000000000000010110001010001",
			2802 => "00000001010000000010110001010001",
			2803 => "00000000000000000010110001010001",
			2804 => "0000000010000000001011111000001000",
			2805 => "0000001111000000000011001000000100",
			2806 => "00000000000000000010110001010001",
			2807 => "00000000011011110010110001010001",
			2808 => "11111111011001010010110001010001",
			2809 => "0000000100000000000000101100000100",
			2810 => "11111111011010100010110001010001",
			2811 => "00000000000000000010110001010001",
			2812 => "0000001111000000000101110100001000",
			2813 => "0000000100000000000011010100000100",
			2814 => "00000000000000000010110001010001",
			2815 => "00000110100001010010110001010001",
			2816 => "0000000001000000001101011100001100",
			2817 => "0000000100000000000100001100000100",
			2818 => "00000000000000000010110001010001",
			2819 => "0000000101000000000111001000000100",
			2820 => "00000000000000000010110001010001",
			2821 => "00000001100011100010110001010001",
			2822 => "00000000000000000010110001010001",
			2823 => "0000000100000000001010010000010000",
			2824 => "0000001001000000000100110100000100",
			2825 => "11111110111100000010110001010001",
			2826 => "0000000001000000001101011100001000",
			2827 => "0000001111000000001110000000000100",
			2828 => "00000000011001010010110001010001",
			2829 => "00000000000000000010110001010001",
			2830 => "11111111111111000010110001010001",
			2831 => "0000001001000000001101101000000100",
			2832 => "11111111011010100010110001010001",
			2833 => "0000000010000000001110000000000100",
			2834 => "00000000110011100010110001010001",
			2835 => "00000000000000000010110001010001",
			2836 => "0000001101000000000100011000000100",
			2837 => "11111110100100000010110011111101",
			2838 => "0000001111000000000110010000111100",
			2839 => "0000000111000000001101100000011000",
			2840 => "0000000110000000001011001100010000",
			2841 => "0000000000000000000010111100000100",
			2842 => "00000000000000000010110011111101",
			2843 => "0000001010000000001010110000001000",
			2844 => "0000000111000000001001110000000100",
			2845 => "00000000000000000010110011111101",
			2846 => "00000010000001010010110011111101",
			2847 => "00000000000000000010110011111101",
			2848 => "0000000000000000000100001000000100",
			2849 => "11111111111010100010110011111101",
			2850 => "00000000000000000010110011111101",
			2851 => "0000000110000000001011001100010100",
			2852 => "0000001100000000001100110000001100",
			2853 => "0000000000000000000000111000000100",
			2854 => "11111111101000010010110011111101",
			2855 => "0000000101000000000011100000000100",
			2856 => "00000000000000000010110011111101",
			2857 => "00000000101110100010110011111101",
			2858 => "0000000110000000001011001100000100",
			2859 => "11111110111000110010110011111101",
			2860 => "00000000000000000010110011111101",
			2861 => "0000000100000000001101110100000100",
			2862 => "00000000000000000010110011111101",
			2863 => "0000001011000000001000000000001000",
			2864 => "0000001000000000000110001000000100",
			2865 => "00000000000000000010110011111101",
			2866 => "00000001010011010010110011111101",
			2867 => "00000000000000000010110011111101",
			2868 => "0000000101000000000100010000001000",
			2869 => "0000001111000000001001100000000100",
			2870 => "00000000000000000010110011111101",
			2871 => "11111110100111010010110011111101",
			2872 => "0000001100000000001010111000001100",
			2873 => "0000000100000000000011010100000100",
			2874 => "00000000000000000010110011111101",
			2875 => "0000001101000000001110101100000100",
			2876 => "00000000000000000010110011111101",
			2877 => "00000000111101000010110011111101",
			2878 => "11111111011001110010110011111101",
			2879 => "0000000111000000001001110000001000",
			2880 => "0000001000000000000000111000000100",
			2881 => "11111111000001100010110110011001",
			2882 => "00000000000000000010110110011001",
			2883 => "0000000111000000001101100000010100",
			2884 => "0000000010000000000110010000010000",
			2885 => "0000001110000000001001110000000100",
			2886 => "00000000000000000010110110011001",
			2887 => "0000001000000000001001101000000100",
			2888 => "00000000000000000010110110011001",
			2889 => "0000001101000000000100011000000100",
			2890 => "00000000000000000010110110011001",
			2891 => "00000001011111110010110110011001",
			2892 => "00000000000000000010110110011001",
			2893 => "0000000100000000000000010100000100",
			2894 => "11111111010000000010110110011001",
			2895 => "0000000000000000000011111100010000",
			2896 => "0000001100000000001110001100000100",
			2897 => "00000000000000000010110110011001",
			2898 => "0000000001000000000101011100001000",
			2899 => "0000000101000000001011011100000100",
			2900 => "00000000000000000010110110011001",
			2901 => "00000000101101000010110110011001",
			2902 => "00000000000000000010110110011001",
			2903 => "0000000110000000001011001100010000",
			2904 => "0000001100000000000110000100001000",
			2905 => "0000000100000000000001100100000100",
			2906 => "00000000000000000010110110011001",
			2907 => "00000000110000110010110110011001",
			2908 => "0000000110000000001011001100000100",
			2909 => "11111111100110110010110110011001",
			2910 => "00000000000000000010110110011001",
			2911 => "0000000100000000001101000000001000",
			2912 => "0000000011000000001000001100000100",
			2913 => "11111111010001010010110110011001",
			2914 => "00000000000000000010110110011001",
			2915 => "0000001000000000001010000000000100",
			2916 => "00000000000010100010110110011001",
			2917 => "00000000000000000010110110011001",
			2918 => "0000001101000000000100011000000100",
			2919 => "11111110011011100010111001000101",
			2920 => "0000001100000000001100110000101100",
			2921 => "0000001100000000001001110000010100",
			2922 => "0000001110000000000100001000001100",
			2923 => "0000000100000000000111011100000100",
			2924 => "11111111111110010010111001000101",
			2925 => "0000000110000000001001100100000100",
			2926 => "00000001110100110010111001000101",
			2927 => "00000000000000000010111001000101",
			2928 => "0000000100000000001101000000000100",
			2929 => "11111110100011110010111001000101",
			2930 => "00000000000000000010111001000101",
			2931 => "0000000000000000000010111100000100",
			2932 => "11111111111101000010111001000101",
			2933 => "0000001010000000000001010000000100",
			2934 => "00000010111100100010111001000101",
			2935 => "0000000000000000000111111000001000",
			2936 => "0000000000000000001010000000000100",
			2937 => "11111111110011010010111001000101",
			2938 => "00000000000000000010111001000101",
			2939 => "0000000001000000001001111000000100",
			2940 => "00000000000000000010111001000101",
			2941 => "00000001100011010010111001000101",
			2942 => "0000000110000000001101011000001000",
			2943 => "0000001100000000001100110000000100",
			2944 => "00000000000000000010111001000101",
			2945 => "11111110001111110010111001000101",
			2946 => "0000000001000000000101011100011100",
			2947 => "0000000000000000000000111000001100",
			2948 => "0000000101000000000101100100000100",
			2949 => "11111111011110110010111001000101",
			2950 => "0000001010000000000110011000000100",
			2951 => "00000000000000000010111001000101",
			2952 => "00000001010111000010111001000101",
			2953 => "0000001111000000000111011000001000",
			2954 => "0000000000000000001000111100000100",
			2955 => "11111111011100010010111001000101",
			2956 => "00000001001101110010111001000101",
			2957 => "0000000001000000001101011100000100",
			2958 => "11111110100000100010111001000101",
			2959 => "00000000000000000010111001000101",
			2960 => "11111110100010110010111001000101",
			2961 => "0000001101000000000100011000000100",
			2962 => "11111110011100000010111011010001",
			2963 => "0000001000000000001001101000000100",
			2964 => "11111110100011010010111011010001",
			2965 => "0000001010000000000001010000011000",
			2966 => "0000001100000000001001110000000100",
			2967 => "11111111101001010010111011010001",
			2968 => "0000000010000000001011111000001000",
			2969 => "0000001000000000001001101000000100",
			2970 => "00000000000000000010111011010001",
			2971 => "00000010000110000010111011010001",
			2972 => "0000000011000000000111100000000100",
			2973 => "00000000000000000010111011010001",
			2974 => "0000000011000000001111101000000100",
			2975 => "00000001000001100010111011010001",
			2976 => "00000000000000000010111011010001",
			2977 => "0000001110000000001101010100010100",
			2978 => "0000001100000000000110000100001100",
			2979 => "0000000100000000000111011100000100",
			2980 => "11111111101001010010111011010001",
			2981 => "0000000001000000001100110100000100",
			2982 => "00000000000000000010111011010001",
			2983 => "00000001100011000010111011010001",
			2984 => "0000000001000000001001111000000100",
			2985 => "11111110110111110010111011010001",
			2986 => "00000000000000000010111011010001",
			2987 => "0000001101000000001010001100001000",
			2988 => "0000000100000000001010101000000100",
			2989 => "11111110010110100010111011010001",
			2990 => "00000000000000000010111011010001",
			2991 => "0000001100000000001010111000001000",
			2992 => "0000001100000000000000001100000100",
			2993 => "11111111111111010010111011010001",
			2994 => "00000000111110100010111011010001",
			2995 => "11111110100111000010111011010001",
			2996 => "0000001101000000000100011000000100",
			2997 => "11111110101011000010111101111101",
			2998 => "0000001000000000000111000100110000",
			2999 => "0000000000000000000010011000001000",
			3000 => "0000000100000000000000010100000100",
			3001 => "11111111001101000010111101111101",
			3002 => "00000000000000000010111101111101",
			3003 => "0000000000000000000010111100010000",
			3004 => "0000001010000000000001010000001100",
			3005 => "0000000101000000001000000000000100",
			3006 => "00000000000000000010111101111101",
			3007 => "0000000001000000000101011100000100",
			3008 => "00000001101001110010111101111101",
			3009 => "00000000000000000010111101111101",
			3010 => "00000000000000000010111101111101",
			3011 => "0000000000000000001110111100010000",
			3012 => "0000001010000000000001010000001000",
			3013 => "0000001100000000001110001100000100",
			3014 => "00000000000000000010111101111101",
			3015 => "00000000110010110010111101111101",
			3016 => "0000001100000000000000001100000100",
			3017 => "11111111001111010010111101111101",
			3018 => "00000000000000000010111101111101",
			3019 => "0000001001000000001101011000000100",
			3020 => "00000001011010110010111101111101",
			3021 => "00000000000000000010111101111101",
			3022 => "0000000110000000000100111100100000",
			3023 => "0000000001000000001111001100011000",
			3024 => "0000001001000000001001011000001100",
			3025 => "0000000011000000001110110000000100",
			3026 => "00000000000000000010111101111101",
			3027 => "0000000000000000001010111100000100",
			3028 => "11111111010000110010111101111101",
			3029 => "00000000000000000010111101111101",
			3030 => "0000000100000000000110110000000100",
			3031 => "00000000000000000010111101111101",
			3032 => "0000000110000000001011001100000100",
			3033 => "00000000000000000010111101111101",
			3034 => "00000001000001100010111101111101",
			3035 => "0000000110000000001001100100000100",
			3036 => "11111111001111110010111101111101",
			3037 => "00000000000000000010111101111101",
			3038 => "11111110110111000010111101111101",
			3039 => "0000001011000000000101101100000100",
			3040 => "11111110011101100011000000001011",
			3041 => "0000000100000000000010111000000100",
			3042 => "11111110100101000011000000001011",
			3043 => "0000001000000000000111000100011000",
			3044 => "0000000001000000000101011100010100",
			3045 => "0000000010000000000011001000000100",
			3046 => "00000010001011110011000000001011",
			3047 => "0000001101000000000101110100001000",
			3048 => "0000000000000000001110111100000100",
			3049 => "11111110111101110011000000001011",
			3050 => "00000000000000000011000000001011",
			3051 => "0000001110000000000111110000000100",
			3052 => "00000000000000000011000000001011",
			3053 => "00000001011110100011000000001011",
			3054 => "11111111010010110011000000001011",
			3055 => "0000001100000000000110000100010000",
			3056 => "0000000100000000000001100100000100",
			3057 => "11111110110011010011000000001011",
			3058 => "0000000010000000000010010100001000",
			3059 => "0000001100000000001100110000000100",
			3060 => "00000001011101100011000000001011",
			3061 => "00000000000000000011000000001011",
			3062 => "11111111100000000011000000001011",
			3063 => "0000001101000000000100000100001100",
			3064 => "0000000101000000001010011100001000",
			3065 => "0000001011000000001010111100000100",
			3066 => "11111101101110000011000000001011",
			3067 => "00000000000000000011000000001011",
			3068 => "00000000000000000011000000001011",
			3069 => "0000001100000000000100001000001000",
			3070 => "0000000000000000000100010100000100",
			3071 => "11111111101000010011000000001011",
			3072 => "00000001000111110011000000001011",
			3073 => "11111111000100010011000000001011",
			3074 => "00000000000000000011000000001101",
			3075 => "00000000000000000011000000010001",
			3076 => "00000000000000000011000000010101",
			3077 => "00000000000000000011000000011001",
			3078 => "00000000000000000011000000011101",
			3079 => "00000000000000000011000000100001",
			3080 => "00000000000000000011000000100101",
			3081 => "00000000000000000011000000101001",
			3082 => "00000000000000000011000000101101",
			3083 => "0000000100000000001110111000000100",
			3084 => "11111111110111010011000000111001",
			3085 => "00000000000000000011000000111001",
			3086 => "0000000110000000001011001100000100",
			3087 => "11111111111001100011000001001101",
			3088 => "0000000110000000001000010000000100",
			3089 => "00000000000010000011000001001101",
			3090 => "00000000000000000011000001001101",
			3091 => "0000000001000000001011101000000100",
			3092 => "11111111111111110011000001100001",
			3093 => "0000000001000000000000111100000100",
			3094 => "00000000000001100011000001100001",
			3095 => "00000000000000000011000001100001",
			3096 => "0000000011000000000101110100001000",
			3097 => "0000000110000000001001100100000100",
			3098 => "11111111110111010011000001110101",
			3099 => "00000000000000000011000001110101",
			3100 => "00000000000000000011000001110101",
			3101 => "0000001110000000001110101100001000",
			3102 => "0000000100000000001101000000000100",
			3103 => "11111111110001000011000010001001",
			3104 => "00000000000000000011000010001001",
			3105 => "00000000000000000011000010001001",
			3106 => "0000001110000000001100101100000100",
			3107 => "00000000000000000011000010011101",
			3108 => "0000001110000000001101101100000100",
			3109 => "00000000000100000011000010011101",
			3110 => "00000000000000000011000010011101",
			3111 => "0000001111000000000110010000001000",
			3112 => "0000001111000000000010001000000100",
			3113 => "00000000000000000011000010111001",
			3114 => "00000000000111100011000010111001",
			3115 => "0000001111000000001011110000000100",
			3116 => "11111111111000000011000010111001",
			3117 => "00000000000000000011000010111001",
			3118 => "0000000010000000000100101000000100",
			3119 => "00000000000000000011000011010101",
			3120 => "0000001110000000001010000100001000",
			3121 => "0000000000000000000100010100000100",
			3122 => "11111111011010000011000011010101",
			3123 => "00000000000000000011000011010101",
			3124 => "00000000000000000011000011010101",
			3125 => "0000000010000000000100101000000100",
			3126 => "00000000000000000011000011110001",
			3127 => "0000000100000000000011011000001000",
			3128 => "0000001111000000001011110000000100",
			3129 => "11111111011101010011000011110001",
			3130 => "00000000000000000011000011110001",
			3131 => "00000000000000000011000011110001",
			3132 => "0000000001000000001101011100001100",
			3133 => "0000000001000000001100110100000100",
			3134 => "00000000000000000011000100001101",
			3135 => "0000000001000000001111001100000100",
			3136 => "00000000001010000011000100001101",
			3137 => "00000000000000000011000100001101",
			3138 => "11111111111111110011000100001101",
			3139 => "0000000011000000000010001000000100",
			3140 => "11111111111011100011000100101001",
			3141 => "0000001001000000000100111100001000",
			3142 => "0000001001000000000001000100000100",
			3143 => "00000000000000000011000100101001",
			3144 => "00000000000101010011000100101001",
			3145 => "00000000000000000011000100101001",
			3146 => "0000001100000000001100110000001000",
			3147 => "0000001101000000000110100100000100",
			3148 => "00000000000000000011000101001101",
			3149 => "00000000000011010011000101001101",
			3150 => "0000001111000000001011110000001000",
			3151 => "0000000111000000000110000100000100",
			3152 => "00000000000000000011000101001101",
			3153 => "11111111110111100011000101001101",
			3154 => "00000000000000000011000101001101",
			3155 => "0000001111000000000010000000001000",
			3156 => "0000001111000000000010001000000100",
			3157 => "00000000000000000011000101110001",
			3158 => "00000000000000100011000101110001",
			3159 => "0000001111000000001000110100001000",
			3160 => "0000001111000000000110010000000100",
			3161 => "00000000000000000011000101110001",
			3162 => "11111111110101010011000101110001",
			3163 => "00000000000000000011000101110001",
			3164 => "0000001100000000000011011100001100",
			3165 => "0000000111000000001001110000000100",
			3166 => "00000000000000000011000110011101",
			3167 => "0000001011000000001100110000000100",
			3168 => "00000000000000000011000110011101",
			3169 => "00000000000100110011000110011101",
			3170 => "0000000011000000000011000000001000",
			3171 => "0000000111000000000110000100000100",
			3172 => "00000000000000000011000110011101",
			3173 => "11111111110111010011000110011101",
			3174 => "00000000000000000011000110011101",
			3175 => "0000000100000000001100111100001100",
			3176 => "0000000010000000000100101000000100",
			3177 => "00000000000000000011000111001001",
			3178 => "0000000010000000001110100100000100",
			3179 => "11111111100011000011000111001001",
			3180 => "00000000000000000011000111001001",
			3181 => "0000001101000000000001011000000100",
			3182 => "00000000000000000011000111001001",
			3183 => "0000001101000000001001010000000100",
			3184 => "00000000000111010011000111001001",
			3185 => "00000000000000000011000111001001",
			3186 => "0000000010000000000100101000000100",
			3187 => "00000000000000000011000111101101",
			3188 => "0000000100000000000010010000001100",
			3189 => "0000001111000000001011110000001000",
			3190 => "0000001111000000000101110100000100",
			3191 => "00000000000000000011000111101101",
			3192 => "11111111010111010011000111101101",
			3193 => "00000000000000000011000111101101",
			3194 => "00000000000000000011000111101101",
			3195 => "0000001100000000001100110000010000",
			3196 => "0000000001000000001100110100000100",
			3197 => "00000000000000000011001000010001",
			3198 => "0000000001000000001111001100001000",
			3199 => "0000001100000000000000101000000100",
			3200 => "00000000000000000011001000010001",
			3201 => "00000000010001100011001000010001",
			3202 => "00000000000000000011001000010001",
			3203 => "11111111111111100011001000010001",
			3204 => "0000000101000000001011011100010000",
			3205 => "0000000100000000001010010000001100",
			3206 => "0000000010000000001010001000000100",
			3207 => "00000000000000000011001000110101",
			3208 => "0000001111000000000101110100000100",
			3209 => "00000000000000000011001000110101",
			3210 => "11111111101010010011001000110101",
			3211 => "00000000000000000011001000110101",
			3212 => "00000000000000000011001000110101",
			3213 => "0000000000000000001110111100001000",
			3214 => "0000000000000000000010111100000100",
			3215 => "00000000000000000011001001100001",
			3216 => "11111111110100110011001001100001",
			3217 => "0000001000000000000001110100001100",
			3218 => "0000000111000000001001110000000100",
			3219 => "00000000000000000011001001100001",
			3220 => "0000000111000000001101010100000100",
			3221 => "00000000010100100011001001100001",
			3222 => "00000000000000000011001001100001",
			3223 => "00000000000000000011001001100001",
			3224 => "0000000000000000001110111100001100",
			3225 => "0000000000000000000010111100000100",
			3226 => "00000000000000000011001010010101",
			3227 => "0000000100000000000000100000000100",
			3228 => "11111111110100010011001010010101",
			3229 => "00000000000000000011001010010101",
			3230 => "0000001000000000000001110100001100",
			3231 => "0000000111000000001001110000000100",
			3232 => "00000000000000000011001010010101",
			3233 => "0000000111000000001101010100000100",
			3234 => "00000000010010010011001010010101",
			3235 => "00000000000000000011001010010101",
			3236 => "00000000000000000011001010010101",
			3237 => "0000000000000000000011111100001100",
			3238 => "0000001010000000000110011000000100",
			3239 => "00000000000000000011001011001001",
			3240 => "0000001010000000000001010000000100",
			3241 => "00000000000100100011001011001001",
			3242 => "00000000000000000011001011001001",
			3243 => "0000001010000000000110011000000100",
			3244 => "00000000000000000011001011001001",
			3245 => "0000000000000000001010111100001000",
			3246 => "0000001100000000000000001100000100",
			3247 => "11111111110111110011001011001001",
			3248 => "00000000000000000011001011001001",
			3249 => "00000000000000000011001011001001",
			3250 => "0000000101000000001011011100010000",
			3251 => "0000000100000000001010010000001100",
			3252 => "0000000010000000001010001000000100",
			3253 => "00000000000000000011001011111101",
			3254 => "0000001111000000000101110100000100",
			3255 => "00000000000000000011001011111101",
			3256 => "11111111101100110011001011111101",
			3257 => "00000000000000000011001011111101",
			3258 => "0000001100000000001010111000001000",
			3259 => "0000001100000000001110001100000100",
			3260 => "00000000000000000011001011111101",
			3261 => "00000000000100000011001011111101",
			3262 => "00000000000000000011001011111101",
			3263 => "0000000100000000000001100100010000",
			3264 => "0000001010000000000001010000000100",
			3265 => "00000000000000000011001100111001",
			3266 => "0000001111000000000101110100000100",
			3267 => "00000000000000000011001100111001",
			3268 => "0000000000000000000010011000000100",
			3269 => "00000000000000000011001100111001",
			3270 => "11111111100111010011001100111001",
			3271 => "0000000001000000001111001100001100",
			3272 => "0000000001000000000010001100000100",
			3273 => "00000000000000000011001100111001",
			3274 => "0000001111000000001000001100000100",
			3275 => "00000000001011000011001100111001",
			3276 => "00000000000000000011001100111001",
			3277 => "00000000000000000011001100111001",
			3278 => "0000000001000000001101011100010100",
			3279 => "0000000001000000001100110100000100",
			3280 => "00000000000000000011001101100101",
			3281 => "0000000000000000000010111100000100",
			3282 => "00000000000000000011001101100101",
			3283 => "0000001010000000000001110000001000",
			3284 => "0000001010000000001001000100000100",
			3285 => "00000000000000000011001101100101",
			3286 => "00000000010000100011001101100101",
			3287 => "00000000000000000011001101100101",
			3288 => "00000000000000000011001101100101",
			3289 => "0000000110000000001101011000001000",
			3290 => "0000000100000000001110111000000100",
			3291 => "11111111110111110011001110100001",
			3292 => "00000000000000000011001110100001",
			3293 => "0000000110000000001001100100010000",
			3294 => "0000000001000000000111100100000100",
			3295 => "00000000000000000011001110100001",
			3296 => "0000000001000000000000111100001000",
			3297 => "0000000100000000001000000100000100",
			3298 => "00000000000000000011001110100001",
			3299 => "00000000010100110011001110100001",
			3300 => "00000000000000000011001110100001",
			3301 => "0000000100000000000011111000000100",
			3302 => "11111111111100010011001110100001",
			3303 => "00000000000000000011001110100001",
			3304 => "0000001001000000000100110100011100",
			3305 => "0000000010000000001110010000001100",
			3306 => "0000000011000000000011100000000100",
			3307 => "00000000000000000011001111101101",
			3308 => "0000001110000000000011100000000100",
			3309 => "00000000000111010011001111101101",
			3310 => "00000000000000000011001111101101",
			3311 => "0000000100000000001010010000001100",
			3312 => "0000001111000000000111110000000100",
			3313 => "00000000000000000011001111101101",
			3314 => "0000000101000000000100010000000100",
			3315 => "11111111011110110011001111101101",
			3316 => "00000000000000000011001111101101",
			3317 => "00000000000000000011001111101101",
			3318 => "0000000001000000001001011000001000",
			3319 => "0000001001000000001010011000000100",
			3320 => "00000000000000000011001111101101",
			3321 => "00000000001010010011001111101101",
			3322 => "00000000000000000011001111101101",
			3323 => "0000001100000000001100110000011000",
			3324 => "0000001100000000000100000000000100",
			3325 => "00000000000000000011010000110001",
			3326 => "0000000100000000001000000100000100",
			3327 => "00000000000000000011010000110001",
			3328 => "0000000011000000000100011000000100",
			3329 => "00000000000000000011010000110001",
			3330 => "0000000010000000000010010100001000",
			3331 => "0000000011000000001001011100000100",
			3332 => "00000000010011000011010000110001",
			3333 => "00000000000000000011010000110001",
			3334 => "00000000000000000011010000110001",
			3335 => "0000000010000000000011000000001000",
			3336 => "0000000010000000000110101100000100",
			3337 => "00000000000000000011010000110001",
			3338 => "11111111110100100011010000110001",
			3339 => "00000000000000000011010000110001",
			3340 => "0000001001000000000001000100001100",
			3341 => "0000001111000000001010010100000100",
			3342 => "00000000000000000011010001111101",
			3343 => "0000001000000000000010011000000100",
			3344 => "11111111101010010011010001111101",
			3345 => "00000000000000000011010001111101",
			3346 => "0000000110000000001000010000010100",
			3347 => "0000001010000000000110011000000100",
			3348 => "00000000000000000011010001111101",
			3349 => "0000000110000000001011001100000100",
			3350 => "00000000000000000011010001111101",
			3351 => "0000001001000000001101011000001000",
			3352 => "0000001100000000000011011100000100",
			3353 => "00000000000000000011010001111101",
			3354 => "00000000110100100011010001111101",
			3355 => "00000000000000000011010001111101",
			3356 => "0000001010000000000001010000000100",
			3357 => "00000000000000000011010001111101",
			3358 => "11111111111111000011010001111101",
			3359 => "0000001001000000001101101000000100",
			3360 => "00000000000000000011010010110001",
			3361 => "0000000100000000001110111000000100",
			3362 => "00000000000000000011010010110001",
			3363 => "0000001001000000000101010000010000",
			3364 => "0000000100000000000100111000001100",
			3365 => "0000000011000000000010010100001000",
			3366 => "0000001011000000000101101100000100",
			3367 => "00000000000000000011010010110001",
			3368 => "00000000010001100011010010110001",
			3369 => "00000000000000000011010010110001",
			3370 => "00000000000000000011010010110001",
			3371 => "00000000000000000011010010110001",
			3372 => "0000000000000000000010111100011000",
			3373 => "0000001000000000001001101000000100",
			3374 => "00000000000000000011010011111101",
			3375 => "0000000001000000000101011100010000",
			3376 => "0000001101000000001001110100000100",
			3377 => "00000000000000000011010011111101",
			3378 => "0000001000000000001011010100001000",
			3379 => "0000000100000000001000000100000100",
			3380 => "00000000000000000011010011111101",
			3381 => "00000000101110100011010011111101",
			3382 => "00000000000000000011010011111101",
			3383 => "00000000000000000011010011111101",
			3384 => "0000000001000000001011101000001100",
			3385 => "0000000100000000001010010000001000",
			3386 => "0000001111000000000010110100000100",
			3387 => "00000000000000000011010011111101",
			3388 => "11111111100001000011010011111101",
			3389 => "00000000000000000011010011111101",
			3390 => "00000000000000000011010011111101",
			3391 => "0000000100000000000011101100001100",
			3392 => "0000000010000000000010011100000100",
			3393 => "00000000000000000011010101010001",
			3394 => "0000000111000000000111010000000100",
			3395 => "11111111010101100011010101010001",
			3396 => "00000000000000000011010101010001",
			3397 => "0000001000000000000010101000010100",
			3398 => "0000000001000000000000111100010000",
			3399 => "0000000000000000001011000100001100",
			3400 => "0000000001000000001100110100000100",
			3401 => "00000000000000000011010101010001",
			3402 => "0000001000000000001001101000000100",
			3403 => "00000000000000000011010101010001",
			3404 => "00000000011100110011010101010001",
			3405 => "00000000000000000011010101010001",
			3406 => "00000000000000000011010101010001",
			3407 => "0000000100000000001101000000000100",
			3408 => "11111111101111010011010101010001",
			3409 => "0000000100000000001111110000000100",
			3410 => "00000000000001010011010101010001",
			3411 => "00000000000000000011010101010001",
			3412 => "0000000100000000000011101100001100",
			3413 => "0000000010000000000010011100000100",
			3414 => "00000000000000000011010110100101",
			3415 => "0000000110000000001000010000000100",
			3416 => "11111111010000110011010110100101",
			3417 => "00000000000000000011010110100101",
			3418 => "0000000110000000000100111100011100",
			3419 => "0000001101000000000101100100010000",
			3420 => "0000001111000000001111010000001000",
			3421 => "0000000011000000001110001100000100",
			3422 => "00000000000000000011010110100101",
			3423 => "00000000000011100011010110100101",
			3424 => "0000001110000000001101010100000100",
			3425 => "00000000000000000011010110100101",
			3426 => "11111111111100000011010110100101",
			3427 => "0000001100000000000100001000001000",
			3428 => "0000001000000000001001101000000100",
			3429 => "00000000000000000011010110100101",
			3430 => "00000000100110100011010110100101",
			3431 => "00000000000000000011010110100101",
			3432 => "00000000000000000011010110100101",
			3433 => "0000001000000000000111000100011100",
			3434 => "0000001011000000000101101100000100",
			3435 => "00000000000000000011010111110001",
			3436 => "0000001000000000001001101000000100",
			3437 => "00000000000000000011010111110001",
			3438 => "0000000001000000000101011100010000",
			3439 => "0000001010000000001100011100001100",
			3440 => "0000001100000000000100000000000100",
			3441 => "00000000000000000011010111110001",
			3442 => "0000000100000000001000000100000100",
			3443 => "00000000000000000011010111110001",
			3444 => "00000000011001100011010111110001",
			3445 => "00000000000000000011010111110001",
			3446 => "00000000000000000011010111110001",
			3447 => "0000000100000000001010010000001000",
			3448 => "0000001011000000001000011000000100",
			3449 => "11111111101101110011010111110001",
			3450 => "00000000000000000011010111110001",
			3451 => "00000000000000000011010111110001",
			3452 => "0000000111000000001100101000011100",
			3453 => "0000001011000000000101101100000100",
			3454 => "00000000000000000011011000111101",
			3455 => "0000000001000000001111001100010100",
			3456 => "0000000000000000000010111100000100",
			3457 => "00000000000000000011011000111101",
			3458 => "0000000001000000000010001100000100",
			3459 => "00000000000000000011011000111101",
			3460 => "0000000010000000000010010100001000",
			3461 => "0000001100000000000100000000000100",
			3462 => "00000000000000000011011000111101",
			3463 => "00000000010101000011011000111101",
			3464 => "00000000000000000011011000111101",
			3465 => "00000000000000000011011000111101",
			3466 => "0000000000000000000010111100000100",
			3467 => "00000000000000000011011000111101",
			3468 => "0000000010000000001000100000000100",
			3469 => "00000000000000000011011000111101",
			3470 => "11111111100011100011011000111101",
			3471 => "0000001111000000000110010000011100",
			3472 => "0000000111000000001001110000000100",
			3473 => "00000000000000000011011010000001",
			3474 => "0000001000000000001001101000000100",
			3475 => "00000000000000000011011010000001",
			3476 => "0000001100000000001100110000010000",
			3477 => "0000000111000000001101111000001100",
			3478 => "0000001000000000001010000000001000",
			3479 => "0000001100000000000000101000000100",
			3480 => "00000000000000000011011010000001",
			3481 => "00000000010101000011011010000001",
			3482 => "00000000000000000011011010000001",
			3483 => "00000000000000000011011010000001",
			3484 => "00000000000000000011011010000001",
			3485 => "0000001100000000000011011100000100",
			3486 => "00000000000000000011011010000001",
			3487 => "11111111110100010011011010000001",
			3488 => "0000000111000000001100101000011100",
			3489 => "0000001101000000000100011000000100",
			3490 => "11111111101000000011011011010101",
			3491 => "0000000110000000001000010000010100",
			3492 => "0000000000000000000010111100000100",
			3493 => "00000000000000000011011011010101",
			3494 => "0000000001000000001100110100000100",
			3495 => "00000000000000000011011011010101",
			3496 => "0000001000000000001001101000000100",
			3497 => "00000000000000000011011011010101",
			3498 => "0000000111000000001001110000000100",
			3499 => "00000000000000000011011011010101",
			3500 => "00000000100101110011011011010101",
			3501 => "00000000000000000011011011010101",
			3502 => "0000001101000000001001010100001100",
			3503 => "0000001011000000001110110000000100",
			3504 => "00000000000000000011011011010101",
			3505 => "0000000010000000000000010000000100",
			3506 => "00000000000000000011011011010101",
			3507 => "11111111010110100011011011010101",
			3508 => "00000000000000000011011011010101",
			3509 => "0000001001000000001010011000100100",
			3510 => "0000000010000000001110010000011000",
			3511 => "0000000011000000000011100000000100",
			3512 => "00000000000000000011011100101001",
			3513 => "0000001110000000000011100000010000",
			3514 => "0000001011000000000101101100000100",
			3515 => "00000000000000000011011100101001",
			3516 => "0000001011000000001110001100001000",
			3517 => "0000001100000000001001110000000100",
			3518 => "00000000001100110011011100101001",
			3519 => "00000000000000000011011100101001",
			3520 => "00000000000000000011011100101001",
			3521 => "00000000000000000011011100101001",
			3522 => "0000000100000000001010010000001000",
			3523 => "0000001110000000001000111000000100",
			3524 => "00000000000000000011011100101001",
			3525 => "11111111011110010011011100101001",
			3526 => "00000000000000000011011100101001",
			3527 => "0000000001000000001001011000000100",
			3528 => "00000000001100010011011100101001",
			3529 => "00000000000000000011011100101001",
			3530 => "0000000010000000000110101100011100",
			3531 => "0000001001000000001101101000000100",
			3532 => "00000000000000000011011101111101",
			3533 => "0000000000000000000010111100000100",
			3534 => "00000000000000000011011101111101",
			3535 => "0000001011000000000101101100000100",
			3536 => "00000000000000000011011101111101",
			3537 => "0000000110000000001001100100001100",
			3538 => "0000000111000000001001110000000100",
			3539 => "00000000000000000011011101111101",
			3540 => "0000001101000000000100011000000100",
			3541 => "00000000000000000011011101111101",
			3542 => "00000000011100110011011101111101",
			3543 => "00000000000000000011011101111101",
			3544 => "0000001111000000001011110000001100",
			3545 => "0000000100000000001010010000001000",
			3546 => "0000000000000000000010111100000100",
			3547 => "00000000000000000011011101111101",
			3548 => "11111111011110000011011101111101",
			3549 => "00000000000000000011011101111101",
			3550 => "00000000000000000011011101111101",
			3551 => "0000000111000000000001111100011100",
			3552 => "0000001101000000000100011000000100",
			3553 => "00000000000000000011011110111001",
			3554 => "0000001010000000000110011100010100",
			3555 => "0000000000000000000010111100000100",
			3556 => "00000000000000000011011110111001",
			3557 => "0000000111000000001001110000000100",
			3558 => "00000000000000000011011110111001",
			3559 => "0000001111000000000000010000001000",
			3560 => "0000001000000000001001101000000100",
			3561 => "00000000000000000011011110111001",
			3562 => "00000000011101010011011110111001",
			3563 => "00000000000000000011011110111001",
			3564 => "00000000000000000011011110111001",
			3565 => "11111111110100010011011110111001",
			3566 => "0000000001000000000110101000000100",
			3567 => "00000000000000000011011111110101",
			3568 => "0000000001000000000101011100011000",
			3569 => "0000001010000000001001000100000100",
			3570 => "00000000000000000011011111110101",
			3571 => "0000000111000000001001110000000100",
			3572 => "00000000000000000011011111110101",
			3573 => "0000001101000000001001110100000100",
			3574 => "00000000000000000011011111110101",
			3575 => "0000001011000000001011110100001000",
			3576 => "0000000101000000001000000000000100",
			3577 => "00000000000000000011011111110101",
			3578 => "00000000010001010011011111110101",
			3579 => "00000000000000000011011111110101",
			3580 => "00000000000000000011011111110101",
			3581 => "0000001110000000001100101100000100",
			3582 => "00000000000000000011100000110001",
			3583 => "0000001111000000000000010000011000",
			3584 => "0000000001000000001101011100010100",
			3585 => "0000001010000000001001000100000100",
			3586 => "00000000000000000011100000110001",
			3587 => "0000001001000000001101101000000100",
			3588 => "00000000000000000011100000110001",
			3589 => "0000001001000000001101011000001000",
			3590 => "0000000110000000001000010000000100",
			3591 => "00000000010110100011100000110001",
			3592 => "00000000000000000011100000110001",
			3593 => "00000000000000000011100000110001",
			3594 => "00000000000000000011100000110001",
			3595 => "00000000000000000011100000110001",
			3596 => "0000000100000000001110111000000100",
			3597 => "11111111001111100011100010001101",
			3598 => "0000001000000000000111000100010000",
			3599 => "0000000111000000001001110000000100",
			3600 => "00000000000000000011100010001101",
			3601 => "0000000010000000000011110000001000",
			3602 => "0000001000000000001001101000000100",
			3603 => "00000000000000000011100010001101",
			3604 => "00000000010011000011100010001101",
			3605 => "00000000000000000011100010001101",
			3606 => "0000000110000000000100111100010100",
			3607 => "0000000100000000000110110000001000",
			3608 => "0000000010000000001100111000000100",
			3609 => "11111111111111100011100010001101",
			3610 => "00000000000000000011100010001101",
			3611 => "0000000110000000001011001100000100",
			3612 => "00000000000000000011100010001101",
			3613 => "0000000000000000000110100100000100",
			3614 => "00000000011011100011100010001101",
			3615 => "00000000000000000011100010001101",
			3616 => "0000001101000000001100100100000100",
			3617 => "11111111100010000011100010001101",
			3618 => "00000000000000000011100010001101",
			3619 => "0000000010000000000110101100011100",
			3620 => "0000001001000000001101101000000100",
			3621 => "00000000000000000011100011101001",
			3622 => "0000000000000000000010111100000100",
			3623 => "00000000000000000011100011101001",
			3624 => "0000001011000000000101101100000100",
			3625 => "00000000000000000011100011101001",
			3626 => "0000000110000000001001100100001100",
			3627 => "0000001000000000001001101000000100",
			3628 => "00000000000000000011100011101001",
			3629 => "0000000111000000001001110000000100",
			3630 => "00000000000000000011100011101001",
			3631 => "00000000011000010011100011101001",
			3632 => "00000000000000000011100011101001",
			3633 => "0000001100000000001100110000000100",
			3634 => "00000000000000000011100011101001",
			3635 => "0000001111000000001011110000001100",
			3636 => "0000000000000000000010111100000100",
			3637 => "00000000000000000011100011101001",
			3638 => "0000000000000000001010111100000100",
			3639 => "11111111011110100011100011101001",
			3640 => "00000000000000000011100011101001",
			3641 => "00000000000000000011100011101001",
			3642 => "0000000000000000000010111100011000",
			3643 => "0000001000000000001001101000000100",
			3644 => "11111111110100100011100101011101",
			3645 => "0000001100000000001000111000000100",
			3646 => "00000000000000000011100101011101",
			3647 => "0000000001000000000101011100001100",
			3648 => "0000001000000000001011010100001000",
			3649 => "0000000100000000001000000100000100",
			3650 => "00000000000000000011100101011101",
			3651 => "00000001010011010011100101011101",
			3652 => "00000000000000000011100101011101",
			3653 => "00000000000000000011100101011101",
			3654 => "0000000010000000000100101000001000",
			3655 => "0000000011000000001010111000000100",
			3656 => "11111111111001010011100101011101",
			3657 => "00000000111001110011100101011101",
			3658 => "0000000100000000001011001000000100",
			3659 => "11111110111110000011100101011101",
			3660 => "0000000010000000000110101100001100",
			3661 => "0000000101000000001001001000000100",
			3662 => "00000000000000000011100101011101",
			3663 => "0000001110000000001101100000000100",
			3664 => "00000000000000000011100101011101",
			3665 => "00000000011011110011100101011101",
			3666 => "0000000000000000001010111100001000",
			3667 => "0000000101000000001011011100000100",
			3668 => "11111111010001000011100101011101",
			3669 => "00000000000000000011100101011101",
			3670 => "00000000000000000011100101011101",
			3671 => "0000000000000000000010111100011000",
			3672 => "0000001000000000001001101000000100",
			3673 => "11111111110110010011100111010001",
			3674 => "0000001100000000001000111000000100",
			3675 => "00000000000000000011100111010001",
			3676 => "0000000001000000000101011100001100",
			3677 => "0000001000000000001011010100001000",
			3678 => "0000000100000000001000000100000100",
			3679 => "00000000000000000011100111010001",
			3680 => "00000001001110110011100111010001",
			3681 => "00000000000000000011100111010001",
			3682 => "00000000000000000011100111010001",
			3683 => "0000000010000000000100101000001000",
			3684 => "0000000011000000001010111000000100",
			3685 => "11111111111010100011100111010001",
			3686 => "00000000110111000011100111010001",
			3687 => "0000000100000000001011001000000100",
			3688 => "11111111000001000011100111010001",
			3689 => "0000000010000000000110101100001000",
			3690 => "0000000001000000000110101000000100",
			3691 => "00000000000000000011100111010001",
			3692 => "00000000011100000011100111010001",
			3693 => "0000000000000000001010111100001100",
			3694 => "0000000101000000001011011100001000",
			3695 => "0000001111000000001110101000000100",
			3696 => "00000000000000000011100111010001",
			3697 => "11111111010101010011100111010001",
			3698 => "00000000000000000011100111010001",
			3699 => "00000000000000000011100111010001",
			3700 => "0000000010000000000100101000010000",
			3701 => "0000000111000000001001110000000100",
			3702 => "00000000000000000011101001010101",
			3703 => "0000001110000000001001110000000100",
			3704 => "00000000000000000011101001010101",
			3705 => "0000001000000000001001101000000100",
			3706 => "00000000000000000011101001010101",
			3707 => "00000000111110010011101001010101",
			3708 => "0000000000000000000010111100011000",
			3709 => "0000001010000000000110011000000100",
			3710 => "00000000000000000011101001010101",
			3711 => "0000000001000000000101011100010000",
			3712 => "0000000011000000000101110100000100",
			3713 => "00000000000000000011101001010101",
			3714 => "0000001000000000001011010100001000",
			3715 => "0000000100000000001000000100000100",
			3716 => "00000000000000000011101001010101",
			3717 => "00000000101011010011101001010101",
			3718 => "00000000000000000011101001010101",
			3719 => "00000000000000000011101001010101",
			3720 => "0000000100000000001101000000001100",
			3721 => "0000001011000000000100011000001000",
			3722 => "0000000010000000000111111100000100",
			3723 => "00000000000000000011101001010101",
			3724 => "11111111001100100011101001010101",
			3725 => "00000000000000000011101001010101",
			3726 => "0000001010000000000111000100001100",
			3727 => "0000001011000000001001110100001000",
			3728 => "0000000110000000001010011000000100",
			3729 => "00000000000000000011101001010101",
			3730 => "00000000011110010011101001010101",
			3731 => "00000000000000000011101001010101",
			3732 => "11111111111111100011101001010101",
			3733 => "0000000100000000001110111000000100",
			3734 => "11111111001010110011101010111001",
			3735 => "0000001000000000000111000100011000",
			3736 => "0000000001000000000101011100010100",
			3737 => "0000000001000000001100110100000100",
			3738 => "00000000000000000011101010111001",
			3739 => "0000001010000000001100011100001100",
			3740 => "0000001010000000000110011000000100",
			3741 => "00000000000000000011101010111001",
			3742 => "0000001101000000000100011000000100",
			3743 => "00000000000000000011101010111001",
			3744 => "00000000100011000011101010111001",
			3745 => "00000000000000000011101010111001",
			3746 => "00000000000000000011101010111001",
			3747 => "0000000110000000000100111100010000",
			3748 => "0000000110000000001011001100000100",
			3749 => "00000000000000000011101010111001",
			3750 => "0000000100000000000110110000000100",
			3751 => "00000000000000000011101010111001",
			3752 => "0000000001000000000010001100000100",
			3753 => "00000000000000000011101010111001",
			3754 => "00000000011111100011101010111001",
			3755 => "0000001101000000001100100100000100",
			3756 => "11111111011110110011101010111001",
			3757 => "00000000000000000011101010111001",
			3758 => "0000001111000000000110010000110100",
			3759 => "0000000111000000001001110000001000",
			3760 => "0000001010000000000110001000000100",
			3761 => "11111111010111100011101100111101",
			3762 => "00000000000000000011101100111101",
			3763 => "0000000111000000001101100000010100",
			3764 => "0000000010000000000110010000010000",
			3765 => "0000001010000000000110011000000100",
			3766 => "00000000000000000011101100111101",
			3767 => "0000001101000000000100011000000100",
			3768 => "00000000000000000011101100111101",
			3769 => "0000000110000000001011001100000100",
			3770 => "00000000111111010011101100111101",
			3771 => "00000000000000000011101100111101",
			3772 => "00000000000000000011101100111101",
			3773 => "0000000100000000001011001000001000",
			3774 => "0000000010000000001010001000000100",
			3775 => "00000000000000000011101100111101",
			3776 => "11111111100111110011101100111101",
			3777 => "0000000001000000001001111000000100",
			3778 => "00000000000000000011101100111101",
			3779 => "0000000110000000001101011000000100",
			3780 => "00000000000000000011101100111101",
			3781 => "0000000111000000000111001000000100",
			3782 => "00000000100100110011101100111101",
			3783 => "00000000000000000011101100111101",
			3784 => "0000001001000000001010011000001000",
			3785 => "0000001111000000001001100000000100",
			3786 => "00000000000000000011101100111101",
			3787 => "11111111000101010011101100111101",
			3788 => "0000000001000000001001011000000100",
			3789 => "00000000010101100011101100111101",
			3790 => "11111111100111000011101100111101",
			3791 => "0000000001000000001011101000011100",
			3792 => "0000001111000000000100101000011000",
			3793 => "0000001101000000000100011000000100",
			3794 => "00000000000000000011101110101001",
			3795 => "0000001100000000000110000100010000",
			3796 => "0000001010000000000110011000000100",
			3797 => "00000000000000000011101110101001",
			3798 => "0000000110000000001111000000001000",
			3799 => "0000000011000000001110001100000100",
			3800 => "00000000000000000011101110101001",
			3801 => "00000000011111110011101110101001",
			3802 => "00000000000000000011101110101001",
			3803 => "00000000000000000011101110101001",
			3804 => "11111111101100100011101110101001",
			3805 => "0000001010000000000110011000000100",
			3806 => "00000000000000000011101110101001",
			3807 => "0000000001000000000101011100010100",
			3808 => "0000001101000000001011011100000100",
			3809 => "00000000000000000011101110101001",
			3810 => "0000000010000000000011110000001100",
			3811 => "0000000110000000000101010000001000",
			3812 => "0000000100000000000000010100000100",
			3813 => "00000000000000000011101110101001",
			3814 => "00000000100111100011101110101001",
			3815 => "00000000000000000011101110101001",
			3816 => "00000000000000000011101110101001",
			3817 => "00000000000000000011101110101001",
			3818 => "0000000101000000000100011000001000",
			3819 => "0000000100000000001101000000000100",
			3820 => "11111110111011110011110000011101",
			3821 => "00000000000000000011110000011101",
			3822 => "0000001100000000000011011100010000",
			3823 => "0000001100000000001000111000000100",
			3824 => "00000000000000000011110000011101",
			3825 => "0000001111000000000000010000001000",
			3826 => "0000001000000000001001101000000100",
			3827 => "00000000000000000011110000011101",
			3828 => "00000001001111000011110000011101",
			3829 => "00000000000000000011110000011101",
			3830 => "0000001010000000000110011000000100",
			3831 => "11111111100101110011110000011101",
			3832 => "0000000111000000001101111000010000",
			3833 => "0000001010000000001100000100001100",
			3834 => "0000000110000000001101011000000100",
			3835 => "00000000000000000011110000011101",
			3836 => "0000001001000000000001111000000100",
			3837 => "11111111100111000011110000011101",
			3838 => "00000000000000000011110000011101",
			3839 => "00000000000000000011110000011101",
			3840 => "0000000011000000001111101000001100",
			3841 => "0000000110000000001101011000000100",
			3842 => "00000000000000000011110000011101",
			3843 => "0000001001000000000001000100000100",
			3844 => "00000000000000000011110000011101",
			3845 => "00000000100011110011110000011101",
			3846 => "00000000000000000011110000011101",
			3847 => "0000001101000000000100011000000100",
			3848 => "11111110011011000011110010000001",
			3849 => "0000001100000000000100001000100000",
			3850 => "0000000110000000001000010000011100",
			3851 => "0000000000000000000010011000000100",
			3852 => "11111110110000000011110010000001",
			3853 => "0000000010000000001110010000001000",
			3854 => "0000001011000000001110001100000100",
			3855 => "00000011010101010011110010000001",
			3856 => "11111111001001110011110010000001",
			3857 => "0000001011000000001110001100001000",
			3858 => "0000000011000000000011100000000100",
			3859 => "00000000101110100011110010000001",
			3860 => "11111110100100010011110010000001",
			3861 => "0000001100000000001100110000000100",
			3862 => "00000001100110110011110010000001",
			3863 => "00000000011110100011110010000001",
			3864 => "11111110011011110011110010000001",
			3865 => "0000000010000000000101000000000100",
			3866 => "11111110011110000011110010000001",
			3867 => "0000001111000000000101000000001000",
			3868 => "0000000000000000000010111100000100",
			3869 => "00000001010001010011110010000001",
			3870 => "11111111111100010011110010000001",
			3871 => "11111110100110100011110010000001",
			3872 => "0000001101000000000100011000000100",
			3873 => "11111110110101010011110011111101",
			3874 => "0000000111000000001100101000101100",
			3875 => "0000001000000000000111000100010100",
			3876 => "0000000000000000000010111100000100",
			3877 => "00000000000000000011110011111101",
			3878 => "0000000111000000001001110000000100",
			3879 => "00000000000000000011110011111101",
			3880 => "0000001100000000001110001100001000",
			3881 => "0000001110000000001110010000000100",
			3882 => "00000001010110010011110011111101",
			3883 => "00000000000000000011110011111101",
			3884 => "00000000000000000011110011111101",
			3885 => "0000000100000000001101000000001100",
			3886 => "0000001100000000000011011100001000",
			3887 => "0000000110000000001101011000000100",
			3888 => "00000000000000000011110011111101",
			3889 => "11111111010010110011110011111101",
			3890 => "00000000000000000011110011111101",
			3891 => "0000000110000000001101011000000100",
			3892 => "00000000000000000011110011111101",
			3893 => "0000000000000000000001001000000100",
			3894 => "00000000101000100011110011111101",
			3895 => "00000000000000000011110011111101",
			3896 => "0000000010000000001000100000001000",
			3897 => "0000001100000000001110001100000100",
			3898 => "00000000000000000011110011111101",
			3899 => "11111111111101110011110011111101",
			3900 => "0000001110000000001010111000000100",
			3901 => "00000000000000000011110011111101",
			3902 => "11111111001101100011110011111101",
			3903 => "0000000101000000000100011000001000",
			3904 => "0000000100000000001101000000000100",
			3905 => "11111110110111110011110110001001",
			3906 => "00000000000000000011110110001001",
			3907 => "0000000010000000000110010000010000",
			3908 => "0000001011000000001110001100001100",
			3909 => "0000001100000000000011011100001000",
			3910 => "0000000000000000000010111100000100",
			3911 => "00000000000000000011110110001001",
			3912 => "00000001100001100011110110001001",
			3913 => "00000000000000000011110110001001",
			3914 => "00000000000000000011110110001001",
			3915 => "0000000111000000001101111000010000",
			3916 => "0000000000000000001100101100001100",
			3917 => "0000001111000000001101000100000100",
			3918 => "00000000000000000011110110001001",
			3919 => "0000001001000000000001111000000100",
			3920 => "11111111010001000011110110001001",
			3921 => "00000000000000000011110110001001",
			3922 => "00000000000000000011110110001001",
			3923 => "0000000100000000001100111100010000",
			3924 => "0000000010000000001110100100001000",
			3925 => "0000000010000000001011111000000100",
			3926 => "00000000000000000011110110001001",
			3927 => "11111111011011010011110110001001",
			3928 => "0000000011000000001111101000000100",
			3929 => "00000000100010000011110110001001",
			3930 => "00000000000000000011110110001001",
			3931 => "0000000111000000000111001000001100",
			3932 => "0000000110000000001101011000000100",
			3933 => "00000000000000000011110110001001",
			3934 => "0000001000000000000110001000000100",
			3935 => "00000000000000000011110110001001",
			3936 => "00000000111111000011110110001001",
			3937 => "00000000000000000011110110001001",
			3938 => "0000000110000000001101011000011100",
			3939 => "0000001001000000001011101000001000",
			3940 => "0000001111000000000101110000000100",
			3941 => "11111110011001100011111000111101",
			3942 => "11111100110011110011111000111101",
			3943 => "0000001111000000000010110100001100",
			3944 => "0000001000000000001001101000000100",
			3945 => "11111110011111010011111000111101",
			3946 => "0000000101000000000011100000000100",
			3947 => "11111110101111100011111000111101",
			3948 => "00000101010001010011111000111101",
			3949 => "0000000011000000001110110000000100",
			3950 => "00000000110100010011111000111101",
			3951 => "11111110010101010011111000111101",
			3952 => "0000001100000000000100001000110000",
			3953 => "0000000010000000000000010000010100",
			3954 => "0000001011000000001110001100000100",
			3955 => "11111110011100110011111000111101",
			3956 => "0000000111000000001001110000000100",
			3957 => "00001000000010110011111000111101",
			3958 => "0000000000000000001100110000000100",
			3959 => "11111110100101010011111000111101",
			3960 => "0000001110000000000110001000000100",
			3961 => "11111111000101010011111000111101",
			3962 => "00000001010110100011111000111101",
			3963 => "0000000110000000001000010000011000",
			3964 => "0000001111000000001010000100010000",
			3965 => "0000001111000000000110010000001000",
			3966 => "0000001110000000000100010000000100",
			3967 => "00000001101011100011111000111101",
			3968 => "00000011101000010011111000111101",
			3969 => "0000001001000000000100111100000100",
			3970 => "00000000001000100011111000111101",
			3971 => "11111110100011010011111000111101",
			3972 => "0000000000000000000010111100000100",
			3973 => "00000000000000000011111000111101",
			3974 => "00000100000000110011111000111101",
			3975 => "11111110001010110011111000111101",
			3976 => "0000001110000000001101101100001100",
			3977 => "0000000011000000000011000000000100",
			3978 => "11111110011011010011111000111101",
			3979 => "0000000011000000001111101000000100",
			3980 => "00000010100101100011111000111101",
			3981 => "11111110111010110011111000111101",
			3982 => "11111110011001100011111000111101",
			3983 => "0000001101000000000100011000000100",
			3984 => "11111110110111100011111011000001",
			3985 => "0000000111000000001100101000110000",
			3986 => "0000001000000000000111000100011000",
			3987 => "0000000000000000000010111100000100",
			3988 => "00000000000000000011111011000001",
			3989 => "0000000111000000001001110000000100",
			3990 => "00000000000000000011111011000001",
			3991 => "0000000111000000001101100000001000",
			3992 => "0000000110000000001011001100000100",
			3993 => "00000001101000010011111011000001",
			3994 => "00000000000000000011111011000001",
			3995 => "0000000011000000000010110100000100",
			3996 => "11111111111110100011111011000001",
			3997 => "00000000111010100011111011000001",
			3998 => "0000000001000000000110101000001100",
			3999 => "0000001111000000001110101000000100",
			4000 => "00000000000000000011111011000001",
			4001 => "0000000000000000001100101100000100",
			4002 => "11111111001010010011111011000001",
			4003 => "00000000000000000011111011000001",
			4004 => "0000000000000000000100000000000100",
			4005 => "00000000000000000011111011000001",
			4006 => "0000001010000000000110001000000100",
			4007 => "00000000011111110011111011000001",
			4008 => "00000000000000000011111011000001",
			4009 => "0000000010000000001000100000001000",
			4010 => "0000001100000000001110001100000100",
			4011 => "00000000000000000011111011000001",
			4012 => "11111111111111100011111011000001",
			4013 => "0000001011000000001110110000000100",
			4014 => "00000000000000000011111011000001",
			4015 => "11111111001110110011111011000001",
			4016 => "0000001001000000001101101000000100",
			4017 => "11111111001011100011111100111101",
			4018 => "0000000010000000000110010000011000",
			4019 => "0000001011000000000101101100000100",
			4020 => "00000000000000000011111100111101",
			4021 => "0000001100000000001100110000010000",
			4022 => "0000001000000000001001101000000100",
			4023 => "00000000000000000011111100111101",
			4024 => "0000000111000000001001110000000100",
			4025 => "00000000000000000011111100111101",
			4026 => "0000000110000000001011001100000100",
			4027 => "00000001000111110011111100111101",
			4028 => "00000000000000000011111100111101",
			4029 => "00000000000000000011111100111101",
			4030 => "0000000001000000001011101000001000",
			4031 => "0000001110000000001010001100000100",
			4032 => "00000000000000000011111100111101",
			4033 => "11111111000110000011111100111101",
			4034 => "0000001101000000001011011100001000",
			4035 => "0000000110000000001111000000000100",
			4036 => "11111111111011000011111100111101",
			4037 => "00000000000000000011111100111101",
			4038 => "0000001100000000000100001000001100",
			4039 => "0000001000000000001011010100000100",
			4040 => "00000000000000000011111100111101",
			4041 => "0000000001000000000000111100000100",
			4042 => "00000000110110010011111100111101",
			4043 => "00000000000000000011111100111101",
			4044 => "0000000110000000001000010000000100",
			4045 => "11111111111011010011111100111101",
			4046 => "00000000000000000011111100111101",
			4047 => "0000000100000000001001000000100100",
			4048 => "0000000100000000001110111000000100",
			4049 => "11111110011000110011111111110001",
			4050 => "0000001000000000000110001000010100",
			4051 => "0000000000000000000011010000001100",
			4052 => "0000000001000000000101011100001000",
			4053 => "0000000111000000001101010100000100",
			4054 => "11111110110111000011111111110001",
			4055 => "00000010010101100011111111110001",
			4056 => "11111110100000000011111111110001",
			4057 => "0000001110000000001011000100000100",
			4058 => "11111111011101100011111111110001",
			4059 => "00000110100001100011111111110001",
			4060 => "0000001011000000000101101100000100",
			4061 => "11111110011001010011111111110001",
			4062 => "0000000101000000001010111000000100",
			4063 => "00000010010110110011111111110001",
			4064 => "11111110011111000011111111110001",
			4065 => "0000001001000000001011101000010000",
			4066 => "0000001111000000000101001000001100",
			4067 => "0000001001000000001101101000000100",
			4068 => "11111110011001010011111111110001",
			4069 => "0000001110000000000110000100000100",
			4070 => "00000001001100100011111111110001",
			4071 => "11111111001101010011111111110001",
			4072 => "11111101001001010011111111110001",
			4073 => "0000000111000000000011100000100100",
			4074 => "0000000000000000001100001000010100",
			4075 => "0000001000000000001011010100001000",
			4076 => "0000000111000000001101010100000100",
			4077 => "11111110011101100011111111110001",
			4078 => "00000011000110010011111111110001",
			4079 => "0000001000000000000010101000001000",
			4080 => "0000000010000000001011111000000100",
			4081 => "00000101110110000011111111110001",
			4082 => "00000010100100000011111111110001",
			4083 => "00000000000000000011111111110001",
			4084 => "0000000000000000001000111100000100",
			4085 => "11111111011001010011111111110001",
			4086 => "0000000100000000001011100100000100",
			4087 => "11111110110110100011111111110001",
			4088 => "0000001010000000000001110000000100",
			4089 => "00000000111110100011111111110001",
			4090 => "00000001110100010011111111110001",
			4091 => "11111110011001110011111111110001",
			4092 => "0000001101000000000100011000000100",
			4093 => "11111110100110000100000001110101",
			4094 => "0000001111000000000010110100010000",
			4095 => "0000001111000000001011011100000100",
			4096 => "00000000000000000100000001110101",
			4097 => "0000000100000000000010111000000100",
			4098 => "00000000000000000100000001110101",
			4099 => "0000001100000000000110000100000100",
			4100 => "00000001101000100100000001110101",
			4101 => "00000000000000000100000001110101",
			4102 => "0000000001000000001011101000001100",
			4103 => "0000000100000000001010010000000100",
			4104 => "11111110111110000100000001110101",
			4105 => "0000000101000000001011011100000100",
			4106 => "00000000011001110100000001110101",
			4107 => "00000000000000000100000001110101",
			4108 => "0000000111000000001100101000001100",
			4109 => "0000001011000000001010111000000100",
			4110 => "00000000000000000100000001110101",
			4111 => "0000001000000000001011010100000100",
			4112 => "00000000000000000100000001110101",
			4113 => "00000001011111100100000001110101",
			4114 => "0000000101000000000101100100001100",
			4115 => "0000000010000000001100111000001000",
			4116 => "0000001100000000001110001100000100",
			4117 => "11111110110011100100000001110101",
			4118 => "00000000000000000100000001110101",
			4119 => "00000000000000000100000001110101",
			4120 => "0000001100000000001010111000001000",
			4121 => "0000001010000000000001010000000100",
			4122 => "00000000000000000100000001110101",
			4123 => "00000000101110000100000001110101",
			4124 => "11111111000100010100000001110101",
			4125 => "0000000111000000001001110000001000",
			4126 => "0000001010000000000110001000000100",
			4127 => "11111110111010010100000100001001",
			4128 => "00000000000000000100000100001001",
			4129 => "0000000010000000000111111100010000",
			4130 => "0000000010000000001001010000000100",
			4131 => "00000000000000000100000100001001",
			4132 => "0000000100000000000010111000000100",
			4133 => "00000000000000000100000100001001",
			4134 => "0000000111000000001110001100000100",
			4135 => "00000001000110010100000100001001",
			4136 => "00000000000000000100000100001001",
			4137 => "0000000100000000001011001000001100",
			4138 => "0000000010000000001110100100000100",
			4139 => "11111111000001000100000100001001",
			4140 => "0000000011000000001111101000000100",
			4141 => "00000000011001100100000100001001",
			4142 => "00000000000000000100000100001001",
			4143 => "0000000000000000001100001000010000",
			4144 => "0000000011000000001001011100001100",
			4145 => "0000000111000000001010111100001000",
			4146 => "0000001100000000001101111000000100",
			4147 => "00000000111110000100000100001001",
			4148 => "00000000000000000100000100001001",
			4149 => "00000000000000000100000100001001",
			4150 => "00000000000000000100000100001001",
			4151 => "0000000100000000001101000000001000",
			4152 => "0000001001000000000100110100000100",
			4153 => "11111111001000010100000100001001",
			4154 => "00000000000000000100000100001001",
			4155 => "0000001110000000001110110000001000",
			4156 => "0000001100000000000110000100000100",
			4157 => "00000000000000000100000100001001",
			4158 => "11111111101000100100000100001001",
			4159 => "0000000011000000001100010000000100",
			4160 => "00000000011000100100000100001001",
			4161 => "00000000000000000100000100001001",
			4162 => "0000000100000000001001000000100000",
			4163 => "0000000100000000001110111000000100",
			4164 => "11111110011000100100000110111101",
			4165 => "0000001000000000000110001000010000",
			4166 => "0000000011000000000010010100001100",
			4167 => "0000001000000000001011010100001000",
			4168 => "0000001100000000000000001100000100",
			4169 => "11111110101010100100000110111101",
			4170 => "00000010001101010100000110111101",
			4171 => "00000111111000110100000110111101",
			4172 => "11111110100100110100000110111101",
			4173 => "0000001101000000000100011000000100",
			4174 => "11111110011000110100000110111101",
			4175 => "0000000011000000001001001000000100",
			4176 => "00000011110111000100000110111101",
			4177 => "11111110011101110100000110111101",
			4178 => "0000001001000000001011101000010000",
			4179 => "0000001111000000000101001000001100",
			4180 => "0000001001000000001101101000000100",
			4181 => "11111110011000110100000110111101",
			4182 => "0000001110000000000110000100000100",
			4183 => "00000001011000100100000110111101",
			4184 => "11111111000111100100000110111101",
			4185 => "11111100101101010100000110111101",
			4186 => "0000000110000000001000010000101000",
			4187 => "0000000100000000000001001100010100",
			4188 => "0000000011000000001000011000000100",
			4189 => "00001110100110100100000110111101",
			4190 => "0000000011000000001101000100001000",
			4191 => "0000000001000000001101011100000100",
			4192 => "00000011111010010100000110111101",
			4193 => "11111110100011000100000110111101",
			4194 => "0000000101000000001011011100000100",
			4195 => "00100011100000100100000110111101",
			4196 => "00000101010000110100000110111101",
			4197 => "0000000110000000001101011000001000",
			4198 => "0000000010000000001011111000000100",
			4199 => "00000001101111010100000110111101",
			4200 => "11111110111000110100000110111101",
			4201 => "0000001111000000001100010100001000",
			4202 => "0000001010000000000001110000000100",
			4203 => "00000001011000100100000110111101",
			4204 => "00000001111011010100000110111101",
			4205 => "00000010111111000100000110111101",
			4206 => "11111110011000110100000110111101",
			4207 => "0000000100000000001001000000110000",
			4208 => "0000001011000000000101101100000100",
			4209 => "11111110011001110100001001011001",
			4210 => "0000001101000000000110100100011000",
			4211 => "0000001101000000001001110100001000",
			4212 => "0000001001000000001011101000000100",
			4213 => "00000010110000000100001001011001",
			4214 => "11111110100010110100001001011001",
			4215 => "0000000000000000000010111100000100",
			4216 => "11111111011001010100001001011001",
			4217 => "0000000000000000000011111100000100",
			4218 => "00011000111010010100001001011001",
			4219 => "0000000111000000001101100000000100",
			4220 => "00000000000000000100001001011001",
			4221 => "00000100000011100100001001011001",
			4222 => "0000000100000000000000010100000100",
			4223 => "11111110011010010100001001011001",
			4224 => "0000000000000000000010011000001100",
			4225 => "0000000001000000001011111100001000",
			4226 => "0000001000000000001100000100000100",
			4227 => "00000000000000000100001001011001",
			4228 => "00000010000000100100001001011001",
			4229 => "11111111111111000100001001011001",
			4230 => "11111110100110110100001001011001",
			4231 => "0000000001000000001100110100000100",
			4232 => "11111110011011000100001001011001",
			4233 => "0000000111000000001110110000011000",
			4234 => "0000000110000000001000010000010100",
			4235 => "0000000111000000001001110000001000",
			4236 => "0000001100000000000100000000000100",
			4237 => "11111110101011000100001001011001",
			4238 => "00000000000000000100001001011001",
			4239 => "0000000010000000001110110100000100",
			4240 => "00000011101000110100001001011001",
			4241 => "0000000110000000001101011000000100",
			4242 => "00000000000000000100001001011001",
			4243 => "00000001100000000100001001011001",
			4244 => "11111110010111010100001001011001",
			4245 => "11111110010110000100001001011001",
			4246 => "0000000100000000001001000000011100",
			4247 => "0000000100000000001110111000000100",
			4248 => "11111110011000100100001100000101",
			4249 => "0000001011000000000101101100000100",
			4250 => "11111110011001000100001100000101",
			4251 => "0000000010000000001100010100000100",
			4252 => "00000111001111110100001100000101",
			4253 => "0000001010000000001010110000001100",
			4254 => "0000000010000000001111100100000100",
			4255 => "11111110101100000100001100000101",
			4256 => "0000000011000000000010010100000100",
			4257 => "00000011010011100100001100000101",
			4258 => "11111110110110010100001100000101",
			4259 => "11111110011101000100001100000101",
			4260 => "0000001001000000001011101000010000",
			4261 => "0000001111000000000101001000001100",
			4262 => "0000001001000000001101101000000100",
			4263 => "11111110011001000100001100000101",
			4264 => "0000000010000000000111011000000100",
			4265 => "11111111001011010100001100000101",
			4266 => "00000001010010000100001100000101",
			4267 => "11111100111100110100001100000101",
			4268 => "0000000110000000001000010000101000",
			4269 => "0000000000000000001100001000011000",
			4270 => "0000000000000000000011010000001000",
			4271 => "0000001111000000000110010000000100",
			4272 => "11111110101101110100001100000101",
			4273 => "00000001110011000100001100000101",
			4274 => "0000000011000000000110100000001000",
			4275 => "0000001110000000001001001000000100",
			4276 => "00000111100011000100001100000101",
			4277 => "00000010011000100100001100000101",
			4278 => "0000000101000000000110110100000100",
			4279 => "00010000001001110100001100000101",
			4280 => "00000010111110110100001100000101",
			4281 => "0000000110000000001101011000000100",
			4282 => "00000000001000000100001100000101",
			4283 => "0000000100000000001101000000000100",
			4284 => "00000000011011010100001100000101",
			4285 => "0000001111000000001100010100000100",
			4286 => "00000001110100100100001100000101",
			4287 => "00000010101011010100001100000101",
			4288 => "11111110011001010100001100000101",
			4289 => "0000000111000000001001110000001000",
			4290 => "0000000010000000001000100000000100",
			4291 => "11111110101001100100001110100001",
			4292 => "00000000000000000100001110100001",
			4293 => "0000000111000000001001110000001100",
			4294 => "0000000010000000000110010000001000",
			4295 => "0000001101000000000100011000000100",
			4296 => "00000000000000000100001110100001",
			4297 => "00000001110011000100001110100001",
			4298 => "00000000000000000100001110100001",
			4299 => "0000001000000000000111000100010100",
			4300 => "0000000100000000000010111000000100",
			4301 => "11111110111111100100001110100001",
			4302 => "0000000001000000000101011100001100",
			4303 => "0000000001000000001001111000000100",
			4304 => "00000000000000000100001110100001",
			4305 => "0000001100000000001000111000000100",
			4306 => "00000000000000000100001110100001",
			4307 => "00000000111000010100001110100001",
			4308 => "00000000000000000100001110100001",
			4309 => "0000001111000000000101110000011000",
			4310 => "0000001110000000001100101100001100",
			4311 => "0000000010000000001111100100001000",
			4312 => "0000001100000000001000111000000100",
			4313 => "00000000000000000100001110100001",
			4314 => "11111111100110010100001110100001",
			4315 => "00000000000000000100001110100001",
			4316 => "0000000100000000000001100100000100",
			4317 => "00000000000000000100001110100001",
			4318 => "0000001100000000001000111000000100",
			4319 => "00000000000000000100001110100001",
			4320 => "00000000100110100100001110100001",
			4321 => "0000000010000000001000100000000100",
			4322 => "00000000000000000100001110100001",
			4323 => "0000001101000000001011110100000100",
			4324 => "11111110110001010100001110100001",
			4325 => "0000000011000000001001011100000100",
			4326 => "00000000000000000100001110100001",
			4327 => "11111111111011000100001110100001",
			4328 => "0000001101000000000100011000000100",
			4329 => "11111110011010100100010000111101",
			4330 => "0000001100000000001110001100011100",
			4331 => "0000000000000000000010111100000100",
			4332 => "11111110101100100100010000111101",
			4333 => "0000000000000000000010111100001000",
			4334 => "0000001000000000001011010100000100",
			4335 => "00000101001011010100010000111101",
			4336 => "00000000000000000100010000111101",
			4337 => "0000000100000000000100001100000100",
			4338 => "11111110101010000100010000111101",
			4339 => "0000000101000000000111001000000100",
			4340 => "00000011100100010100010000111101",
			4341 => "0000000100000000001011001000000100",
			4342 => "11111111011100010100010000111101",
			4343 => "00000001000101010100010000111101",
			4344 => "0000001100000000000100001000011100",
			4345 => "0000001101000000001110101100010100",
			4346 => "0000001101000000001011110100001100",
			4347 => "0000000111000000001100101000001000",
			4348 => "0000000111000000001100101000000100",
			4349 => "11111111011010110100010000111101",
			4350 => "00000000000000000100010000111101",
			4351 => "11111110100101100100010000111101",
			4352 => "0000000001000000001001011000000100",
			4353 => "00000000111010100100010000111101",
			4354 => "11111110110010100100010000111101",
			4355 => "0000000100000000001010110100000100",
			4356 => "00000000000000000100010000111101",
			4357 => "00000001101101010100010000111101",
			4358 => "0000000010000000000101000000000100",
			4359 => "11111110011010000100010000111101",
			4360 => "0000001100000000001010111000000100",
			4361 => "00000001001101100100010000111101",
			4362 => "0000000010000000000101000000001000",
			4363 => "0000001100000000001001110100000100",
			4364 => "00000000011011100100010000111101",
			4365 => "00000000000000000100010000111101",
			4366 => "11111110100001110100010000111101",
			4367 => "0000001101000000000100011000000100",
			4368 => "11111110100101000100010011100001",
			4369 => "0000000010000000000110010000011000",
			4370 => "0000000101000000001001001000010000",
			4371 => "0000001000000000000111000100001100",
			4372 => "0000000000000000000010111100000100",
			4373 => "00000000000000000100010011100001",
			4374 => "0000001100000000000011011100000100",
			4375 => "00000001111000010100010011100001",
			4376 => "00000000000000000100010011100001",
			4377 => "00000000000000000100010011100001",
			4378 => "0000001010000000000110011100000100",
			4379 => "11111111110001010100010011100001",
			4380 => "00000000000000000100010011100001",
			4381 => "0000000001000000001101101000011000",
			4382 => "0000001110000000000100000100010100",
			4383 => "0000000101000000001001110100001000",
			4384 => "0000001110000000000110000100000100",
			4385 => "00000000000000000100010011100001",
			4386 => "11111111000000110100010011100001",
			4387 => "0000000110000000001101011000000100",
			4388 => "00000000000000000100010011100001",
			4389 => "0000000000000000000101110100000100",
			4390 => "00000000110000110100010011100001",
			4391 => "00000000000000000100010011100001",
			4392 => "11111110100100110100010011100001",
			4393 => "0000000001000000001001011000010000",
			4394 => "0000000010000000001100001100001100",
			4395 => "0000000110000000001011001100000100",
			4396 => "00000000000000000100010011100001",
			4397 => "0000000001000000001011101000000100",
			4398 => "00000000000000000100010011100001",
			4399 => "00000000111010010100010011100001",
			4400 => "11111111110100110100010011100001",
			4401 => "0000000010000000000110001100000100",
			4402 => "11111111001101100100010011100001",
			4403 => "0000001010000000000001010000001000",
			4404 => "0000001001000000001001111100000100",
			4405 => "00000000010111010100010011100001",
			4406 => "00000000000000000100010011100001",
			4407 => "00000000000000000100010011100001",
			4408 => "0000000010000000001000001100101000",
			4409 => "0000000001000000000010001100000100",
			4410 => "11111110011000010100010110110101",
			4411 => "0000001010000000000101000100011100",
			4412 => "0000001111000000000000110100011000",
			4413 => "0000001010000000001010110000010000",
			4414 => "0000001111000000000000110100001000",
			4415 => "0000001010000000000110011000000100",
			4416 => "11111110011010100100010110110101",
			4417 => "11111111001101110100010110110101",
			4418 => "0000001010000000001001000100000100",
			4419 => "11111111100011000100010110110101",
			4420 => "00000101111000100100010110110101",
			4421 => "0000000011000000001110110000000100",
			4422 => "11111110101001100100010110110101",
			4423 => "00001100110010000100010110110101",
			4424 => "11111110011011010100010110110101",
			4425 => "0000001011000000001100101100000100",
			4426 => "11111110111000110100010110110101",
			4427 => "00000001110100100100010110110101",
			4428 => "0000001100000000000100001000110100",
			4429 => "0000000110000000000100111100101000",
			4430 => "0000001101000000000100010000010100",
			4431 => "0000001001000000001011101000001000",
			4432 => "0000000010000000001000001100000100",
			4433 => "00000000001001100100010110110101",
			4434 => "11111110010100110100010110110101",
			4435 => "0000001010000000001010110000000100",
			4436 => "11111110101001000100010110110101",
			4437 => "0000000110000000001101011000000100",
			4438 => "11111111101110000100010110110101",
			4439 => "00000010000000000100010110110101",
			4440 => "0000001001000000001000010000010000",
			4441 => "0000001110000000000111110000001000",
			4442 => "0000001001000000001101011000000100",
			4443 => "00000011001011110100010110110101",
			4444 => "11111111001001010100010110110101",
			4445 => "0000001000000000001011010100000100",
			4446 => "00000011111011110100010110110101",
			4447 => "00000111011110100100010110110101",
			4448 => "11111110100111110100010110110101",
			4449 => "0000000101000000001110101100001000",
			4450 => "0000001000000000001101010000000100",
			4451 => "11111110011001000100010110110101",
			4452 => "11111100100100110100010110110101",
			4453 => "00000001101101000100010110110101",
			4454 => "0000001110000000001101101100001100",
			4455 => "0000000010000000000101000000000100",
			4456 => "11111110011001100100010110110101",
			4457 => "0000001000000000000001110100000100",
			4458 => "00000101010000110100010110110101",
			4459 => "11111111000001110100010110110101",
			4460 => "11111110011000100100010110110101",
			4461 => "0000001101000000000100011000000100",
			4462 => "11111110011101000100011001101001",
			4463 => "0000001100000000000011011100011100",
			4464 => "0000001110000000000100001000001100",
			4465 => "0000000100000000001110111000000100",
			4466 => "00000000000000000100011001101001",
			4467 => "0000000110000000001111000000000100",
			4468 => "00000001101001100100011001101001",
			4469 => "00000000000000000100011001101001",
			4470 => "0000001100000000000011011100001000",
			4471 => "0000000100000000001101000000000100",
			4472 => "11111110101010100100011001101001",
			4473 => "00000000000101000100011001101001",
			4474 => "0000001001000000000001000100000100",
			4475 => "00000000000000000100011001101001",
			4476 => "00000001110001110100011001101001",
			4477 => "0000000110000000001011001100001100",
			4478 => "0000001100000000001100110000001000",
			4479 => "0000001110000000001010111100000100",
			4480 => "00000000000010110100011001101001",
			4481 => "00000000000000000100011001101001",
			4482 => "11111101111101000100011001101001",
			4483 => "0000000110000000001111000000011100",
			4484 => "0000000100000000001101110100001100",
			4485 => "0000001101000000001001010100000100",
			4486 => "11111111000010100100011001101001",
			4487 => "0000000001000000000000111100000100",
			4488 => "00000000111100010100011001101001",
			4489 => "11111111011010110100011001101001",
			4490 => "0000000001000000001101011100001000",
			4491 => "0000001001000000001111001100000100",
			4492 => "00000000000000000100011001101001",
			4493 => "00000001010110000100011001101001",
			4494 => "0000000010000000001111100100000100",
			4495 => "00000000010111010100011001101001",
			4496 => "11111111011000100100011001101001",
			4497 => "0000000010000000001000011100001000",
			4498 => "0000000011000000000010110100000100",
			4499 => "00000000000000000100011001101001",
			4500 => "11111110100000000100011001101001",
			4501 => "0000000011000000001111101000001000",
			4502 => "0000001010000000000101000100000100",
			4503 => "00000001000101100100011001101001",
			4504 => "00000000000000000100011001101001",
			4505 => "11111110111110010100011001101001",
			4506 => "0000001101000000000100011000000100",
			4507 => "11111110011011110100011100010101",
			4508 => "0000001100000000001100110000101100",
			4509 => "0000001100000000001001110000011000",
			4510 => "0000001110000000000100001000010000",
			4511 => "0000000100000000000111011100000100",
			4512 => "11111111111110100100011100010101",
			4513 => "0000000110000000001001100100001000",
			4514 => "0000001101000000001000011000000100",
			4515 => "00000001110011100100011100010101",
			4516 => "00000000000000000100011100010101",
			4517 => "00000000000000000100011100010101",
			4518 => "0000000100000000001101000000000100",
			4519 => "11111110100101100100011100010101",
			4520 => "00000000000000000100011100010101",
			4521 => "0000001111000000000110010000010000",
			4522 => "0000001000000000001001101000000100",
			4523 => "00000000000000000100011100010101",
			4524 => "0000000001000000001001111000000100",
			4525 => "00000000000000000100011100010101",
			4526 => "0000001010000000000001010000000100",
			4527 => "00000010100100010100011100010101",
			4528 => "00000001010000000100011100010101",
			4529 => "00000000000000000100011100010101",
			4530 => "0000000110000000001101011000001000",
			4531 => "0000001100000000001100110000000100",
			4532 => "00000000000000000100011100010101",
			4533 => "11111110010000110100011100010101",
			4534 => "0000000001000000000101011100011100",
			4535 => "0000001010000000001010110000001100",
			4536 => "0000001101000000000101110100000100",
			4537 => "11111111011010110100011100010101",
			4538 => "0000001010000000000110011000000100",
			4539 => "11111111111011010100011100010101",
			4540 => "00000001010001000100011100010101",
			4541 => "0000001111000000000111011000001000",
			4542 => "0000001010000000000101000100000100",
			4543 => "11111111100010000100011100010101",
			4544 => "00000001000000100100011100010101",
			4545 => "0000001001000000001001100100000100",
			4546 => "11111110100010000100011100010101",
			4547 => "00000000000000000100011100010101",
			4548 => "11111110100100000100011100010101",
			4549 => "0000001101000000000100011000000100",
			4550 => "11111110101000100100011110100001",
			4551 => "0000000010000000000010011100001100",
			4552 => "0000001011000000000110000100001000",
			4553 => "0000000100000000001111100100000100",
			4554 => "00000000000000000100011110100001",
			4555 => "00000001100111110100011110100001",
			4556 => "00000000000000000100011110100001",
			4557 => "0000000100000000000011010100000100",
			4558 => "11111110101111110100011110100001",
			4559 => "0000001010000000000110011100011100",
			4560 => "0000001100000000001110001100001100",
			4561 => "0000001100000000001000111000000100",
			4562 => "00000000000000000100011110100001",
			4563 => "0000001010000000000110011000000100",
			4564 => "00000000000000000100011110100001",
			4565 => "00000001001000100100011110100001",
			4566 => "0000001111000000000111011000001000",
			4567 => "0000001111000000001100010100000100",
			4568 => "00000000000000000100011110100001",
			4569 => "11111111100011000100011110100001",
			4570 => "0000000001000000000101011100000100",
			4571 => "00000000111001000100011110100001",
			4572 => "00000000000000000100011110100001",
			4573 => "0000000110000000000100111100010000",
			4574 => "0000000110000000001001100100001000",
			4575 => "0000001100000000001100110000000100",
			4576 => "00000000001110110100011110100001",
			4577 => "11111111010110010100011110100001",
			4578 => "0000000100000000000110110000000100",
			4579 => "00000000000000000100011110100001",
			4580 => "00000000101110100100011110100001",
			4581 => "0000000001000000001101011100000100",
			4582 => "11111110101011000100011110100001",
			4583 => "00000000000000000100011110100001",
			4584 => "0000001011000000000101101100000100",
			4585 => "11111110011101110100100000101101",
			4586 => "0000000100000000000010111000000100",
			4587 => "11111110100110100100100000101101",
			4588 => "0000001000000000000111000100011000",
			4589 => "0000000001000000000101011100010100",
			4590 => "0000001100000000000011011100000100",
			4591 => "00000001110111010100100000101101",
			4592 => "0000001100000000001110001100001000",
			4593 => "0000001101000000000101110100000100",
			4594 => "11111111010111010100100000101101",
			4595 => "00000000000000000100100000101101",
			4596 => "0000001101000000000101110100000100",
			4597 => "00000000000000000100100000101101",
			4598 => "00000001001111000100100000101101",
			4599 => "11111111010110100100100000101101",
			4600 => "0000000110000000001011001100010100",
			4601 => "0000001100000000001100110000001100",
			4602 => "0000000100000000000001100100000100",
			4603 => "11111111011110100100100000101101",
			4604 => "0000000001000000000010001100000100",
			4605 => "00000000000000000100100000101101",
			4606 => "00000001000000000100100000101101",
			4607 => "0000001110000000000100011000000100",
			4608 => "11111101111100100100100000101101",
			4609 => "00000000000000000100100000101101",
			4610 => "0000000110000000001111000000001100",
			4611 => "0000000100000000000010010000000100",
			4612 => "11111111001101000100100000101101",
			4613 => "0000000001000000001111001100000100",
			4614 => "00000001011011010100100000101101",
			4615 => "00000000000000000100100000101101",
			4616 => "0000001111000000001100010100000100",
			4617 => "00000000000000000100100000101101",
			4618 => "11111110110111100100100000101101",
			4619 => "0000000001000000001001111000000100",
			4620 => "11111110011111100100100011011011",
			4621 => "0000001010000000000110011100100100",
			4622 => "0000000000000000001111000100000100",
			4623 => "11111110110000000100100011011011",
			4624 => "0000001100000000001000111000000100",
			4625 => "11111111001000010100100011011011",
			4626 => "0000001010000000000001010000001100",
			4627 => "0000000001000000000000111100001000",
			4628 => "0000001010000000001001000100000100",
			4629 => "00000000000000000100100011011011",
			4630 => "00000001101110100100100011011011",
			4631 => "00000000000000000100100011011011",
			4632 => "0000000100000000001100111100001000",
			4633 => "0000001100000000000000001100000100",
			4634 => "11111111001010000100100011011011",
			4635 => "00000000000000000100100011011011",
			4636 => "0000001110000000000100010000000100",
			4637 => "00000000000000000100100011011011",
			4638 => "00000001100100100100100011011011",
			4639 => "0000000000000000001100101100101000",
			4640 => "0000001100000000001110001100011100",
			4641 => "0000001100000000001100110000010000",
			4642 => "0000000101000000001001110100001000",
			4643 => "0000000110000000001011001100000100",
			4644 => "00000000000000000100100011011011",
			4645 => "11111111101110110100100011011011",
			4646 => "0000000110000000001000010000000100",
			4647 => "00000000010100000100100011011011",
			4648 => "00000000000000000100100011011011",
			4649 => "0000000010000000001111100100000100",
			4650 => "00000000000000000100100011011011",
			4651 => "0000000010000000000011000000000100",
			4652 => "11111101111101100100100011011011",
			4653 => "00000000000000000100100011011011",
			4654 => "0000001100000000000100001000001000",
			4655 => "0000001001000000000111101000000100",
			4656 => "00000000000000000100100011011011",
			4657 => "00000000110001100100100011011011",
			4658 => "11111111101010010100100011011011",
			4659 => "0000000010000000001100001100000100",
			4660 => "00000001000000100100100011011011",
			4661 => "00000000000000000100100011011011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1522, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(3074, initial_addr_3'length));
	end generate gen_rom_13;

	gen_rom_14: if SELECT_ROM = 14 generate
		bank <= (
			0 => "0000000111000000001101111001011000",
			1 => "0000000100000000001011100101010100",
			2 => "0000000110000000000001000100010100",
			3 => "0000000011000000000000111000001000",
			4 => "0000001111000000001000000000000100",
			5 => "00000010010111110000000011010101",
			6 => "11111111010101010000000011010101",
			7 => "0000000011000000000111111000001000",
			8 => "0000001110000000001010101100000100",
			9 => "11111110101011110000000011010101",
			10 => "00000000011101000000000011010101",
			11 => "11111110011000100000000011010101",
			12 => "0000000111000000001100001000100000",
			13 => "0000000011000000001101100000010000",
			14 => "0000000111000000000111111000001000",
			15 => "0000000010000000000010000000000100",
			16 => "00000001111110110000000011010101",
			17 => "11111110011000010000000011010101",
			18 => "0000001010000000000111110100000100",
			19 => "00000010100100100000000011010101",
			20 => "00000000011001000000000011010101",
			21 => "0000000010000000001001010000001000",
			22 => "0000000100000000000010111000000100",
			23 => "00000001100001000000000011010101",
			24 => "00000011000111010000000011010101",
			25 => "0000001010000000000110011000000100",
			26 => "00000000001101100000000011010101",
			27 => "00000001001010110000000011010101",
			28 => "0000001110000000001101111000010000",
			29 => "0000000010000000001100010100001000",
			30 => "0000000110000000000001111000000100",
			31 => "11111110111101110000000011010101",
			32 => "00000000011101110000000011010101",
			33 => "0000000111000000001000111000000100",
			34 => "11111111000110100000000011010101",
			35 => "00000001001111110000000011010101",
			36 => "0000000111000000001000111000001000",
			37 => "0000001110000000000100000100000100",
			38 => "00000001001101110000000011010101",
			39 => "11111110100001010000000011010101",
			40 => "0000000110000000001111000000000100",
			41 => "00000000100001000000000011010101",
			42 => "11111110111111000000000011010101",
			43 => "11111110010111100000000011010101",
			44 => "0000001010000000000111110100010000",
			45 => "0000001111000000001000101000001100",
			46 => "0000000111000000001100101000001000",
			47 => "0000001000000000000000001000000100",
			48 => "11111110101111010000000011010101",
			49 => "00000001010110100000000011010101",
			50 => "11111110010111110000000011010101",
			51 => "00000011100101110000000011010101",
			52 => "11111110010111100000000011010101",
			53 => "0000000000000000001100001010001000",
			54 => "0000000101000000001000111100011100",
			55 => "0000000000000000000111111000001100",
			56 => "0000001001000000001100110100001000",
			57 => "0000000101000000001100001000000100",
			58 => "00000000000000000000001001011001",
			59 => "11111111101110000000001001011001",
			60 => "00000010000010110000001001011001",
			61 => "0000000100000000001111100000000100",
			62 => "11111110101101110000001001011001",
			63 => "0000001011000000001010000000000100",
			64 => "00000000000000000000001001011001",
			65 => "0000001010000000000001010000000100",
			66 => "00000000000000000000001001011001",
			67 => "00000001110000100000001001011001",
			68 => "0000000001000000001110100000110000",
			69 => "0000001001000000001001111000100000",
			70 => "0000000010000000001001010000010000",
			71 => "0000000110000000001101111100001000",
			72 => "0000001111000000001011011100000100",
			73 => "11111111101101110000001001011001",
			74 => "00000011000011110000001001011001",
			75 => "0000000001000000000110000000000100",
			76 => "00000000001101000000001001011001",
			77 => "00000010001011100000001001011001",
			78 => "0000000010000000000101110000001000",
			79 => "0000000000000000000000111000000100",
			80 => "00000001111100110000001001011001",
			81 => "11111110011010110000001001011001",
			82 => "0000000001000000000110000000000100",
			83 => "00000000100001000000001001011001",
			84 => "11111111010100100000001001011001",
			85 => "0000000101000000000011011100001000",
			86 => "0000001110000000001110111100000100",
			87 => "11111110010100100000001001011001",
			88 => "00000000111000100000001001011001",
			89 => "0000001010000000001010110000000100",
			90 => "11111101110011010000001001011001",
			91 => "11111111101100100000001001011001",
			92 => "0000001101000000001100101100011100",
			93 => "0000000011000000000101101100001100",
			94 => "0000001011000000001100001000001000",
			95 => "0000001011000000000000101000000100",
			96 => "11111111111110110000001001011001",
			97 => "00000000110100110000001001011001",
			98 => "11111101011101100000001001011001",
			99 => "0000000010000000001100010100001000",
			100 => "0000000000000000000000111000000100",
			101 => "00000000011111010000001001011001",
			102 => "00000001101001100000001001011001",
			103 => "0000001001000000000110101000000100",
			104 => "00000000110100000000001001011001",
			105 => "11111110001000100000001001011001",
			106 => "0000000001000000001100110100010000",
			107 => "0000001011000000000100000000001000",
			108 => "0000001101000000001101111000000100",
			109 => "11111111101011100000001001011001",
			110 => "11111110001000000000001001011001",
			111 => "0000000001000000001110100000000100",
			112 => "00000001110111110000001001011001",
			113 => "11111111110110110000001001011001",
			114 => "0000001001000000000111100100001000",
			115 => "0000000011000000001101111000000100",
			116 => "00000000001111100000001001011001",
			117 => "00000001011101110000001001011001",
			118 => "0000000001000000001100110100000100",
			119 => "11111111100001000000001001011001",
			120 => "00000000000000100000001001011001",
			121 => "0000000010000000000010000000100100",
			122 => "0000001110000000000000101000100000",
			123 => "0000000011000000000100000000010100",
			124 => "0000001111000000000110110100010000",
			125 => "0000001010000000000110011100001000",
			126 => "0000001110000000000011111100000100",
			127 => "11111110011101010000001001011001",
			128 => "00000000011000110000001001011001",
			129 => "0000000000000000001000111100000100",
			130 => "00000000100110010000001001011001",
			131 => "11111111011011000000001001011001",
			132 => "00000010110010000000001001011001",
			133 => "0000001010000000000001010100000100",
			134 => "11111110100001010000001001011001",
			135 => "0000001111000000001011011100000100",
			136 => "00000000111100010000001001011001",
			137 => "11111111011000100000001001011001",
			138 => "00000001001100010000001001011001",
			139 => "0000000001000000000010001100010000",
			140 => "0000001000000000001000110000000100",
			141 => "11111110010100010000001001011001",
			142 => "0000000001000000001110100000001000",
			143 => "0000001111000000000101110100000100",
			144 => "11111111111000100000001001011001",
			145 => "00000001100001000000001001011001",
			146 => "11111110101111000000001001011001",
			147 => "0000001011000000001100110000000100",
			148 => "00000001000111010000001001011001",
			149 => "11111110111010110000001001011001",
			150 => "0000001001000000001001111001010000",
			151 => "0000001100000000000100010100101100",
			152 => "0000001100000000000100010100101000",
			153 => "0000000010000000000010000000100000",
			154 => "0000000100000000000001101100010000",
			155 => "0000001110000000001111000100001000",
			156 => "0000001011000000000100010100000100",
			157 => "11111111111001110000001110111101",
			158 => "11111110011010000000001110111101",
			159 => "0000001100000000000000110000000100",
			160 => "11111111100100010000001110111101",
			161 => "00000000011101100000001110111101",
			162 => "0000001010000000000001010100001000",
			163 => "0000001101000000001000111000000100",
			164 => "00000011010001110000001110111101",
			165 => "00000000111110110000001110111101",
			166 => "0000001011000000000111111000000100",
			167 => "11111111010101100000001110111101",
			168 => "00000001001011000000001110111101",
			169 => "0000000100000000000100001100000100",
			170 => "00000000011000000000001110111101",
			171 => "11111101111100010000001110111101",
			172 => "11111110010101110000001110111101",
			173 => "0000000001000000000110000000001100",
			174 => "0000001110000000000000111000001000",
			175 => "0000000001000000000000011000000100",
			176 => "00000000000000000000001110111101",
			177 => "11111110010111110000001110111101",
			178 => "00000000010011010000001110111101",
			179 => "0000001100000000000000101000010100",
			180 => "0000001110000000001110111100010000",
			181 => "0000001101000000001100110000001000",
			182 => "0000001001000000000010001100000100",
			183 => "00000001110111000000001110111101",
			184 => "00000000010111000000001110111101",
			185 => "0000001011000000001011000100000100",
			186 => "11111111000011010000001110111101",
			187 => "00000000110000110000001110111101",
			188 => "00000010101101110000001110111101",
			189 => "11111110011010110000001110111101",
			190 => "0000000001000000001110100000110000",
			191 => "0000001100000000000000110000000100",
			192 => "00000001100100100000001110111101",
			193 => "0000000010000000001001011100010100",
			194 => "0000000100000000001011100000010000",
			195 => "0000001110000000000100010100001000",
			196 => "0000000111000000000111111000000100",
			197 => "00000001011000010000001110111101",
			198 => "11111111100001010000001110111101",
			199 => "0000000001000000001110100000000100",
			200 => "11111111110101100000001110111101",
			201 => "00000001010001110000001110111101",
			202 => "00000001101111110000001110111101",
			203 => "0000001001000000001001111000001100",
			204 => "0000001001000000001001111000001000",
			205 => "0000001111000000001011110100000100",
			206 => "11111110000001100000001110111101",
			207 => "11111111111010000000001110111101",
			208 => "00000000100100010000001110111101",
			209 => "0000000110000000000100110100000100",
			210 => "11111110000010000000001110111101",
			211 => "0000000000000000001011000100000100",
			212 => "00000000000011110000001110111101",
			213 => "11111110001100100000001110111101",
			214 => "0000000111000000000111111000000100",
			215 => "00000001011100110000001110111101",
			216 => "0000001100000000001010000000010100",
			217 => "0000001101000000000110000100001100",
			218 => "0000000001000000001110100000001000",
			219 => "0000001110000000000100010100000100",
			220 => "11111110011100010000001110111101",
			221 => "00000000001011110000001110111101",
			222 => "00000001011011100000001110111101",
			223 => "0000000100000000001110111000000100",
			224 => "11111110001100000000001110111101",
			225 => "11111111110000000000001110111101",
			226 => "0000001100000000001110111100001100",
			227 => "0000000010000000001111010000000100",
			228 => "11111111011011000000001110111101",
			229 => "0000000111000000000100010100000100",
			230 => "00000010101011100000001110111101",
			231 => "00000000100101100000001110111101",
			232 => "0000001101000000001100110000001000",
			233 => "0000000100000000001110111000000100",
			234 => "11111110000100100000001110111101",
			235 => "00000000010001010000001110111101",
			236 => "0000001100000000001000111000000100",
			237 => "00000000000100010000001110111101",
			238 => "11111111101110110000001110111101",
			239 => "0000001100000000000100000010010100",
			240 => "0000000111000000001001110001100100",
			241 => "0000000111000000001000111000111100",
			242 => "0000001100000000000100000000100000",
			243 => "0000000010000000000100101000010000",
			244 => "0000000010000000000100101000001000",
			245 => "0000000001000000000010001100000100",
			246 => "00000000000010100000010101110001",
			247 => "00000000110110000000010101110001",
			248 => "0000001010000000001010110000000100",
			249 => "00000001011010110000010101110001",
			250 => "11111111100010110000010101110001",
			251 => "0000001010000000001010110000001000",
			252 => "0000001110000000001101100000000100",
			253 => "11111111100101110000010101110001",
			254 => "11111111111110000000010101110001",
			255 => "0000001100000000000100010100000100",
			256 => "11111111100011100000010101110001",
			257 => "00000000011011100000010101110001",
			258 => "0000001010000000001100011100010000",
			259 => "0000001011000000000100000000001000",
			260 => "0000000010000000001001010000000100",
			261 => "11111111111010110000010101110001",
			262 => "00000001100010010000010101110001",
			263 => "0000001111000000000110100000000100",
			264 => "11111110111110000000010101110001",
			265 => "11111111111110100000010101110001",
			266 => "0000001010000000001100011100000100",
			267 => "00000001111101000000010101110001",
			268 => "0000000110000000001101011000000100",
			269 => "11111111000011000000010101110001",
			270 => "00000001001011010000010101110001",
			271 => "0000000000000000000111111000100000",
			272 => "0000001000000000000110001000010000",
			273 => "0000001111000000001100100100001000",
			274 => "0000001100000000000000101000000100",
			275 => "11111111100100000000010101110001",
			276 => "00000001010000010000010101110001",
			277 => "0000001010000000000001010000000100",
			278 => "11111110001101100000010101110001",
			279 => "00000001000101010000010101110001",
			280 => "0000001010000000001010110000001000",
			281 => "0000001101000000001010111000000100",
			282 => "00000010010010010000010101110001",
			283 => "00000001010011100000010101110001",
			284 => "0000000011000000000001101000000100",
			285 => "11111111100011100000010101110001",
			286 => "00000001110000100000010101110001",
			287 => "0000001101000000000111001000000100",
			288 => "11111101111010110000010101110001",
			289 => "00000000100011000000010101110001",
			290 => "0000000010000000000010000100011100",
			291 => "0000000001000000000110101000010000",
			292 => "0000000010000000000101110000000100",
			293 => "00000000111111010000010101110001",
			294 => "0000000111000000001101100000000100",
			295 => "11111101111001100000010101110001",
			296 => "0000001110000000001110110000000100",
			297 => "11111111111011110000010101110001",
			298 => "11111101111100010000010101110001",
			299 => "0000001101000000001001001000000100",
			300 => "00000001100000010000010101110001",
			301 => "0000000111000000001101100000000100",
			302 => "11111110001011000000010101110001",
			303 => "00000000011000100000010101110001",
			304 => "0000000000000000000000111000001000",
			305 => "0000001011000000001110001100000100",
			306 => "11111101111111100000010101110001",
			307 => "00000000000101000000010101110001",
			308 => "0000000110000000001011001100000100",
			309 => "00000001111011010000010101110001",
			310 => "0000000111000000001101100000000100",
			311 => "11111110011011000000010101110001",
			312 => "00000000110101000000010101110001",
			313 => "0000001100000000000100000000011000",
			314 => "0000000010000000000011001000001000",
			315 => "0000000010000000001111010000000100",
			316 => "00000000000000000000010101110001",
			317 => "00000010001010010000010101110001",
			318 => "0000000010000000001100010100000100",
			319 => "11111111010010010000010101110001",
			320 => "0000001101000000001010111100000100",
			321 => "11111111110001000000010101110001",
			322 => "0000000001000000001001111000000100",
			323 => "00000010000000010000010101110001",
			324 => "00000000000000000000010101110001",
			325 => "0000000000000000000100010100101000",
			326 => "0000001000000000000010101000100000",
			327 => "0000001100000000001000111100010000",
			328 => "0000001100000000001000111100001000",
			329 => "0000001110000000001010111000000100",
			330 => "11111111101101110000010101110001",
			331 => "00000001011000010000010101110001",
			332 => "0000000110000000001010011000000100",
			333 => "11111111110110100000010101110001",
			334 => "11111110001000010000010101110001",
			335 => "0000000001000000000010001100001000",
			336 => "0000000110000000001010011000000100",
			337 => "00000000000000000000010101110001",
			338 => "11111101111100110000010101110001",
			339 => "0000000110000000001010011000000100",
			340 => "00000000111010100000010101110001",
			341 => "00000000000001010000010101110001",
			342 => "0000000010000000000111010100000100",
			343 => "00000011001011100000010101110001",
			344 => "00000000000000000000010101110001",
			345 => "0000001011000000001001110000000100",
			346 => "00000000000011010000010101110001",
			347 => "11111110011000000000010101110001",
			348 => "0000000111000000000101101101111000",
			349 => "0000000001000000000000011000001000",
			350 => "0000000110000000000100110100000100",
			351 => "11111110010101100000011011010101",
			352 => "00000000111011010000011011010101",
			353 => "0000000100000000001110111000111100",
			354 => "0000000110000000001101111100100000",
			355 => "0000000010000000000101110000010000",
			356 => "0000000000000000000000110000001000",
			357 => "0000000110000000001101111100000100",
			358 => "00000000101101100000011011010101",
			359 => "00000001100111110000011011010101",
			360 => "0000000100000000000101010100000100",
			361 => "11111110100001010000011011010101",
			362 => "00000000011111110000011011010101",
			363 => "0000000000000000001111000100001000",
			364 => "0000000100000000001011110000000100",
			365 => "00000000000000000000011011010101",
			366 => "11111110000001110000011011010101",
			367 => "0000000011000000001101111000000100",
			368 => "11111111101101010000011011010101",
			369 => "00000001001110000000011011010101",
			370 => "0000001100000000000100000000001100",
			371 => "0000000001000000000110101000001000",
			372 => "0000000100000000000011001100000100",
			373 => "00000010000000010000011011010101",
			374 => "00000001011001110000011011010101",
			375 => "11111110000110100000011011010101",
			376 => "0000001100000000000100000000001000",
			377 => "0000000100000000000011001100000100",
			378 => "11111101001111100000011011010101",
			379 => "11111110011101010000011011010101",
			380 => "0000000110000000001001100100000100",
			381 => "00000000111010010000011011010101",
			382 => "11111110100001000000011011010101",
			383 => "0000001100000000000100010100010100",
			384 => "0000001010000000000110011000000100",
			385 => "11111110010110110000011011010101",
			386 => "0000001001000000001001111000001000",
			387 => "0000000011000000001100001000000100",
			388 => "00000000111000100000011011010101",
			389 => "00000011000001010000011011010101",
			390 => "0000000011000000001001110000000100",
			391 => "11111111110101000000011011010101",
			392 => "00000001001001000000011011010101",
			393 => "0000000110000000001100011000010000",
			394 => "0000000010000000001001011100001000",
			395 => "0000000111000000000100010100000100",
			396 => "11111110100100110000011011010101",
			397 => "00000000011010010000011011010101",
			398 => "0000001001000000000111100100000100",
			399 => "11111111010111010000011011010101",
			400 => "11111101111011010000011011010101",
			401 => "0000000100000000000010100100001000",
			402 => "0000001001000000000110101000000100",
			403 => "00000001101111100000011011010101",
			404 => "00000000011110010000011011010101",
			405 => "0000001100000000000100010100000100",
			406 => "00000000101000110000011011010101",
			407 => "11111111001010100000011011010101",
			408 => "0000001100000000000110000100100100",
			409 => "0000001101000000000111010000010000",
			410 => "0000001110000000001001001000000100",
			411 => "11111110010100100000011011010101",
			412 => "0000001110000000000100000100001000",
			413 => "0000000000000000001101010000000100",
			414 => "11111110101000010000011011010101",
			415 => "00000001110110100000011011010101",
			416 => "11111110001111110000011011010101",
			417 => "0000000100000000001001001100010000",
			418 => "0000000000000000001001101000000100",
			419 => "11111110011100110000011011010101",
			420 => "0000000110000000001111000000000100",
			421 => "00000011100100000000011011010101",
			422 => "0000001010000000001100011100000100",
			423 => "11111110011101000000011011010101",
			424 => "00000000010100100000011011010101",
			425 => "11111110011000100000011011010101",
			426 => "0000001100000000001010111100010100",
			427 => "0000000111000000000110100100010000",
			428 => "0000000111000000001101111000001100",
			429 => "0000000111000000001110001100000100",
			430 => "11111110100000100000011011010101",
			431 => "0000001100000000000110000100000100",
			432 => "00000000110011000000011011010101",
			433 => "11111111000001000000011011010101",
			434 => "11111110010111100000011011010101",
			435 => "00000100100111110000011011010101",
			436 => "11111110010101010000011011010101",
			437 => "0000001110000000001000000010010000",
			438 => "0000001001000000001111001101011100",
			439 => "0000000001000000001001111000110000",
			440 => "0000001001000000001011101000100000",
			441 => "0000000110000000001100011000010000",
			442 => "0000000010000000001100010100001000",
			443 => "0000001100000000000000101000000100",
			444 => "11111111111110010000100010101001",
			445 => "00000000011010100000100010101001",
			446 => "0000001001000000001101101000000100",
			447 => "11111111101100000000100010101001",
			448 => "11111110011000110000100010101001",
			449 => "0000001100000000000100000000001000",
			450 => "0000000011000000000101101100000100",
			451 => "11111111101011010000100010101001",
			452 => "00000000011101000000100010101001",
			453 => "0000000011000000000100011000000100",
			454 => "11111111000111010000100010101001",
			455 => "00000000111110000000100010101001",
			456 => "0000000100000000000011010100001100",
			457 => "0000000101000000000111001000001000",
			458 => "0000000000000000001110111100000100",
			459 => "11111111110011110000100010101001",
			460 => "11111101111110000000100010101001",
			461 => "11111101100011000000100010101001",
			462 => "00000001001101000000100010101001",
			463 => "0000000100000000000011110000010100",
			464 => "0000000110000000000001111000001000",
			465 => "0000001001000000001011101000000100",
			466 => "00000000000000000000100010101001",
			467 => "00000100100000100000100010101001",
			468 => "0000000011000000001110110000001000",
			469 => "0000000111000000001000111000000100",
			470 => "00000001101011010000100010101001",
			471 => "00000000000000000000100010101001",
			472 => "00000001110100110000100010101001",
			473 => "0000000011000000001000000000001100",
			474 => "0000001001000000001011101000000100",
			475 => "00000001101111100000100010101001",
			476 => "0000000000000000000000110000000100",
			477 => "11111111101011100000100010101001",
			478 => "11111110001000000000100010101001",
			479 => "0000000100000000000100001100001000",
			480 => "0000000001000000001001111000000100",
			481 => "00000010101100100000100010101001",
			482 => "00000000110110100000100010101001",
			483 => "11111111110000100000100010101001",
			484 => "0000000000000000000000110000011100",
			485 => "0000000001000000001001111000000100",
			486 => "11111110010110100000100010101001",
			487 => "0000000100000000001000001000001100",
			488 => "0000000001000000000110101000001000",
			489 => "0000000011000000001001001000000100",
			490 => "11111111000100110000100010101001",
			491 => "00000000100000110000100010101001",
			492 => "11111101110011110000100010101001",
			493 => "0000000100000000000010111000000100",
			494 => "00000001111111110000100010101001",
			495 => "0000000010000000000110010000000100",
			496 => "11111110110010010000100010101001",
			497 => "00000001000111100000100010101001",
			498 => "0000001001000000001001011000010000",
			499 => "0000000110000000001001100100000100",
			500 => "11111110010011100000100010101001",
			501 => "0000000101000000000100011000000100",
			502 => "11111110111101110000100010101001",
			503 => "0000000001000000001001111000000100",
			504 => "00000001011001100000100010101001",
			505 => "00000000000000000000100010101001",
			506 => "0000001011000000000000001100000100",
			507 => "00000001010111000000100010101001",
			508 => "00000000000000000000100010101001",
			509 => "0000000110000000001001100101000100",
			510 => "0000001100000000001000111100100100",
			511 => "0000001100000000000000101000001000",
			512 => "0000000100000000000011110000000100",
			513 => "00000001101100110000100010101001",
			514 => "11111101100100110000100010101001",
			515 => "0000001000000000000110001000010000",
			516 => "0000001000000000001001101000001000",
			517 => "0000000010000000000111111100000100",
			518 => "00000000000000000000100010101001",
			519 => "00000001100001000000100010101001",
			520 => "0000001000000000001011010100000100",
			521 => "11111110111110010000100010101001",
			522 => "00000000100010100000100010101001",
			523 => "0000001100000000000100000000001000",
			524 => "0000001100000000001100001000000100",
			525 => "00000001000001010000100010101001",
			526 => "00000010100010100000100010101001",
			527 => "00000000110001000000100010101001",
			528 => "0000001100000000001000111100000100",
			529 => "11111101110000100000100010101001",
			530 => "0000000011000000001111011100001100",
			531 => "0000000111000000000101101100000100",
			532 => "11111110100111010000100010101001",
			533 => "0000000101000000000001101000000100",
			534 => "00000001010101100000100010101001",
			535 => "00000000000000000000100010101001",
			536 => "0000000011000000000100000100001000",
			537 => "0000001100000000000011011100000100",
			538 => "00000001111000000000100010101001",
			539 => "11111111000011110000100010101001",
			540 => "0000001101000000000001101000000100",
			541 => "11111111100101110000100010101001",
			542 => "00000000101101000000100010101001",
			543 => "0000001101000000001000000000001000",
			544 => "0000001110000000001000011000000100",
			545 => "11111111011100110000100010101001",
			546 => "00000001001100110000100010101001",
			547 => "0000000110000000000100111100000100",
			548 => "11111110010111100000100010101001",
			549 => "0000000010000000001111010100001000",
			550 => "0000000101000000000110100100000100",
			551 => "00000000000000000000100010101001",
			552 => "00000001100010010000100010101001",
			553 => "11111110101101000000100010101001",
			554 => "0000001100000000000110000110001000",
			555 => "0000000001000000000000011000001100",
			556 => "0000000110000000000100110100000100",
			557 => "11111110010110100000100111100101",
			558 => "0000000111000000000111111000000100",
			559 => "00000001101001000000100111100101",
			560 => "11111110111001100000100111100101",
			561 => "0000001001000000001001111001000000",
			562 => "0000000011000000000100000000100000",
			563 => "0000001001000000001001111000010000",
			564 => "0000000011000000000100010100001000",
			565 => "0000001100000000000000110000000100",
			566 => "00000001101010100000100111100101",
			567 => "11111111111010000000100111100101",
			568 => "0000001111000000000110100100000100",
			569 => "00000100101000100000100111100101",
			570 => "00000000101001000000100111100101",
			571 => "0000000001000000001110100000001000",
			572 => "0000001100000000000111111000000100",
			573 => "11111111100010010000100111100101",
			574 => "11111110001000000000100111100101",
			575 => "0000001111000000001010001100000100",
			576 => "00000001110110100000100111100101",
			577 => "11111110111111100000100111100101",
			578 => "0000001111000000000101100100010000",
			579 => "0000001110000000000000110000001000",
			580 => "0000001010000000000001010000000100",
			581 => "11111111010010110000100111100101",
			582 => "00000010111110110000100111100101",
			583 => "0000000000000000001111000100000100",
			584 => "11111111001111010000100111100101",
			585 => "00000011100011010000100111100101",
			586 => "0000001000000000001001101000001000",
			587 => "0000001110000000000100010100000100",
			588 => "11111110001000110000100111100101",
			589 => "00000000011111100000100111100101",
			590 => "0000000011000000001001110000000100",
			591 => "00000000001010000000100111100101",
			592 => "00000001100111000000100111100101",
			593 => "0000001110000000001000111100011100",
			594 => "0000000011000000001110001100010000",
			595 => "0000000011000000001100101100001000",
			596 => "0000000011000000001100101100000100",
			597 => "00000000001000010000100111100101",
			598 => "11111110001100010000100111100101",
			599 => "0000000010000000001001011100000100",
			600 => "00000001110011000000100111100101",
			601 => "11111111101100100000100111100101",
			602 => "0000001000000000001010101100001000",
			603 => "0000001111000000000101100100000100",
			604 => "00000000100100100000100111100101",
			605 => "11111110111000000000100111100101",
			606 => "00000100111010010000100111100101",
			607 => "0000001001000000001101101000010000",
			608 => "0000000010000000000010000000001000",
			609 => "0000000111000000001100001000000100",
			610 => "00000000101011010000100111100101",
			611 => "00000001010110000000100111100101",
			612 => "0000000110000000001100011000000100",
			613 => "11111111000110000000100111100101",
			614 => "00000000100010110000100111100101",
			615 => "0000001110000000001101111000001000",
			616 => "0000001101000000001101111000000100",
			617 => "00000010000111000000100111100101",
			618 => "11111111101111100000100111100101",
			619 => "0000001001000000001111001100000100",
			620 => "00000000101111100000100111100101",
			621 => "11111111111110010000100111100101",
			622 => "0000001100000000001010111100010100",
			623 => "0000001101000000001001010000010000",
			624 => "0000000111000000001101111000001100",
			625 => "0000000111000000001110001100000100",
			626 => "11111110101101000000100111100101",
			627 => "0000001100000000000110000100000100",
			628 => "00000000011000010000100111100101",
			629 => "00000000000000000000100111100101",
			630 => "11111110011010110000100111100101",
			631 => "00000011000001110000100111100101",
			632 => "11111110011001010000100111100101",
			633 => "0000000111000000000101101101101100",
			634 => "0000000001000000001100100000000100",
			635 => "11111110010110100000101101000001",
			636 => "0000000100000000001110111000111000",
			637 => "0000000111000000001001110000100000",
			638 => "0000000110000000001101111100010000",
			639 => "0000000010000000000111111100001000",
			640 => "0000001110000000001000111100000100",
			641 => "00000000100110100000101101000001",
			642 => "00000001010111110000101101000001",
			643 => "0000000000000000000010111100000100",
			644 => "11111110101100110000101101000001",
			645 => "00000000010000000000101101000001",
			646 => "0000000111000000001100001000001000",
			647 => "0000001111000000001011110100000100",
			648 => "00000010011000100000101101000001",
			649 => "00000001100010110000101101000001",
			650 => "0000001110000000000110000100000100",
			651 => "00000000101001110000101101000001",
			652 => "00000001100000100000101101000001",
			653 => "0000001000000000000111000100001100",
			654 => "0000000110000000001001100100001000",
			655 => "0000001111000000001010010100000100",
			656 => "11111110101110010000101101000001",
			657 => "00000001000100110000101101000001",
			658 => "11111110010110100000101101000001",
			659 => "0000000100000000001001001100001000",
			660 => "0000000010000000000110111100000100",
			661 => "11111101111100100000101101000001",
			662 => "00000000000000000000101101000001",
			663 => "11111111111101110000101101000001",
			664 => "0000001001000000000110101000010100",
			665 => "0000000110000000000111101000000100",
			666 => "11111110010111110000101101000001",
			667 => "0000001110000000001011000100001000",
			668 => "0000000111000000000111111000000100",
			669 => "00000001100010100000101101000001",
			670 => "00000000011011100000101101000001",
			671 => "0000000010000000001100010100000100",
			672 => "00000010101110100000101101000001",
			673 => "00000001000010000000101101000001",
			674 => "0000000011000000000101101100001100",
			675 => "0000001101000000000110000100000100",
			676 => "00000001111101100000101101000001",
			677 => "0000000010000000001111010000000100",
			678 => "00000000000111010000101101000001",
			679 => "11111110101010110000101101000001",
			680 => "0000000110000000001100011000001000",
			681 => "0000001110000000001001110000000100",
			682 => "00000000000000110000101101000001",
			683 => "11111110010110110000101101000001",
			684 => "0000000100000000001111100000000100",
			685 => "00000000110101000000101101000001",
			686 => "11111111111001100000101101000001",
			687 => "0000000111000000001100101000100100",
			688 => "0000001110000000001001001000000100",
			689 => "11111110010101110000101101000001",
			690 => "0000000010000000000111010100011100",
			691 => "0000001101000000000111010000001100",
			692 => "0000001110000000000100000100001000",
			693 => "0000000000000000001101010000000100",
			694 => "11111110100111000000101101000001",
			695 => "00000001001110000000101101000001",
			696 => "11111110010010000000101101000001",
			697 => "0000000110000000000100110100001000",
			698 => "0000001011000000001010111000000100",
			699 => "11111110011001100000101101000001",
			700 => "00000000000000000000101101000001",
			701 => "0000001011000000001101010100000100",
			702 => "00000011111111010000101101000001",
			703 => "00000000110111010000101101000001",
			704 => "11111110011001110000101101000001",
			705 => "0000001000000000000110011100011100",
			706 => "0000000100000000001011110000010000",
			707 => "0000000111000000000001111100001100",
			708 => "0000000111000000000001111100001000",
			709 => "0000000111000000001100101000000100",
			710 => "00000000000000000000101101000001",
			711 => "11111111110010100000101101000001",
			712 => "00000000110111000000101101000001",
			713 => "11111110010110100000101101000001",
			714 => "0000000000000000000111000100000100",
			715 => "00000100110111000000101101000001",
			716 => "0000000100000000001000110100000100",
			717 => "11111110100000110000101101000001",
			718 => "00000001110100010000101101000001",
			719 => "11111110010110000000101101000001",
			720 => "0000001001000000001001111001101000",
			721 => "0000001100000000000100010100111000",
			722 => "0000001100000000000100010100110100",
			723 => "0000000100000000000001101100011100",
			724 => "0000001110000000001111000100001100",
			725 => "0000001011000000000100010100001000",
			726 => "0000000010000000000010110100000100",
			727 => "00000000110010010000110011011101",
			728 => "11111111100000010000110011011101",
			729 => "11111110010111010000110011011101",
			730 => "0000001111000000000000011100001000",
			731 => "0000001000000000000111000100000100",
			732 => "00000000010101110000110011011101",
			733 => "00000001011110000000110011011101",
			734 => "0000001100000000000111111000000100",
			735 => "11111111111001000000110011011101",
			736 => "00000010010000000000110011011101",
			737 => "0000001010000000000001010100001100",
			738 => "0000000010000000001101000100000100",
			739 => "00000101110110110000110011011101",
			740 => "0000000100000000001100111100000100",
			741 => "00000001111000000000110011011101",
			742 => "11111111111111110000110011011101",
			743 => "0000001010000000000001110000000100",
			744 => "11111110011000000000110011011101",
			745 => "0000000100000000000011111000000100",
			746 => "00000000111101000000110011011101",
			747 => "11111111011100010000110011011101",
			748 => "11111110010010000000110011011101",
			749 => "0000000001000000000110000000001000",
			750 => "0000001110000000000000111000000100",
			751 => "11111110011010110000110011011101",
			752 => "00000000011100100000110011011101",
			753 => "0000000010000000000001000000010100",
			754 => "0000000010000000001110101000001100",
			755 => "0000000111000000000100010100001000",
			756 => "0000000110000000000001111000000100",
			757 => "00000001000011000000110011011101",
			758 => "11111110100001110000110011011101",
			759 => "00000010011101000000110011011101",
			760 => "0000000100000000001110111000000100",
			761 => "11111110001100100000110011011101",
			762 => "00000000011001100000110011011101",
			763 => "0000001100000000000100010100001100",
			764 => "0000001101000000001101100000000100",
			765 => "00000011000111010000110011011101",
			766 => "0000001110000000000000111000000100",
			767 => "11111111101001100000110011011101",
			768 => "00000010101101100000110011011101",
			769 => "0000001010000000001100011100000100",
			770 => "00000001100001000000110011011101",
			771 => "11111111001011100000110011011101",
			772 => "0000000001000000001110100000101000",
			773 => "0000001100000000000000110000000100",
			774 => "00000001101100110000110011011101",
			775 => "0000000010000000001001011100010100",
			776 => "0000000100000000001011100000010000",
			777 => "0000001110000000000100010100001000",
			778 => "0000001011000000000100010100000100",
			779 => "00000000000010110000110011011101",
			780 => "11111111010000110000110011011101",
			781 => "0000000110000000000001111000000100",
			782 => "00000001100000010000110011011101",
			783 => "11111111111010110000110011011101",
			784 => "00000001111011110000110011011101",
			785 => "0000001001000000001001111000001100",
			786 => "0000001010000000000001010000000100",
			787 => "11111101110110100000110011011101",
			788 => "0000000000000000000100010100000100",
			789 => "00000000001101000000110011011101",
			790 => "11111110101011110000110011011101",
			791 => "11111101111011000000110011011101",
			792 => "0000000111000000000111111000000100",
			793 => "00000001100110010000110011011101",
			794 => "0000001100000000001000111000100000",
			795 => "0000001010000000001001000100010000",
			796 => "0000001010000000001001000100001000",
			797 => "0000001110000000001000111100000100",
			798 => "11111111101100110000110011011101",
			799 => "00000000001101100000110011011101",
			800 => "0000000100000000001000110100000100",
			801 => "11111101100011010000110011011101",
			802 => "11111111100000100000110011011101",
			803 => "0000001000000000001011010100001000",
			804 => "0000001111000000001110101100000100",
			805 => "00000001000110000000110011011101",
			806 => "11111111110110010000110011011101",
			807 => "0000001010000000000110011000000100",
			808 => "11111111101110010000110011011101",
			809 => "00000000000111100000110011011101",
			810 => "0000000100000000001110111000010000",
			811 => "0000000100000000000011110000001000",
			812 => "0000001000000000001011010100000100",
			813 => "11111111110100000000110011011101",
			814 => "11111101110101110000110011011101",
			815 => "0000000000000000001110111100000100",
			816 => "00000000100010000000110011011101",
			817 => "11111110100100100000110011011101",
			818 => "0000001000000000000001110100000100",
			819 => "11111110000110010000110011011101",
			820 => "0000000000000000000100010100000100",
			821 => "00000000110101000000110011011101",
			822 => "11111110101001000000110011011101",
			823 => "0000000010000000000010110101100100",
			824 => "0000000010000000000001001000101000",
			825 => "0000000000000000001000110000011000",
			826 => "0000000011000000001101100000001100",
			827 => "0000000001000000000110000000000100",
			828 => "11111111100011010000111011011001",
			829 => "0000001110000000000000111000000100",
			830 => "00000000101100010000111011011001",
			831 => "00000010001011000000111011011001",
			832 => "0000001111000000001010011100000100",
			833 => "11111110100000110000111011011001",
			834 => "0000000100000000001110010000000100",
			835 => "00000000000000000000111011011001",
			836 => "00000000100001010000111011011001",
			837 => "0000001100000000001010000000001100",
			838 => "0000000111000000000111111000001000",
			839 => "0000000111000000001110111100000100",
			840 => "11111111111000010000111011011001",
			841 => "00000001001110100000111011011001",
			842 => "11111110111101000000111011011001",
			843 => "11111110010010110000111011011001",
			844 => "0000001010000000001000010100011000",
			845 => "0000000100000000001110100100010000",
			846 => "0000000011000000001000111100000100",
			847 => "11111110101000110000111011011001",
			848 => "0000000000000000001000110000001000",
			849 => "0000000010000000001110101100000100",
			850 => "11111111110011110000111011011001",
			851 => "00000001101001110000111011011001",
			852 => "00000001110111100000111011011001",
			853 => "0000000001000000001110100000000100",
			854 => "00000000010010100000111011011001",
			855 => "00000011101000100000111011011001",
			856 => "0000001010000000001001000100001000",
			857 => "0000000100000000000010110000000100",
			858 => "11111101110110010000111011011001",
			859 => "00000000000000000000111011011001",
			860 => "0000000110000000000001111000001100",
			861 => "0000001100000000001010000000001000",
			862 => "0000001100000000001010000000000100",
			863 => "11111111111111010000111011011001",
			864 => "00000001100111100000111011011001",
			865 => "11111110011001000000111011011001",
			866 => "0000001100000000001010000000001000",
			867 => "0000000001000000000000011000000100",
			868 => "00000000000001110000111011011001",
			869 => "11111110011111000000111011011001",
			870 => "0000000111000000000111111000000100",
			871 => "00000011010000010000111011011001",
			872 => "00000001000001110000111011011001",
			873 => "0000001110000000001111000101011000",
			874 => "0000001111000000000110100100100100",
			875 => "0000000011000000000111111000011000",
			876 => "0000000001000000000110000000010000",
			877 => "0000000011000000000011111100001000",
			878 => "0000001101000000000100000000000100",
			879 => "00000000000000000000111011011001",
			880 => "11111110100110010000111011011001",
			881 => "0000001010000000000110011100000100",
			882 => "11111111110010110000111011011001",
			883 => "00000010101000000000111011011001",
			884 => "0000000100000000001001001100000100",
			885 => "00000000000000000000111011011001",
			886 => "11111110011011000000111011011001",
			887 => "0000000011000000000111111000000100",
			888 => "00000010000111010000111011011001",
			889 => "0000000110000000001100011000000100",
			890 => "00000000000111010000111011011001",
			891 => "00000000000000000000111011011001",
			892 => "0000001110000000001000110000100000",
			893 => "0000001111000000001000011000010000",
			894 => "0000000110000000000001111000001000",
			895 => "0000001010000000001010110000000100",
			896 => "00000000000000000000111011011001",
			897 => "00000001000111100000111011011001",
			898 => "0000001110000000000111000100000100",
			899 => "00000000011010110000111011011001",
			900 => "11111110010110010000111011011001",
			901 => "0000000000000000001011000100001000",
			902 => "0000000000000000001110111100000100",
			903 => "00000000000000000000111011011001",
			904 => "00000010010111000000111011011001",
			905 => "0000000111000000001011000100000100",
			906 => "11111111011010010000111011011001",
			907 => "00000000111101110000111011011001",
			908 => "0000000001000000001110100000001100",
			909 => "0000001001000000001100110100001000",
			910 => "0000001111000000001111011100000100",
			911 => "00000001000001110000111011011001",
			912 => "11111110011010000000111011011001",
			913 => "11111110001000110000111011011001",
			914 => "0000000100000000001111100000000100",
			915 => "00000000011101100000111011011001",
			916 => "11111111011010100000111011011001",
			917 => "0000001111000000000110100100000100",
			918 => "00000001110011110000111011011001",
			919 => "0000001010000000001001000100100000",
			920 => "0000001010000000001000010100010000",
			921 => "0000000110000000001100011000001000",
			922 => "0000000000000000000010111100000100",
			923 => "11111111101111000000111011011001",
			924 => "00000000101001010000111011011001",
			925 => "0000001100000000001000111000000100",
			926 => "00000001110111100000111011011001",
			927 => "00000000000000000000111011011001",
			928 => "0000000110000000001101111100001000",
			929 => "0000001000000000001001101000000100",
			930 => "00000001010010000000111011011001",
			931 => "11111111010010000000111011011001",
			932 => "0000001101000000000100001000000100",
			933 => "11111110000110010000111011011001",
			934 => "11111111110001010000111011011001",
			935 => "0000001100000000000100010100010000",
			936 => "0000000001000000001100110100001000",
			937 => "0000000111000000001011000100000100",
			938 => "00000000001010100000111011011001",
			939 => "11111111101001110000111011011001",
			940 => "0000001000000000000110001000000100",
			941 => "00000000000111010000111011011001",
			942 => "00000001000110110000111011011001",
			943 => "0000001100000000000100010100001000",
			944 => "0000000001000000001100110100000100",
			945 => "11111111111011100000111011011001",
			946 => "11111111000011010000111011011001",
			947 => "0000001100000000000100010100000100",
			948 => "00000000110010000000111011011001",
			949 => "11111111111110100000111011011001",
			950 => "0000000111000000001101111010000000",
			951 => "0000000100000000000011111001111100",
			952 => "0000000111000000000100010100111100",
			953 => "0000000011000000000000101000100000",
			954 => "0000001001000000001100110100010000",
			955 => "0000000011000000000000111000001000",
			956 => "0000000010000000001101000100000100",
			957 => "11111111010101100000111111111101",
			958 => "00000001110110100000111111111101",
			959 => "0000000110000000000111101000000100",
			960 => "11111110100101110000111111111101",
			961 => "00000010111000110000111111111101",
			962 => "0000000010000000001110101100001000",
			963 => "0000000011000000001110111100000100",
			964 => "00000000000010110000111111111101",
			965 => "00000010110010000000111111111101",
			966 => "0000001010000000000101000100000100",
			967 => "11111111000101010000111111111101",
			968 => "00000001010111100000111111111101",
			969 => "0000001010000000001001000100010000",
			970 => "0000000010000000000111100000001000",
			971 => "0000001011000000001011000100000100",
			972 => "11111111010011110000111111111101",
			973 => "00000010000101000000111111111101",
			974 => "0000001010000000001000010100000100",
			975 => "00000000000011010000111111111101",
			976 => "11111101010011010000111111111101",
			977 => "0000000010000000001110101000000100",
			978 => "00000100111111000000111111111101",
			979 => "0000001001000000000010001100000100",
			980 => "00000010000111110000111111111101",
			981 => "00000000111101000000111111111101",
			982 => "0000000110000000000100110100100000",
			983 => "0000000010000000001010001000010000",
			984 => "0000000111000000000100000000001000",
			985 => "0000001110000000000101101100000100",
			986 => "00000000010000100000111111111101",
			987 => "00000001010110100000111111111101",
			988 => "0000000100000000001000001000000100",
			989 => "11111111101110010000111111111101",
			990 => "11111101110001010000111111111101",
			991 => "0000001001000000001001111000001000",
			992 => "0000001000000000001111001000000100",
			993 => "11111111110110000000111111111101",
			994 => "00000011100100100000111111111101",
			995 => "0000001011000000001000111100000100",
			996 => "11111111000010100000111111111101",
			997 => "11111101111010110000111111111101",
			998 => "0000001001000000000110101000010000",
			999 => "0000001101000000001110001100001000",
			1000 => "0000000010000000001001010000000100",
			1001 => "00000001100110100000111111111101",
			1002 => "00000000010001110000111111111101",
			1003 => "0000001010000000000101000100000100",
			1004 => "00000010100010100000111111111101",
			1005 => "11111110011111110000111111111101",
			1006 => "0000000011000000001100101100001000",
			1007 => "0000001010000000000110011000000100",
			1008 => "11111100110000010000111111111101",
			1009 => "11111111011000100000111111111101",
			1010 => "0000001001000000000111100100000100",
			1011 => "00000001100011110000111111111101",
			1012 => "00000000010111100000111111111101",
			1013 => "11111110011001100000111111111101",
			1014 => "0000001010000000000111110100010000",
			1015 => "0000001111000000001000101000001100",
			1016 => "0000000111000000000001111100001000",
			1017 => "0000000110000000001011111100000100",
			1018 => "11111110101110100000111111111101",
			1019 => "00000001110011010000111111111101",
			1020 => "11111110011001010000111111111101",
			1021 => "00000011011100110000111111111101",
			1022 => "11111110011000110000111111111101",
			1023 => "0000001110000000001100110010101000",
			1024 => "0000001101000000000001111101110100",
			1025 => "0000001111000000000101110101000000",
			1026 => "0000001110000000000100000000100000",
			1027 => "0000001111000000000101100100010000",
			1028 => "0000000011000000001100001000001000",
			1029 => "0000001011000000000100010100000100",
			1030 => "00000000001100000001001000001001",
			1031 => "11111111100111110001001000001001",
			1032 => "0000001001000000001001111000000100",
			1033 => "00000001100011110001001000001001",
			1034 => "00000000001101100001001000001001",
			1035 => "0000000001000000001100110100001000",
			1036 => "0000001110000000000100010100000100",
			1037 => "11111111100111000001001000001001",
			1038 => "00000000001000000001001000001001",
			1039 => "0000001110000000001100001000000100",
			1040 => "11111111010111110001001000001001",
			1041 => "11111101010110100001001000001001",
			1042 => "0000000100000000001100001100010000",
			1043 => "0000001111000000000010001000001000",
			1044 => "0000000110000000000111101000000100",
			1045 => "11111110110111000001001000001001",
			1046 => "00000001001100010001001000001001",
			1047 => "0000000111000000001100001000000100",
			1048 => "00000000010000010001001000001001",
			1049 => "11111101110110110001001000001001",
			1050 => "0000001100000000000000101000001000",
			1051 => "0000000111000000000100000000000100",
			1052 => "00000001000001000001001000001001",
			1053 => "11111110111011010001001000001001",
			1054 => "0000001011000000001000111000000100",
			1055 => "00000010110111010001001000001001",
			1056 => "00000000100111100001001000001001",
			1057 => "0000001100000000000000101000100000",
			1058 => "0000001100000000001110111100010000",
			1059 => "0000001100000000001010000000001000",
			1060 => "0000001111000000000000110100000100",
			1061 => "11111111010000000001001000001001",
			1062 => "00000001101010100001001000001001",
			1063 => "0000000110000000001100011000000100",
			1064 => "00000010010001100001001000001001",
			1065 => "00000000101010100001001000001001",
			1066 => "0000001000000000001011010100001000",
			1067 => "0000001101000000001100101100000100",
			1068 => "11111101111011110001001000001001",
			1069 => "11111111101001110001001000001001",
			1070 => "0000000000000000000011010000000100",
			1071 => "00000010010111000001001000001001",
			1072 => "11111111110000000001001000001001",
			1073 => "0000001100000000000000101000000100",
			1074 => "00000100000100000001001000001001",
			1075 => "0000001100000000000100000000001000",
			1076 => "0000001111000000000111110000000100",
			1077 => "11111111010000000001001000001001",
			1078 => "11111101111110000001001000001001",
			1079 => "0000001110000000001000111000000100",
			1080 => "11111111010101110001001000001001",
			1081 => "00000001000010000001001000001001",
			1082 => "0000001100000000001000111000100100",
			1083 => "0000001111000000000000110100011100",
			1084 => "0000000011000000000100001000010000",
			1085 => "0000001110000000001100001000001000",
			1086 => "0000001110000000000000101000000100",
			1087 => "11111111010100000001001000001001",
			1088 => "00000000001011000001001000001001",
			1089 => "0000001100000000000100000000000100",
			1090 => "11111101011001000001001000001001",
			1091 => "11111110100010100001001000001001",
			1092 => "0000000111000000000100000000000100",
			1093 => "00000001000000110001001000001001",
			1094 => "0000001110000000000011011100000100",
			1095 => "11111111100101010001001000001001",
			1096 => "11111101110011010001001000001001",
			1097 => "0000001001000000001011101000000100",
			1098 => "00000000010100000001001000001001",
			1099 => "00000010110010010001001000001001",
			1100 => "0000001111000000000111110000001000",
			1101 => "0000000010000000000110100000000100",
			1102 => "00000001100100110001001000001001",
			1103 => "11111110110111010001001000001001",
			1104 => "0000001110000000000011011100000100",
			1105 => "00000101110111100001001000001001",
			1106 => "11111111110010110001001000001001",
			1107 => "0000001101000000000000001100100000",
			1108 => "0000000010000000000110010000010100",
			1109 => "0000000001000000001110100000000100",
			1110 => "11111101010001100001001000001001",
			1111 => "0000000111000000000100010100000100",
			1112 => "11111111101101000001001000001001",
			1113 => "0000001011000000001000111100001000",
			1114 => "0000001011000000000100000000000100",
			1115 => "00000001010111100001001000001001",
			1116 => "11111111101110010001001000001001",
			1117 => "00000010100100000001001000001001",
			1118 => "0000001111000000001100100100001000",
			1119 => "0000000111000000001100001000000100",
			1120 => "00000001011111100001001000001001",
			1121 => "11111110100110100001001000001001",
			1122 => "11111110000010000001001000001001",
			1123 => "0000000011000000000000001100001100",
			1124 => "0000001011000000000100000000000100",
			1125 => "00000000100110100001001000001001",
			1126 => "0000000001000000000010001100000100",
			1127 => "11111100100101010001001000001001",
			1128 => "00000000011000110001001000001001",
			1129 => "0000001000000000001010101100011000",
			1130 => "0000000100000000000010100100010000",
			1131 => "0000000000000000001111000100001000",
			1132 => "0000000100000000001000110100000100",
			1133 => "11111111111110100001001000001001",
			1134 => "11111110101101110001001000001001",
			1135 => "0000001000000000001001101000000100",
			1136 => "00000001011000000001001000001001",
			1137 => "00000000001000110001001000001001",
			1138 => "0000001101000000000100001000000100",
			1139 => "00000000000000000001001000001001",
			1140 => "11111110010000000001001000001001",
			1141 => "0000001100000000000100000000001100",
			1142 => "0000001111000000001110101100000100",
			1143 => "00000110111110110001001000001001",
			1144 => "0000001111000000001100100100000100",
			1145 => "11111111000010100001001000001001",
			1146 => "00000010101000110001001000001001",
			1147 => "0000001110000000000110100100001000",
			1148 => "0000000111000000001000111000000100",
			1149 => "00000000011110000001001000001001",
			1150 => "11111110100101010001001000001001",
			1151 => "0000000110000000001000010000000100",
			1152 => "00000010010010000001001000001001",
			1153 => "11111111001000110001001000001001",
			1154 => "0000001100000000000110000110101100",
			1155 => "0000001001000000001001111001011000",
			1156 => "0000000011000000001000111100111100",
			1157 => "0000001000000000000110001000100000",
			1158 => "0000000100000000000010111000010000",
			1159 => "0000001100000000000111111000001000",
			1160 => "0000001000000000001011010100000100",
			1161 => "00000001101101100001001101110101",
			1162 => "11111111011111110001001101110101",
			1163 => "0000001110000000000011010000000100",
			1164 => "11111110011100010001001101110101",
			1165 => "00000000001011010001001101110101",
			1166 => "0000000101000000001001110000001000",
			1167 => "0000000010000000001110101000000100",
			1168 => "00000000111100010001001101110101",
			1169 => "11111110111011010001001101110101",
			1170 => "0000000101000000000011011100000100",
			1171 => "00000100011100000001001101110101",
			1172 => "00000000011110000001001101110101",
			1173 => "0000000101000000001100110000010000",
			1174 => "0000001001000000000010001100001000",
			1175 => "0000000011000000001010000000000100",
			1176 => "11111111101100010001001101110101",
			1177 => "00000000110111010001001101110101",
			1178 => "0000001000000000001111001000000100",
			1179 => "11111110010111110001001101110101",
			1180 => "11111111101001100001001101110101",
			1181 => "0000001000000000000010101000000100",
			1182 => "00000101000011110001001101110101",
			1183 => "0000001101000000001100101100000100",
			1184 => "11111111100000000001001101110101",
			1185 => "00000010101110110001001101110101",
			1186 => "0000001011000000001100001000011000",
			1187 => "0000000010000000000010011100001100",
			1188 => "0000000000000000000010011000000100",
			1189 => "11111110111100010001001101110101",
			1190 => "0000001000000000000110001000000100",
			1191 => "00000011110011000001001101110101",
			1192 => "00000001101011000001001101110101",
			1193 => "0000000000000000000000111000000100",
			1194 => "11111110000110100001001101110101",
			1195 => "0000000101000000001100110000000100",
			1196 => "00000000100110100001001101110101",
			1197 => "00000010001000010001001101110101",
			1198 => "11111101111101100001001101110101",
			1199 => "0000000001000000001110100000011000",
			1200 => "0000000101000000000011011100000100",
			1201 => "00000000101001100001001101110101",
			1202 => "0000000001000000001110100000001000",
			1203 => "0000001110000000000111111000000100",
			1204 => "11111110011100010001001101110101",
			1205 => "11111100110100100001001101110101",
			1206 => "0000001110000000000100010100001000",
			1207 => "0000000000000000000100010100000100",
			1208 => "11111101111110100001001101110101",
			1209 => "11111111110000000001001101110101",
			1210 => "00000000100100010001001101110101",
			1211 => "0000001100000000000111111000100000",
			1212 => "0000001001000000001001111000010000",
			1213 => "0000000101000000001101100000001000",
			1214 => "0000001100000000000111111000000100",
			1215 => "00000000101010000001001101110101",
			1216 => "11111110001110110001001101110101",
			1217 => "0000001000000000001111001000000100",
			1218 => "00000010110001000001001101110101",
			1219 => "00000001101010110001001101110101",
			1220 => "0000000010000000000011001000001000",
			1221 => "0000000010000000000100101000000100",
			1222 => "11111111110111010001001101110101",
			1223 => "11111111000011110001001101110101",
			1224 => "0000000101000000001101100000000100",
			1225 => "00000010100110010001001101110101",
			1226 => "11111111111001110001001101110101",
			1227 => "0000001100000000000100010100010000",
			1228 => "0000000101000000001110001100001000",
			1229 => "0000001001000000000110101000000100",
			1230 => "00000000100001000001001101110101",
			1231 => "00000010000100100001001101110101",
			1232 => "0000001011000000001000111100000100",
			1233 => "11111110011001100001001101110101",
			1234 => "00000001100101010001001101110101",
			1235 => "0000000101000000000011011100000100",
			1236 => "00000010011100100001001101110101",
			1237 => "0000001011000000001011000100000100",
			1238 => "11111110110111110001001101110101",
			1239 => "00000000000100110001001101110101",
			1240 => "0000001010000000000111110100001000",
			1241 => "0000000010000000000001011100000100",
			1242 => "11111110100011110001001101110101",
			1243 => "00000001011101010001001101110101",
			1244 => "11111110011100100001001101110101",
			1245 => "0000001000000000001001101010001100",
			1246 => "0000001000000000001001101001000000",
			1247 => "0000001101000000000101101100100100",
			1248 => "0000000111000000000100010100010100",
			1249 => "0000000110000000000001111000010000",
			1250 => "0000001110000000001110111100001000",
			1251 => "0000001011000000000100010100000100",
			1252 => "00000000110110100001010110100001",
			1253 => "11111110110101100001010110100001",
			1254 => "0000000100000000001110000000000100",
			1255 => "11111111011001110001010110100001",
			1256 => "00000010000101100001010110100001",
			1257 => "11111110111010010001010110100001",
			1258 => "0000000010000000001101000100001100",
			1259 => "0000000011000000000100010100000100",
			1260 => "00000000000010010001010110100001",
			1261 => "0000000010000000000010110100000100",
			1262 => "00000010111010000001010110100001",
			1263 => "00000001011010100001010110100001",
			1264 => "11111111100010110001010110100001",
			1265 => "0000001110000000000000110000000100",
			1266 => "11111110010011110001010110100001",
			1267 => "0000000111000000000100010100001000",
			1268 => "0000000001000000001110100000000100",
			1269 => "11111111110110010001010110100001",
			1270 => "00000010100000000001010110100001",
			1271 => "0000001011000000000000101000001000",
			1272 => "0000000100000000000110001100000100",
			1273 => "11111110011110110001010110100001",
			1274 => "00000000011110000001010110100001",
			1275 => "0000000101000000001100101100000100",
			1276 => "00000000101010110001010110100001",
			1277 => "11111111111100010001010110100001",
			1278 => "0000000010000000000010011100101000",
			1279 => "0000001010000000001000010100010000",
			1280 => "0000001010000000001000010100000100",
			1281 => "00000000001111110001010110100001",
			1282 => "0000000110000000000001111000001000",
			1283 => "0000001011000000001100001000000100",
			1284 => "11111110100101100001010110100001",
			1285 => "00000000011100100001010110100001",
			1286 => "11111101101000000001010110100001",
			1287 => "0000000001000000001110100000001000",
			1288 => "0000001001000000001001111000000100",
			1289 => "11111111101100000001010110100001",
			1290 => "11111110001101010001010110100001",
			1291 => "0000000101000000001101111000001000",
			1292 => "0000001100000000000000101000000100",
			1293 => "00000000100010100001010110100001",
			1294 => "00000010100000100001010110100001",
			1295 => "0000000101000000000000001100000100",
			1296 => "11111110011011110001010110100001",
			1297 => "00000000011101010001010110100001",
			1298 => "0000001011000000000100010100001000",
			1299 => "0000001100000000000000111000000100",
			1300 => "00000000000000000001010110100001",
			1301 => "00000010100011010001010110100001",
			1302 => "0000000001000000001100110100001100",
			1303 => "0000000111000000001011000100000100",
			1304 => "11111101001101000001010110100001",
			1305 => "0000001110000000001000111100000100",
			1306 => "11111101111111110001010110100001",
			1307 => "11111111101101000001010110100001",
			1308 => "0000001101000000000000001100001000",
			1309 => "0000000001000000001100110100000100",
			1310 => "00000000010101000001010110100001",
			1311 => "00000010001010100001010110100001",
			1312 => "0000000001000000001001111000000100",
			1313 => "11111110011100100001010110100001",
			1314 => "00000000000001100001010110100001",
			1315 => "0000001000000000001011010100110100",
			1316 => "0000000110000000001010011000101000",
			1317 => "0000000100000000001000001000010100",
			1318 => "0000001101000000001110001100001100",
			1319 => "0000001011000000000000101000000100",
			1320 => "00000001010011110001010110100001",
			1321 => "0000000100000000000110001100000100",
			1322 => "00000001000110100001010110100001",
			1323 => "11111110110011110001010110100001",
			1324 => "0000000010000000001010001000000100",
			1325 => "00000010000100100001010110100001",
			1326 => "00000001000110000001010110100001",
			1327 => "0000000010000000000101110000001100",
			1328 => "0000000100000000000011001100000100",
			1329 => "00000000001100000001010110100001",
			1330 => "0000000110000000000001111000000100",
			1331 => "00000000100110000001010110100001",
			1332 => "00000010101011000001010110100001",
			1333 => "0000000111000000000100010100000100",
			1334 => "00000001101001010001010110100001",
			1335 => "11111110000111010001010110100001",
			1336 => "0000000010000000001111010100000100",
			1337 => "11111101101010000001010110100001",
			1338 => "0000000011000000001101000100000100",
			1339 => "00000010000111110001010110100001",
			1340 => "00000000000000000001010110100001",
			1341 => "0000000101000000000100011001000000",
			1342 => "0000001001000000001011101000100000",
			1343 => "0000000001000000000010001100010000",
			1344 => "0000000010000000000010000000001000",
			1345 => "0000000011000000001101111000000100",
			1346 => "00000000000011100001010110100001",
			1347 => "00000000011111000001010110100001",
			1348 => "0000000111000000000100000000000100",
			1349 => "11111111010111100001010110100001",
			1350 => "00000000101010010001010110100001",
			1351 => "0000001011000000000100000000001000",
			1352 => "0000001001000000001101101000000100",
			1353 => "11111101011010100001010110100001",
			1354 => "00000000010010000001010110100001",
			1355 => "0000001001000000001101101000000100",
			1356 => "00000010010111010001010110100001",
			1357 => "00000000100101010001010110100001",
			1358 => "0000001110000000001101010100010000",
			1359 => "0000001100000000001000111000001000",
			1360 => "0000001000000000001011010100000100",
			1361 => "11111101000110010001010110100001",
			1362 => "11111111010100010001010110100001",
			1363 => "0000000100000000001110111000000100",
			1364 => "00000001101100100001010110100001",
			1365 => "11111110101100100001010110100001",
			1366 => "0000001001000000001111001100001000",
			1367 => "0000000110000000001010011000000100",
			1368 => "11111111111100010001010110100001",
			1369 => "00000001010001010001010110100001",
			1370 => "0000001010000000000001010000000100",
			1371 => "00000000111011010001010110100001",
			1372 => "11111111000010000001010110100001",
			1373 => "0000000100000000000010100100010100",
			1374 => "0000001110000000001101010100000100",
			1375 => "00000011010111110001010110100001",
			1376 => "0000000100000000001000001000001000",
			1377 => "0000000111000000001001110000000100",
			1378 => "00000001110000000001010110100001",
			1379 => "11111111000100000001010110100001",
			1380 => "0000001100000000000100000000000100",
			1381 => "11111111010110110001010110100001",
			1382 => "00000001010111000001010110100001",
			1383 => "11111110011111110001010110100001",
			1384 => "0000000101000000000011100010110000",
			1385 => "0000000100000000000011010101100000",
			1386 => "0000001110000000000100010100110000",
			1387 => "0000001110000000001010000000010100",
			1388 => "0000000100000000000111010100000100",
			1389 => "00000110011000010001011101110101",
			1390 => "0000000110000000001101111100001000",
			1391 => "0000001011000000000100010100000100",
			1392 => "00000001001100110001011101110101",
			1393 => "11111111101111110001011101110101",
			1394 => "0000000000000000000100010100000100",
			1395 => "00000011000000100001011101110101",
			1396 => "11111110111010000001011101110101",
			1397 => "0000001000000000001100000100001100",
			1398 => "0000000110000000000001111000001000",
			1399 => "0000000101000000000101101100000100",
			1400 => "00000000100100010001011101110101",
			1401 => "11111110011100100001011101110101",
			1402 => "00000011010000000001011101110101",
			1403 => "0000000010000000001110101000001000",
			1404 => "0000000000000000000010111100000100",
			1405 => "00000010100010110001011101110101",
			1406 => "00000111000101010001011101110101",
			1407 => "0000001001000000001001111000000100",
			1408 => "00000100010101110001011101110101",
			1409 => "00000001011001010001011101110101",
			1410 => "0000000110000000000111101000010000",
			1411 => "0000001000000000000001010100001100",
			1412 => "0000000011000000001101100000000100",
			1413 => "11111111111100110001011101110101",
			1414 => "0000001100000000000111111000000100",
			1415 => "11111110111011110001011101110101",
			1416 => "11111110010001000001011101110101",
			1417 => "00000010101011010001011101110101",
			1418 => "0000000100000000001010110100010000",
			1419 => "0000000110000000001001100100001000",
			1420 => "0000000110000000001101111100000100",
			1421 => "00000010111100010001011101110101",
			1422 => "00000100101110000001011101110101",
			1423 => "0000001010000000001100011100000100",
			1424 => "11111110001100010001011101110101",
			1425 => "00000001010101000001011101110101",
			1426 => "0000001100000000000100000000001000",
			1427 => "0000001110000000001100110000000100",
			1428 => "00000010010011010001011101110101",
			1429 => "00000011111011100001011101110101",
			1430 => "0000000010000000001100010000000100",
			1431 => "11111111110101000001011101110101",
			1432 => "00000010110001010001011101110101",
			1433 => "0000000110000000001101111100010100",
			1434 => "0000000100000000000011110100000100",
			1435 => "00000010010101010001011101110101",
			1436 => "0000000001000000000000011000000100",
			1437 => "11111110001110100001011101110101",
			1438 => "0000001001000000000010001100001000",
			1439 => "0000000100000000000011101100000100",
			1440 => "11111110011110000001011101110101",
			1441 => "00000000011101110001011101110101",
			1442 => "11111110011000110001011101110101",
			1443 => "0000001011000000001100001000100000",
			1444 => "0000000000000000001011000100010000",
			1445 => "0000001100000000000111111000001000",
			1446 => "0000000100000000000011110100000100",
			1447 => "00000011111000110001011101110101",
			1448 => "00000111101001000001011101110101",
			1449 => "0000000101000000000101101100000100",
			1450 => "00000010100110010001011101110101",
			1451 => "11111111001111110001011101110101",
			1452 => "0000000100000000000001101100001000",
			1453 => "0000001001000000001100110100000100",
			1454 => "00000011000000010001011101110101",
			1455 => "00000000001010000001011101110101",
			1456 => "0000001010000000001100000100000100",
			1457 => "00000100101001000001011101110101",
			1458 => "11111110010000100001011101110101",
			1459 => "0000001111000000001100100100010000",
			1460 => "0000000010000000001001011100001000",
			1461 => "0000000011000000000101101100000100",
			1462 => "11111111100110110001011101110101",
			1463 => "00000011111000100001011101110101",
			1464 => "0000001100000000000111111000000100",
			1465 => "00000001100010000001011101110101",
			1466 => "11111110111001100001011101110101",
			1467 => "0000000000000000000100010100000100",
			1468 => "11111110001101100001011101110101",
			1469 => "0000000100000000000011101100000100",
			1470 => "00000011101011110001011101110101",
			1471 => "11111111010111010001011101110101",
			1472 => "0000001100000000000110000100100100",
			1473 => "0000000101000000000100010000100000",
			1474 => "0000000011000000001000011000000100",
			1475 => "11111110010011110001011101110101",
			1476 => "0000000110000000001101011000001100",
			1477 => "0000000110000000000001111000000100",
			1478 => "11111110010110000001011101110101",
			1479 => "0000000010000000001100010100000100",
			1480 => "00000101110010100001011101110101",
			1481 => "00000001111000000001011101110101",
			1482 => "0000000110000000001001100100001000",
			1483 => "0000000010000000001100010000000100",
			1484 => "11111110111001000001011101110101",
			1485 => "00000000110001010001011101110101",
			1486 => "0000001100000000001100001000000100",
			1487 => "11111111011010100001011101110101",
			1488 => "11111110010010110001011101110101",
			1489 => "00000101110001100001011101110101",
			1490 => "0000001100000000000110000100010100",
			1491 => "0000001000000000001111001000010000",
			1492 => "0000001000000000000110001000001100",
			1493 => "0000001000000000000110011100000100",
			1494 => "11111110011000110001011101110101",
			1495 => "0000001000000000001100000100000100",
			1496 => "00000000100110000001011101110101",
			1497 => "11111110100011010001011101110101",
			1498 => "00000001111011100001011101110101",
			1499 => "11111110010011100001011101110101",
			1500 => "11111110001110100001011101110101",
			1501 => "0000000010000000001100010110001100",
			1502 => "0000000100000000000011011001100000",
			1503 => "0000000110000000001010011001000000",
			1504 => "0000000110000000001100011000100000",
			1505 => "0000000110000000001100011000010000",
			1506 => "0000000010000000001110101000001000",
			1507 => "0000000110000000000001111000000100",
			1508 => "00000000000000100001100110011001",
			1509 => "00000000101111010001100110011001",
			1510 => "0000000110000000001101111100000100",
			1511 => "11111111101101110001100110011001",
			1512 => "00000000000100110001100110011001",
			1513 => "0000000100000000000011001100001000",
			1514 => "0000000001000000001100110100000100",
			1515 => "11111110111101010001100110011001",
			1516 => "00000000110001010001100110011001",
			1517 => "0000001000000000001111001000000100",
			1518 => "11111101010011000001100110011001",
			1519 => "11111111100001000001100110011001",
			1520 => "0000000011000000001101111000010000",
			1521 => "0000000001000000001100110100001000",
			1522 => "0000000011000000001100101100000100",
			1523 => "00000000001011010001100110011001",
			1524 => "00000001010000110001100110011001",
			1525 => "0000001000000000000001110100000100",
			1526 => "11111101110000010001100110011001",
			1527 => "00000000001011010001100110011001",
			1528 => "0000001100000000000100000000001000",
			1529 => "0000001110000000001001110000000100",
			1530 => "00000000010000100001100110011001",
			1531 => "00000001001010010001100110011001",
			1532 => "0000000110000000001010011000000100",
			1533 => "00000000100001010001100110011001",
			1534 => "11111110011111010001100110011001",
			1535 => "0000001000000000001011010100001100",
			1536 => "0000001100000000001000111000001000",
			1537 => "0000001000000000001001101000000100",
			1538 => "11111111000011000001100110011001",
			1539 => "11111011110100010001100110011001",
			1540 => "00000000100100000001100110011001",
			1541 => "0000001010000000000001010000000100",
			1542 => "00000011010111100001100110011001",
			1543 => "0000000111000000000100000000001000",
			1544 => "0000000010000000000011001000000100",
			1545 => "11111111100010110001100110011001",
			1546 => "00000001111100100001100110011001",
			1547 => "0000001101000000001100101000000100",
			1548 => "00000001010110000001100110011001",
			1549 => "11111110111110100001100110011001",
			1550 => "0000000001000000001110100000100100",
			1551 => "0000001101000000000110000100011100",
			1552 => "0000000000000000001100110000010000",
			1553 => "0000000011000000001110111100001000",
			1554 => "0000001010000000000101000100000100",
			1555 => "11111111001101010001100110011001",
			1556 => "00000001111100010001100110011001",
			1557 => "0000000110000000000001111000000100",
			1558 => "00000000000000000001100110011001",
			1559 => "00000011000100110001100110011001",
			1560 => "0000000100000000000110110000000100",
			1561 => "11111110010001110001100110011001",
			1562 => "0000000100000000000011111000000100",
			1563 => "00000001010001000001100110011001",
			1564 => "11111110101000100001100110011001",
			1565 => "0000001110000000000011111100000100",
			1566 => "11111110010100010001100110011001",
			1567 => "11111111111111010001100110011001",
			1568 => "0000001100000000000000101000000100",
			1569 => "00000110101110100001100110011001",
			1570 => "11111110111000110001100110011001",
			1571 => "0000000110000000001100011001001100",
			1572 => "0000001111000000001110101000101000",
			1573 => "0000001110000000001101111000100000",
			1574 => "0000000000000000000000110000010000",
			1575 => "0000001011000000000000101000001000",
			1576 => "0000001100000000001010000000000100",
			1577 => "00000000000000000001100110011001",
			1578 => "00000000111001100001100110011001",
			1579 => "0000000111000000001100001000000100",
			1580 => "11111101001010110001100110011001",
			1581 => "11111110011011100001100110011001",
			1582 => "0000000111000000001100001000001000",
			1583 => "0000001101000000001100101100000100",
			1584 => "11111111011010000001100110011001",
			1585 => "00000001000101100001100110011001",
			1586 => "0000000111000000000100000000000100",
			1587 => "11111110000100100001100110011001",
			1588 => "00000000001001000001100110011001",
			1589 => "0000000001000000000010001100000100",
			1590 => "00000010000110010001100110011001",
			1591 => "11111111001110110001100110011001",
			1592 => "0000001110000000000011011100000100",
			1593 => "00000100011111010001100110011001",
			1594 => "0000001101000000001010111000010000",
			1595 => "0000001100000000000000101000001000",
			1596 => "0000001000000000001100000100000100",
			1597 => "00000001110100000001100110011001",
			1598 => "11111110010000000001100110011001",
			1599 => "0000000000000000000000110000000100",
			1600 => "11111100100110000001100110011001",
			1601 => "11111101110001010001100110011001",
			1602 => "0000000110000000001100011000001000",
			1603 => "0000000100000000000001011100000100",
			1604 => "11111111111100010001100110011001",
			1605 => "11111110010110000001100110011001",
			1606 => "0000000010000000001110110100000100",
			1607 => "00000001100111100001100110011001",
			1608 => "11111111001011010001100110011001",
			1609 => "0000000110000000001111000000110000",
			1610 => "0000001111000000000000110100010000",
			1611 => "0000000110000000001010011000001000",
			1612 => "0000000011000000001110001100000100",
			1613 => "11111110100000100001100110011001",
			1614 => "00000001100110000001100110011001",
			1615 => "0000000001000000000010001100000100",
			1616 => "11111110001001100001100110011001",
			1617 => "00000000000000000001100110011001",
			1618 => "0000001000000000001111001000010000",
			1619 => "0000000100000000001000001000001000",
			1620 => "0000001101000000001010111000000100",
			1621 => "00000001111100010001100110011001",
			1622 => "11111111110011110001100110011001",
			1623 => "0000000010000000000010000000000100",
			1624 => "00000000101101110001100110011001",
			1625 => "11111110011111110001100110011001",
			1626 => "0000000100000000001110111000001000",
			1627 => "0000001111000000000101110000000100",
			1628 => "00000000100101010001100110011001",
			1629 => "00000010001010000001100110011001",
			1630 => "0000000000000000001110111100000100",
			1631 => "11111111000110100001100110011001",
			1632 => "00000000010001100001100110011001",
			1633 => "0000001101000000001011000000001000",
			1634 => "0000000010000000001111010100000100",
			1635 => "11111111011011000001100110011001",
			1636 => "00000001001111010001100110011001",
			1637 => "11111110010110110001100110011001",
			1638 => "0000001100000000000100000010101100",
			1639 => "0000001100000000000000101001110000",
			1640 => "0000000010000000000110010000111000",
			1641 => "0000000001000000000010001100100000",
			1642 => "0000000111000000001100001000010000",
			1643 => "0000000111000000000000101000001000",
			1644 => "0000000111000000000000101000000100",
			1645 => "00000000000011100001110000001101",
			1646 => "11111111010101110001110000001101",
			1647 => "0000001110000000001101111000000100",
			1648 => "00000000010000110001110000001101",
			1649 => "00000001100110010001110000001101",
			1650 => "0000000111000000001100001000001000",
			1651 => "0000001010000000001100011100000100",
			1652 => "11111110100110000001110000001101",
			1653 => "00000000111100100001110000001101",
			1654 => "0000001000000000000001110100000100",
			1655 => "11111111111001110001110000001101",
			1656 => "00000000111110010001110000001101",
			1657 => "0000001001000000001101011100010000",
			1658 => "0000000111000000001000111000001000",
			1659 => "0000000100000000001000101000000100",
			1660 => "11111111010101110001110000001101",
			1661 => "00000001010001010001110000001101",
			1662 => "0000001010000000000001010000000100",
			1663 => "11111110101001000001110000001101",
			1664 => "00000000111010010001110000001101",
			1665 => "0000001110000000001000000000000100",
			1666 => "11111110000101010001110000001101",
			1667 => "00000000000101010001110000001101",
			1668 => "0000001001000000001101101000100000",
			1669 => "0000001111000000001101000100010000",
			1670 => "0000001010000000001100011100001000",
			1671 => "0000001000000000000110001000000100",
			1672 => "00000000110110010001110000001101",
			1673 => "11111110011010010001110000001101",
			1674 => "0000001110000000001000111100000100",
			1675 => "11111110100101000001110000001101",
			1676 => "00000000100001000001110000001101",
			1677 => "0000001111000000001110000100001000",
			1678 => "0000001100000000000100010100000100",
			1679 => "11111111110100010001110000001101",
			1680 => "00000001100100110001110000001101",
			1681 => "0000001111000000000010011100000100",
			1682 => "11111110010000010001110000001101",
			1683 => "00000000000000000001110000001101",
			1684 => "0000000100000000000010110000001000",
			1685 => "0000000100000000000110001100000100",
			1686 => "11111110111110000001110000001101",
			1687 => "00000001100110110001110000001101",
			1688 => "0000001000000000000111000100001000",
			1689 => "0000000001000000001001111000000100",
			1690 => "11111101111101110001110000001101",
			1691 => "00000000000000000001110000001101",
			1692 => "0000000100000000000100001100000100",
			1693 => "00000000001111110001110000001101",
			1694 => "11111110010011110001110000001101",
			1695 => "0000001100000000000000101000011000",
			1696 => "0000000100000000001101001000001100",
			1697 => "0000000011000000000000001100000100",
			1698 => "11111110101100110001110000001101",
			1699 => "0000001110000000000001111100000100",
			1700 => "00000001110111000001110000001101",
			1701 => "00000000010000000001110000001101",
			1702 => "0000001011000000001000111000001000",
			1703 => "0000001000000000000001110100000100",
			1704 => "00000011100000000001110000001101",
			1705 => "00000010001100100001110000001101",
			1706 => "00000000111000000001110000001101",
			1707 => "0000001000000000000001110000010000",
			1708 => "0000001010000000000111110100001000",
			1709 => "0000001001000000001111001100000100",
			1710 => "11111110100000110001110000001101",
			1711 => "00000001010111110001110000001101",
			1712 => "0000000001000000000010001100000100",
			1713 => "00000001000011000001110000001101",
			1714 => "00000010001010100001110000001101",
			1715 => "0000001010000000001000010100001000",
			1716 => "0000001010000000001000100100000100",
			1717 => "00000000011010000001110000001101",
			1718 => "11111100110000110001110000001101",
			1719 => "0000001010000000001000010100000100",
			1720 => "00000010001111100001110000001101",
			1721 => "0000001000000000001011010100000100",
			1722 => "11111111100010110001110000001101",
			1723 => "00000000010010000001110000001101",
			1724 => "0000001100000000000100000000111000",
			1725 => "0000000111000000000100000000001100",
			1726 => "0000000111000000000100000000000100",
			1727 => "11111110100000010001110000001101",
			1728 => "0000001111000000000001001000000100",
			1729 => "00000000011100110001110000001101",
			1730 => "00000010000011000001110000001101",
			1731 => "0000000001000000001001111000011000",
			1732 => "0000000010000000000110010000010000",
			1733 => "0000001001000000001101101000001000",
			1734 => "0000001011000000001000111000000100",
			1735 => "11111110010011000001110000001101",
			1736 => "11111100100101000001110000001101",
			1737 => "0000000001000000000010001100000100",
			1738 => "11111111101100010001110000001101",
			1739 => "11111101100010110001110000001101",
			1740 => "0000000101000000001100101000000100",
			1741 => "11111110010010110001110000001101",
			1742 => "00000000000000000001110000001101",
			1743 => "0000001110000000001110110000001000",
			1744 => "0000000111000000001001110000000100",
			1745 => "00000001110010000001110000001101",
			1746 => "11111111101101010001110000001101",
			1747 => "0000001111000000001001011100001000",
			1748 => "0000000000000000000010011000000100",
			1749 => "11111100111110010001110000001101",
			1750 => "11111110101111100001110000001101",
			1751 => "00000000100011000001110000001101",
			1752 => "0000001100000000000100000000011100",
			1753 => "0000000101000000000000001100001000",
			1754 => "0000000101000000001101111000000100",
			1755 => "00000001010000100001110000001101",
			1756 => "00000010101011000001110000001101",
			1757 => "0000000101000000000100001000000100",
			1758 => "11111110111101100001110000001101",
			1759 => "0000000101000000001010111000001000",
			1760 => "0000001110000000001100101000000100",
			1761 => "00000000101010110001110000001101",
			1762 => "00000010001110100001110000001101",
			1763 => "0000001111000000000100101000000100",
			1764 => "11111110010001000001110000001101",
			1765 => "00000000101110110001110000001101",
			1766 => "0000001100000000001000111100011100",
			1767 => "0000001100000000001000111100010000",
			1768 => "0000001110000000001010111000001000",
			1769 => "0000000111000000001000111000000100",
			1770 => "11111111111101010001110000001101",
			1771 => "11111110100011000001110000001101",
			1772 => "0000000010000000000110010000000100",
			1773 => "00000010001010000001110000001101",
			1774 => "11111110100001100001110000001101",
			1775 => "0000001110000000001110001100000100",
			1776 => "00000000000100000001110000001101",
			1777 => "0000000010000000001100000000000100",
			1778 => "11111101101100010001110000001101",
			1779 => "00000000001110000001110000001101",
			1780 => "0000001100000000001000111000010000",
			1781 => "0000000011000000000001011000001000",
			1782 => "0000001110000000000000001100000100",
			1783 => "11111111110111010001110000001101",
			1784 => "00000010000000110001110000001101",
			1785 => "0000000001000000001101101000000100",
			1786 => "11111110010111110001110000001101",
			1787 => "00000001000010110001110000001101",
			1788 => "0000001100000000001000111000001000",
			1789 => "0000000010000000001000001100000100",
			1790 => "11111110011011110001110000001101",
			1791 => "00000001100110010001110000001101",
			1792 => "0000000101000000001101010100000100",
			1793 => "00000000111011000001110000001101",
			1794 => "11111111111010110001110000001101",
			1795 => "0000001100000000001000111011011100",
			1796 => "0000001100000000000111111001110100",
			1797 => "0000001001000000000110101001000000",
			1798 => "0000000011000000001001110000100000",
			1799 => "0000001001000000001001111000010000",
			1800 => "0000000011000000001011000100001000",
			1801 => "0000001111000000000111010000000100",
			1802 => "11111111111111110001111001011001",
			1803 => "11111110011101100001111001011001",
			1804 => "0000000101000000000011011100000100",
			1805 => "00000000101110010001111001011001",
			1806 => "11111111101111000001111001011001",
			1807 => "0000000100000000000011110000001000",
			1808 => "0000001110000000000000110000000100",
			1809 => "11111111000111100001111001011001",
			1810 => "00000001110000000001111001011001",
			1811 => "0000001010000000000001010000000100",
			1812 => "11111110100010000001111001011001",
			1813 => "11111111101111110001111001011001",
			1814 => "0000001111000000000010001000010000",
			1815 => "0000001110000000000100010100001000",
			1816 => "0000000111000000000100010100000100",
			1817 => "11111111110100010001111001011001",
			1818 => "00000001101101100001111001011001",
			1819 => "0000000110000000000111101000000100",
			1820 => "00000000000000000001111001011001",
			1821 => "00000010011000000001111001011001",
			1822 => "0000001010000000000001010000001000",
			1823 => "0000001110000000000100000000000100",
			1824 => "11111110111001100001111001011001",
			1825 => "00000000011100010001111001011001",
			1826 => "0000001010000000001100011100000100",
			1827 => "00000001010110110001111001011001",
			1828 => "11111110100010100001111001011001",
			1829 => "0000000101000000001100110000010100",
			1830 => "0000001011000000000000101000001100",
			1831 => "0000001100000000000111111000001000",
			1832 => "0000001110000000000000101000000100",
			1833 => "11111110000010100001111001011001",
			1834 => "11111111111111100001111001011001",
			1835 => "00000000111111010001111001011001",
			1836 => "0000001001000000000110101000000100",
			1837 => "11111110100011110001111001011001",
			1838 => "11111100100110100001111001011001",
			1839 => "0000001010000000001001000100010000",
			1840 => "0000000100000000001000110100001000",
			1841 => "0000001010000000001000100100000100",
			1842 => "11111111010110000001111001011001",
			1843 => "00000001010111000001111001011001",
			1844 => "0000000010000000000101001000000100",
			1845 => "11111101111111110001111001011001",
			1846 => "11111111011011010001111001011001",
			1847 => "0000001100000000000111111000001000",
			1848 => "0000000101000000001100101100000100",
			1849 => "00000001101010100001111001011001",
			1850 => "11111110111000000001111001011001",
			1851 => "0000000010000000000010011100000100",
			1852 => "00000000100101110001111001011001",
			1853 => "11111111011101000001111001011001",
			1854 => "0000001100000000000100010100101000",
			1855 => "0000000100000000001000001000010100",
			1856 => "0000001100000000000111111000001100",
			1857 => "0000000111000000000100010100000100",
			1858 => "00000001100010100001111001011001",
			1859 => "0000000111000000001100001000000100",
			1860 => "11111101110111110001111001011001",
			1861 => "00000000000000000001111001011001",
			1862 => "0000001001000000000110101000000100",
			1863 => "11111111111000010001111001011001",
			1864 => "00000010000010000001111001011001",
			1865 => "0000001011000000001110111100000100",
			1866 => "11111110010010000001111001011001",
			1867 => "0000000010000000000011001000001000",
			1868 => "0000001110000000000100010100000100",
			1869 => "00000001000000100001111001011001",
			1870 => "00000010100010100001111001011001",
			1871 => "0000001110000000001001110000000100",
			1872 => "11111110111000100001111001011001",
			1873 => "00000001010010010001111001011001",
			1874 => "0000000011000000001100110000100000",
			1875 => "0000001001000000000110101000010000",
			1876 => "0000001101000000001110001100001000",
			1877 => "0000000101000000000110000100000100",
			1878 => "11111111111111110001111001011001",
			1879 => "11111110111000000001111001011001",
			1880 => "0000001111000000000101100100000100",
			1881 => "00000001110010100001111001011001",
			1882 => "11111110110010100001111001011001",
			1883 => "0000001111000000000100000100001000",
			1884 => "0000000011000000001001110000000100",
			1885 => "11111110100001000001111001011001",
			1886 => "00000000101011010001111001011001",
			1887 => "0000000010000000001001010000000100",
			1888 => "11111101101011000001111001011001",
			1889 => "11111111101101110001111001011001",
			1890 => "0000001001000000000111100100010000",
			1891 => "0000001100000000000100010100001000",
			1892 => "0000001101000000000000001100000100",
			1893 => "00000000001111010001111001011001",
			1894 => "11111101011101100001111001011001",
			1895 => "0000000101000000000101101100000100",
			1896 => "00000010001001010001111001011001",
			1897 => "00000000100110110001111001011001",
			1898 => "0000001110000000001000111100001000",
			1899 => "0000001010000000000001010000000100",
			1900 => "11111111111100010001111001011001",
			1901 => "11111110111010010001111001011001",
			1902 => "0000001111000000001010010100000100",
			1903 => "00000000011011110001111001011001",
			1904 => "11111111111110100001111001011001",
			1905 => "0000001111000000001101000100011000",
			1906 => "0000000101000000001000000000001100",
			1907 => "0000001110000000000110000100001000",
			1908 => "0000000100000000001010110100000100",
			1909 => "00000001001000000001111001011001",
			1910 => "11111110011111110001111001011001",
			1911 => "11111101110111110001111001011001",
			1912 => "0000000101000000001000000000001000",
			1913 => "0000000110000000001100011000000100",
			1914 => "00000000000000000001111001011001",
			1915 => "00000011000000010001111001011001",
			1916 => "11111110110110100001111001011001",
			1917 => "0000000110000000001101011000011000",
			1918 => "0000000100000000001000001000010100",
			1919 => "0000000010000000000011001000001000",
			1920 => "0000000111000000000100001000000100",
			1921 => "00000001101100110001111001011001",
			1922 => "11111111101110010001111001011001",
			1923 => "0000001001000000001001100100000100",
			1924 => "11111110010111110001111001011001",
			1925 => "0000001010000000000010101100000100",
			1926 => "11111111001011110001111001011001",
			1927 => "00000001000010000001111001011001",
			1928 => "00000010111101100001111001011001",
			1929 => "0000001010000000000110011100010000",
			1930 => "0000001011000000001101111000000100",
			1931 => "11111110001100110001111001011001",
			1932 => "0000001001000000000101011100000100",
			1933 => "00000001001010010001111001011001",
			1934 => "0000000010000000001100000000000100",
			1935 => "11111111111100010001111001011001",
			1936 => "11111110100110100001111001011001",
			1937 => "0000001111000000000010011100001000",
			1938 => "0000000111000000000101101100000100",
			1939 => "00000100000111110001111001011001",
			1940 => "00000000000000000001111001011001",
			1941 => "11111110101100010001111001011001",
			1942 => "0000001001000000001001111010001000",
			1943 => "0000000101000000001101100001001000",
			1944 => "0000000101000000000011011101000000",
			1945 => "0000000010000000001001010000100000",
			1946 => "0000000011000000000100010100010000",
			1947 => "0000001011000000001011000100001000",
			1948 => "0000001010000000000101000100000100",
			1949 => "00000000000100100010000010111101",
			1950 => "00000001000100010010000010111101",
			1951 => "0000000110000000000001111000000100",
			1952 => "11111111111011000010000010111101",
			1953 => "11111110011101000010000010111101",
			1954 => "0000000111000000000111111000001000",
			1955 => "0000000011000000001100001000000100",
			1956 => "11111110110010100010000010111101",
			1957 => "11111111101101000010000010111101",
			1958 => "0000001011000000000100010100000100",
			1959 => "00000001110000110010000010111101",
			1960 => "00000000101100000010000010111101",
			1961 => "0000000001000000000110000000010000",
			1962 => "0000000011000000001100001000001000",
			1963 => "0000001100000000001010000000000100",
			1964 => "00000000100011100010000010111101",
			1965 => "11111110100011000010000010111101",
			1966 => "0000000011000000001100001000000100",
			1967 => "00000010000111100010000010111101",
			1968 => "00000000000001000010000010111101",
			1969 => "0000001011000000000100010100001000",
			1970 => "0000001000000000000001110100000100",
			1971 => "11111101111101100010000010111101",
			1972 => "11111111101010110010000010111101",
			1973 => "0000001100000000000111111000000100",
			1974 => "00000000110010000010000010111101",
			1975 => "11111110110000000010000010111101",
			1976 => "0000001111000000000110100100000100",
			1977 => "00000000010010010010000010111101",
			1978 => "11111110001111110010000010111101",
			1979 => "0000000110000000001101111100100100",
			1980 => "0000001101000000001101100000001100",
			1981 => "0000001100000000000100010100001000",
			1982 => "0000001000000000001011010100000100",
			1983 => "00000001001101100010000010111101",
			1984 => "11111110011111000010000010111101",
			1985 => "00000010010100010010000010111101",
			1986 => "0000000001000000000110000000010000",
			1987 => "0000001000000000001011010100001000",
			1988 => "0000000010000000000110100000000100",
			1989 => "11111111010110010010000010111101",
			1990 => "00000010001101000010000010111101",
			1991 => "0000000010000000000010000000000100",
			1992 => "11111110010110100010000010111101",
			1993 => "00000000001011100010000010111101",
			1994 => "0000001011000000001011000100000100",
			1995 => "11111110001110000010000010111101",
			1996 => "11111111011101010010000010111101",
			1997 => "0000000111000000001100001000011000",
			1998 => "0000001110000000000000111000001100",
			1999 => "0000001111000000000101100100001000",
			2000 => "0000000010000000001110000100000100",
			2001 => "00000000001000000010000010111101",
			2002 => "00000001100110100010000010111101",
			2003 => "11111110010100100010000010111101",
			2004 => "0000001101000000001101100000000100",
			2005 => "00000000010100110010000010111101",
			2006 => "0000001101000000000101101100000100",
			2007 => "00000010101001010010000010111101",
			2008 => "00000001011001100010000010111101",
			2009 => "11111110101011010010000010111101",
			2010 => "0000000011000000000101101101001100",
			2011 => "0000000011000000000101101100110100",
			2012 => "0000000011000000001100110000100000",
			2013 => "0000001001000000000111100100010000",
			2014 => "0000001100000000000111111000001000",
			2015 => "0000001011000000000000101000000100",
			2016 => "11111111110101000010000010111101",
			2017 => "11111110111110110010000010111101",
			2018 => "0000001100000000000100010100000100",
			2019 => "00000000010011010010000010111101",
			2020 => "11111111110100100010000010111101",
			2021 => "0000001001000000000111100100001000",
			2022 => "0000001010000000001010110000000100",
			2023 => "11111101111100010010000010111101",
			2024 => "11111111111101000010000010111101",
			2025 => "0000001111000000001011011100000100",
			2026 => "11111111111111000010000010111101",
			2027 => "11111110001111010010000010111101",
			2028 => "0000000110000000000100110100001100",
			2029 => "0000001100000000000100010100001000",
			2030 => "0000001100000000000100010100000100",
			2031 => "00000000010010000010000010111101",
			2032 => "11111110100101100010000010111101",
			2033 => "00000001010100000010000010111101",
			2034 => "0000000010000000001110010000000100",
			2035 => "00000010000000010010000010111101",
			2036 => "00000000101011110010000010111101",
			2037 => "0000001010000000000110011000001000",
			2038 => "0000000110000000000001111000000100",
			2039 => "11111110101001110010000010111101",
			2040 => "00000000011101110010000010111101",
			2041 => "0000001010000000001010110000001000",
			2042 => "0000001011000000001100001000000100",
			2043 => "11111110100000100010000010111101",
			2044 => "11111101100001000010000010111101",
			2045 => "0000000010000000001001011100000100",
			2046 => "00000000010101110010000010111101",
			2047 => "11111110010111100010000010111101",
			2048 => "0000001001000000000110101000110000",
			2049 => "0000001111000000000101110100010100",
			2050 => "0000001010000000001000010100001000",
			2051 => "0000001111000000001011011100000100",
			2052 => "00000000100101110010000010111101",
			2053 => "11111111101110000010000010111101",
			2054 => "0000001001000000000110101000000100",
			2055 => "00000000001000100010000010111101",
			2056 => "0000001011000000001100001000000100",
			2057 => "00000001010011000010000010111101",
			2058 => "00000010010010100010000010111101",
			2059 => "0000000101000000001100101100010000",
			2060 => "0000001100000000000111111000001000",
			2061 => "0000000011000000001100101100000100",
			2062 => "00000010001100010010000010111101",
			2063 => "00000000010011110010000010111101",
			2064 => "0000001100000000000100010100000100",
			2065 => "11111111110001000010000010111101",
			2066 => "00000001010001010010000010111101",
			2067 => "0000001001000000000110101000000100",
			2068 => "00000000000000000010000010111101",
			2069 => "0000001110000000001000111000000100",
			2070 => "11111101101010110010000010111101",
			2071 => "11111111010111100010000010111101",
			2072 => "0000001100000000000111111000010100",
			2073 => "0000001001000000000110101000000100",
			2074 => "11111110011001110010000010111101",
			2075 => "0000001111000000001010010100001000",
			2076 => "0000001101000000001110001100000100",
			2077 => "00000001110111000010000010111101",
			2078 => "11111111010001010010000010111101",
			2079 => "0000000010000000001110010000000100",
			2080 => "11111101111011110010000010111101",
			2081 => "00000000000000000010000010111101",
			2082 => "0000001100000000000111111000001100",
			2083 => "0000000111000000001011000100000100",
			2084 => "11111111010101010010000010111101",
			2085 => "0000000101000000001110001100000100",
			2086 => "00000000111101110010000010111101",
			2087 => "00000010100101010010000010111101",
			2088 => "0000000011000000001100101100001000",
			2089 => "0000000011000000001100101100000100",
			2090 => "11111111111100000010000010111101",
			2091 => "11111110101001010010000010111101",
			2092 => "0000001001000000000111100100000100",
			2093 => "00000000010100100010000010111101",
			2094 => "11111111111110100010000010111101",
			2095 => "0000001110000000000101101110100100",
			2096 => "0000001111000000000101100101010100",
			2097 => "0000000110000000000111101000100100",
			2098 => "0000001101000000001100101100011000",
			2099 => "0000000011000000001000111000010000",
			2100 => "0000000110000000000111101000001000",
			2101 => "0000001101000000001100110000000100",
			2102 => "00000001010111010010001101000001",
			2103 => "11111111011111110010001101000001",
			2104 => "0000000111000000000111111000000100",
			2105 => "00000001101011010010001101000001",
			2106 => "11111110110111010010001101000001",
			2107 => "0000001110000000001110111100000100",
			2108 => "00000000011001000010001101000001",
			2109 => "00000010010000100010001101000001",
			2110 => "0000001110000000001000111000000100",
			2111 => "11111110010001010010001101000001",
			2112 => "0000001110000000000011011100000100",
			2113 => "00000000000000000010001101000001",
			2114 => "11111111010001110010001101000001",
			2115 => "0000000011000000000101101100100000",
			2116 => "0000000010000000000010110100010000",
			2117 => "0000000010000000000000110100001000",
			2118 => "0000000111000000000100010100000100",
			2119 => "11111110011001110010001101000001",
			2120 => "00000000100111010010001101000001",
			2121 => "0000001111000000001001001000000100",
			2122 => "00000000011000000010001101000001",
			2123 => "00000010001001000010001101000001",
			2124 => "0000001001000000000111100100001000",
			2125 => "0000000011000000001101100000000100",
			2126 => "00000000000101100010001101000001",
			2127 => "00000001011110100010001101000001",
			2128 => "0000001111000000000100000100000100",
			2129 => "00000000100011100010001101000001",
			2130 => "11111110000011100010001101000001",
			2131 => "0000001101000000000001111100001100",
			2132 => "0000001001000000000110101000000100",
			2133 => "00000000000000110010001101000001",
			2134 => "0000000001000000001100110100000100",
			2135 => "00000001010101100010001101000001",
			2136 => "00000010011000100010001101000001",
			2137 => "11111111110111010010001101000001",
			2138 => "0000001001000000001011101000111100",
			2139 => "0000000011000000000011011100011100",
			2140 => "0000001001000000001001111000001100",
			2141 => "0000000111000000000000101000001000",
			2142 => "0000000011000000001000111000000100",
			2143 => "11111111110000010010001101000001",
			2144 => "00000000111100010010001101000001",
			2145 => "11111101111111110010001101000001",
			2146 => "0000000001000000001110100000001000",
			2147 => "0000001111000000000110110100000100",
			2148 => "11111111100101000010001101000001",
			2149 => "11111101111010000010001101000001",
			2150 => "0000001101000000001100101100000100",
			2151 => "00000000000110100010001101000001",
			2152 => "11111110101111000010001101000001",
			2153 => "0000001001000000000110101000010000",
			2154 => "0000001010000000000001010000001000",
			2155 => "0000000010000000001001010000000100",
			2156 => "00000000010110010010001101000001",
			2157 => "11111111011101110010001101000001",
			2158 => "0000000010000000000010000000000100",
			2159 => "00000000101001000010001101000001",
			2160 => "11111111101000110010001101000001",
			2161 => "0000000011000000000110000100001000",
			2162 => "0000001111000000000100010000000100",
			2163 => "11111111100000010010001101000001",
			2164 => "11111101111000000010001101000001",
			2165 => "0000001111000000001010010100000100",
			2166 => "00000000001010000010001101000001",
			2167 => "11111111100100100010001101000001",
			2168 => "0000000001000000000010001100000100",
			2169 => "11111101100001000010001101000001",
			2170 => "0000001111000000000000110100001000",
			2171 => "0000001110000000001100110000000100",
			2172 => "11111101111011100010001101000001",
			2173 => "11111111111010100010001101000001",
			2174 => "0000000010000000001011101100000100",
			2175 => "00000011010011100010001101000001",
			2176 => "00000000000000000010001101000001",
			2177 => "0000000000000000001111000101010100",
			2178 => "0000000100000000001011110000101100",
			2179 => "0000000000000000001101010000011100",
			2180 => "0000001000000000000001110000010000",
			2181 => "0000001010000000000111110100001000",
			2182 => "0000000100000000001011101100000100",
			2183 => "00000000001110000010001101000001",
			2184 => "11111110100000010010001101000001",
			2185 => "0000000111000000001000111000000100",
			2186 => "00000001111100010010001101000001",
			2187 => "11111111111100110010001101000001",
			2188 => "0000001001000000001011101000000100",
			2189 => "11111100111001110010001101000001",
			2190 => "0000001110000000000001101000000100",
			2191 => "00000000101110100010001101000001",
			2192 => "11111101111011110010001101000001",
			2193 => "0000000100000000000011000000000100",
			2194 => "11111110011000110010001101000001",
			2195 => "0000000101000000000000001100000100",
			2196 => "00000000001010010010001101000001",
			2197 => "0000000010000000001001100000000100",
			2198 => "00000010001111000010001101000001",
			2199 => "00000000000000000010001101000001",
			2200 => "0000000111000000001000111000010100",
			2201 => "0000000101000000001010111100010000",
			2202 => "0000000011000000001010111100001000",
			2203 => "0000001000000000000001110000000100",
			2204 => "11111110100001000010001101000001",
			2205 => "00000000100100010010001101000001",
			2206 => "0000001000000000001100000100000100",
			2207 => "11111110001101000010001101000001",
			2208 => "11111100010000010010001101000001",
			2209 => "00000000011111010010001101000001",
			2210 => "0000000101000000001101010100000100",
			2211 => "00000001101110100010001101000001",
			2212 => "0000000010000000000010000100001000",
			2213 => "0000000100000000001000000100000100",
			2214 => "11111111100000010010001101000001",
			2215 => "11111101100111100010001101000001",
			2216 => "0000000111000000000110100100000100",
			2217 => "00000000111000000010001101000001",
			2218 => "11111110111001000010001101000001",
			2219 => "0000001000000000001001101000010100",
			2220 => "0000000100000000000110001100001100",
			2221 => "0000000001000000000010001100001000",
			2222 => "0000001111000000001110101100000100",
			2223 => "00000001110101010010001101000001",
			2224 => "00000000010100010010001101000001",
			2225 => "00000010000110000010001101000001",
			2226 => "0000000000000000000010111100000100",
			2227 => "11111110001101110010001101000001",
			2228 => "00000010011011100010001101000001",
			2229 => "0000001001000000001011101000011100",
			2230 => "0000000000000000000011111100001100",
			2231 => "0000000010000000001110010000001000",
			2232 => "0000001110000000000110000100000100",
			2233 => "11111101110101110010001101000001",
			2234 => "00000000101100010010001101000001",
			2235 => "11111101101011110010001101000001",
			2236 => "0000000010000000001001100000001000",
			2237 => "0000001111000000001101000100000100",
			2238 => "00000000100011000010001101000001",
			2239 => "00000001111000000010001101000001",
			2240 => "0000001000000000000111000100000100",
			2241 => "11111111001011010010001101000001",
			2242 => "00000000011100110010001101000001",
			2243 => "0000000011000000001000000000010000",
			2244 => "0000000000000000000011111100001000",
			2245 => "0000001111000000001110101100000100",
			2246 => "00000001110110110010001101000001",
			2247 => "11111111111100000010001101000001",
			2248 => "0000000100000000001111100000000100",
			2249 => "11111110100100110010001101000001",
			2250 => "00000010011101110010001101000001",
			2251 => "0000001111000000001001100000001000",
			2252 => "0000001101000000000100000100000100",
			2253 => "00000000010100010010001101000001",
			2254 => "00000011000100010010001101000001",
			2255 => "11111110011000100010001101000001",
			2256 => "0000000101000000000011100011000000",
			2257 => "0000000100000000000011010101110100",
			2258 => "0000001110000000000100010100110100",
			2259 => "0000000011000000001001110000010100",
			2260 => "0000000000000000000100010100010000",
			2261 => "0000000110000000001101111100001000",
			2262 => "0000001011000000000100010100000100",
			2263 => "00000001011100110010010101010101",
			2264 => "00000000000000100010010101010101",
			2265 => "0000000000000000001010000000000100",
			2266 => "00000100111001000010010101010101",
			2267 => "00000001011110000010010101010101",
			2268 => "11111110001011100010010101010101",
			2269 => "0000001001000000000110101000010000",
			2270 => "0000000110000000001101111100001000",
			2271 => "0000000010000000001100100100000100",
			2272 => "00000011011100010010010101010101",
			2273 => "11111111111111000010010101010101",
			2274 => "0000001111000000000010001000000100",
			2275 => "00000110001010100010010101010101",
			2276 => "00000010001011100010010101010101",
			2277 => "0000000000000000000000111000001000",
			2278 => "0000001000000000000001110000000100",
			2279 => "11111111000100000010010101010101",
			2280 => "00000010101000100010010101010101",
			2281 => "0000000011000000001100110000000100",
			2282 => "11111111000011000010010101010101",
			2283 => "00000001110100110010010101010101",
			2284 => "0000000110000000000111101000100000",
			2285 => "0000001000000000000001010100010000",
			2286 => "0000001010000000000011101000001000",
			2287 => "0000001100000000000100010100000100",
			2288 => "11111111000011010010010101010101",
			2289 => "11111110010001100010010101010101",
			2290 => "0000000100000000001111101000000100",
			2291 => "00000011101101010010010101010101",
			2292 => "11111110110110010010010101010101",
			2293 => "0000001001000000000110101000001000",
			2294 => "0000000100000000001100001100000100",
			2295 => "00000101010111110010010101010101",
			2296 => "11111110011000000010010101010101",
			2297 => "0000001100000000000100010100000100",
			2298 => "11111110010100100010010101010101",
			2299 => "11111111100001100010010101010101",
			2300 => "0000000010000000000101110000010000",
			2301 => "0000001110000000000100000000001000",
			2302 => "0000001001000000000111100100000100",
			2303 => "00000011011111000010010101010101",
			2304 => "00000001101000110010010101010101",
			2305 => "0000000110000000001010011000000100",
			2306 => "00000100010001100010010101010101",
			2307 => "00000000100110000010010101010101",
			2308 => "0000001110000000001101100000001000",
			2309 => "0000001100000000000100010100000100",
			2310 => "00000010010101010010010101010101",
			2311 => "00000000110101010010010101010101",
			2312 => "0000001011000000000011011100000100",
			2313 => "00000011011101110010010101010101",
			2314 => "00000001100111100010010101010101",
			2315 => "0000000110000000001101111100010000",
			2316 => "0000000100000000000011110100000100",
			2317 => "00000010000001100010010101010101",
			2318 => "0000000001000000000000011000000100",
			2319 => "11111110010000010010010101010101",
			2320 => "0000001000000000000001110100000100",
			2321 => "11111110010101010010010101010101",
			2322 => "00000000111110000010010101010101",
			2323 => "0000001011000000001100001000100000",
			2324 => "0000000010000000000101001000010000",
			2325 => "0000001011000000000100010100001000",
			2326 => "0000000011000000001110111100000100",
			2327 => "00000000010111100010010101010101",
			2328 => "00000011111010110010010101010101",
			2329 => "0000000011000000000100010100000100",
			2330 => "11111110110101010010010101010101",
			2331 => "00000000110001100010010101010101",
			2332 => "0000001001000000000010001100001000",
			2333 => "0000000110000000000100110100000100",
			2334 => "00000101010000010010010101010101",
			2335 => "11111111000111110010010101010101",
			2336 => "0000001100000000000000101000000100",
			2337 => "00000001000101000010010101010101",
			2338 => "00000110111111000010010101010101",
			2339 => "0000001111000000001001010000010000",
			2340 => "0000000010000000001001011100001000",
			2341 => "0000000000000000000000101000000100",
			2342 => "00000001011001010010010101010101",
			2343 => "11111110110100000010010101010101",
			2344 => "0000001010000000000110011100000100",
			2345 => "11111110100111100010010101010101",
			2346 => "11111111100110000010010101010101",
			2347 => "0000001011000000000110000100001000",
			2348 => "0000000011000000000001101000000100",
			2349 => "11111111011011110010010101010101",
			2350 => "00000101000000010010010101010101",
			2351 => "11111110010111000010010101010101",
			2352 => "0000001100000000000110000100110100",
			2353 => "0000000011000000001000011000000100",
			2354 => "11111110010100110010010101010101",
			2355 => "0000000110000000001101011000010100",
			2356 => "0000000110000000000001111000000100",
			2357 => "11111110010111100010010101010101",
			2358 => "0000000101000000001000000000001000",
			2359 => "0000000110000000001101011000000100",
			2360 => "00000001110111010010010101010101",
			2361 => "11111111010001010010010101010101",
			2362 => "0000001011000000001010111000000100",
			2363 => "00000011100100010010010101010101",
			2364 => "00000110101011110010010101010101",
			2365 => "0000000110000000001001100100010000",
			2366 => "0000000010000000001100010000001000",
			2367 => "0000001001000000000001000100000100",
			2368 => "11111110010001010010010101010101",
			2369 => "11111111101111110010010101010101",
			2370 => "0000000010000000001000001100000100",
			2371 => "00000010010100100010010101010101",
			2372 => "11111110010111110010010101010101",
			2373 => "0000001100000000001100001000000100",
			2374 => "11111111100001100010010101010101",
			2375 => "0000000110000000001111000000000100",
			2376 => "11111110111000010010010101010101",
			2377 => "11111110001111110010010101010101",
			2378 => "0000001100000000000110000100010100",
			2379 => "0000001000000000001111001000010000",
			2380 => "0000001000000000000110001000001100",
			2381 => "0000001000000000000110011100000100",
			2382 => "11111110011010110010010101010101",
			2383 => "0000001000000000001100000100000100",
			2384 => "00000000100000000010010101010101",
			2385 => "11111110100101100010010101010101",
			2386 => "00000001101010100010010101010101",
			2387 => "11111110010101010010010101010101",
			2388 => "11111110010000100010010101010101",
			2389 => "0000001001000000000110101010000000",
			2390 => "0000000001000000001100110101110000",
			2391 => "0000000101000000001100101101000000",
			2392 => "0000001011000000000000101000100000",
			2393 => "0000001000000000000111000000010000",
			2394 => "0000000100000000001011100000001000",
			2395 => "0000000000000000001011000100000100",
			2396 => "00000000001000100010011101011001",
			2397 => "11111111011111100010011101011001",
			2398 => "0000001111000000000110100100000100",
			2399 => "11111110011100100010011101011001",
			2400 => "00000001010010010010011101011001",
			2401 => "0000001111000000000111010000001000",
			2402 => "0000000010000000001111010000000100",
			2403 => "11111111010111000010011101011001",
			2404 => "00000001100001010010011101011001",
			2405 => "0000000001000000000000011000000100",
			2406 => "00000000010000010010011101011001",
			2407 => "11111110000101010010011101011001",
			2408 => "0000001110000000001010000000010000",
			2409 => "0000001001000000001001111000001000",
			2410 => "0000001010000000001010110000000100",
			2411 => "11111111011011100010011101011001",
			2412 => "00000010011011010010011101011001",
			2413 => "0000000111000000000100010100000100",
			2414 => "00000000110001100010011101011001",
			2415 => "11111110111001010010011101011001",
			2416 => "0000000010000000001110010000001000",
			2417 => "0000000110000000000100110100000100",
			2418 => "00000001000101110010011101011001",
			2419 => "00000010010010000010011101011001",
			2420 => "0000000110000000000100110100000100",
			2421 => "11111110101011000010011101011001",
			2422 => "00000000101110110010011101011001",
			2423 => "0000000110000000000100110100010100",
			2424 => "0000001101000000001100101100000100",
			2425 => "00000000010100100010011101011001",
			2426 => "0000000111000000001100001000001000",
			2427 => "0000000100000000000101000000000100",
			2428 => "11111111001010110010011101011001",
			2429 => "11111101110011000010011101011001",
			2430 => "0000000100000000000101010100000100",
			2431 => "00000000001111010010011101011001",
			2432 => "11111101110110010010011101011001",
			2433 => "0000000010000000000101110000001100",
			2434 => "0000000010000000000001000000000100",
			2435 => "00000000000000000010011101011001",
			2436 => "0000001000000000001110001100000100",
			2437 => "00000010100010000010011101011001",
			2438 => "00000000000000000010011101011001",
			2439 => "0000000010000000000010000100001000",
			2440 => "0000000010000000001110010000000100",
			2441 => "00000000000110110010011101011001",
			2442 => "11111110010100000010011101011001",
			2443 => "0000001010000000000010101000000100",
			2444 => "00000011110000110010011101011001",
			2445 => "11111111101100010010011101011001",
			2446 => "0000000101000000000101101100000100",
			2447 => "11111111011010110010011101011001",
			2448 => "0000000010000000000101110000001000",
			2449 => "0000001011000000001100001000000100",
			2450 => "00000010101011000010011101011001",
			2451 => "00000000001110000010011101011001",
			2452 => "00000011101101100010011101011001",
			2453 => "0000000001000000001110100000001100",
			2454 => "0000001011000000001100001000001000",
			2455 => "0000000111000000000100010100000100",
			2456 => "11111111111100110010011101011001",
			2457 => "11111101111011000010011101011001",
			2458 => "11111100111011000010011101011001",
			2459 => "0000001110000000000100010100111100",
			2460 => "0000001011000000000000101000011100",
			2461 => "0000000100000000000101010100010000",
			2462 => "0000000100000000000010110000001000",
			2463 => "0000000111000000001011000100000100",
			2464 => "00000000000010100010011101011001",
			2465 => "11111101101011010010011101011001",
			2466 => "0000000001000000001110100000000100",
			2467 => "00000001011100000010011101011001",
			2468 => "00000011010011110010011101011001",
			2469 => "0000000100000000000011010100001000",
			2470 => "0000001111000000000010001000000100",
			2471 => "11111101110001100010011101011001",
			2472 => "11111111100110100010011101011001",
			2473 => "00000000110000100010011101011001",
			2474 => "0000001111000000000001011000010000",
			2475 => "0000000100000000000100001100001000",
			2476 => "0000001110000000000111111000000100",
			2477 => "11111110101011100010011101011001",
			2478 => "00000000001011110010011101011001",
			2479 => "0000001010000000000110011100000100",
			2480 => "00000100110101100010011101011001",
			2481 => "11111110110100010010011101011001",
			2482 => "0000000010000000001110000100001000",
			2483 => "0000001111000000000101100100000100",
			2484 => "11111110011010110010011101011001",
			2485 => "11111101000100010010011101011001",
			2486 => "0000000100000000001001001100000100",
			2487 => "00000000000000000010011101011001",
			2488 => "11111110010011100010011101011001",
			2489 => "0000000010000000001110000100011100",
			2490 => "0000000110000000000001111000010000",
			2491 => "0000001110000000000100000000001000",
			2492 => "0000000100000000000010010100000100",
			2493 => "00000000010111000010011101011001",
			2494 => "11111101110001110010011101011001",
			2495 => "0000001010000000000011101000000100",
			2496 => "11111110111001100010011101011001",
			2497 => "00000001000010000010011101011001",
			2498 => "0000000100000000000010111000001000",
			2499 => "0000000000000000000011010000000100",
			2500 => "00000000111111110010011101011001",
			2501 => "11111110100011100010011101011001",
			2502 => "00000010110000100010011101011001",
			2503 => "0000001000000000000001110100010000",
			2504 => "0000001001000000000110101000001000",
			2505 => "0000001111000000000101110100000100",
			2506 => "00000001000100100010011101011001",
			2507 => "11111111111101100010011101011001",
			2508 => "0000001110000000001000111000000100",
			2509 => "11111111100000010010011101011001",
			2510 => "11111111111110100010011101011001",
			2511 => "0000000000000000000111111000001000",
			2512 => "0000000110000000001011001100000100",
			2513 => "00000011000100000010011101011001",
			2514 => "00000000011000100010011101011001",
			2515 => "0000000001000000001001111000000100",
			2516 => "00000000010110000010011101011001",
			2517 => "11111110101001000010011101011001",
			2518 => "0000001100000000000100001010101100",
			2519 => "0000000011000000001011000100111000",
			2520 => "0000001111000000000001011000110100",
			2521 => "0000000111000000000111111000011000",
			2522 => "0000001000000000001001101000001000",
			2523 => "0000000011000000001010000000000100",
			2524 => "00000001010001110010100010110101",
			2525 => "00000100010110110010100010110101",
			2526 => "0000000111000000000111111000001000",
			2527 => "0000001100000000000111111000000100",
			2528 => "11111111010011110010100010110101",
			2529 => "00000001011110100010100010110101",
			2530 => "0000001100000000000111111000000100",
			2531 => "00000010111010000010100010110101",
			2532 => "11111110101001010010100010110101",
			2533 => "0000000011000000000111111000010000",
			2534 => "0000001010000000000110011100001000",
			2535 => "0000000110000000000001111000000100",
			2536 => "00000000000111110010100010110101",
			2537 => "11111110100110100010100010110101",
			2538 => "0000001010000000000001110000000100",
			2539 => "00000000101111000010100010110101",
			2540 => "11111110110001010010100010110101",
			2541 => "0000001011000000001110111100000100",
			2542 => "00000010110010110010100010110101",
			2543 => "0000000100000000000000010100000100",
			2544 => "11111111010011110010100010110101",
			2545 => "00000000011101000010100010110101",
			2546 => "11111110000011000010100010110101",
			2547 => "0000001111000000000010001000111100",
			2548 => "0000000101000000000011011100011100",
			2549 => "0000001010000000001010110000010000",
			2550 => "0000001101000000001100110000001000",
			2551 => "0000001011000000001011000100000100",
			2552 => "00000000110100010010100010110101",
			2553 => "11111110101011000010100010110101",
			2554 => "0000000011000000000100000000000100",
			2555 => "00000001010100000010100010110101",
			2556 => "00000100011011010010100010110101",
			2557 => "0000000101000000000011011100001000",
			2558 => "0000001100000000000111111000000100",
			2559 => "00000011000000000010100010110101",
			2560 => "00000000001101110010100010110101",
			2561 => "00000100100101000010100010110101",
			2562 => "0000000011000000000100000000010000",
			2563 => "0000001111000000000110100100001000",
			2564 => "0000001101000000001100101100000100",
			2565 => "00000100111000100010100010110101",
			2566 => "11111111100001000010100010110101",
			2567 => "0000000001000000001110100000000100",
			2568 => "11111111011111000010100010110101",
			2569 => "00000010001010110010100010110101",
			2570 => "0000001101000000001100101000001000",
			2571 => "0000000011000000001100110000000100",
			2572 => "00000000010011000010100010110101",
			2573 => "00000000111111110010100010110101",
			2574 => "0000000011000000001110001100000100",
			2575 => "11111110110110010010100010110101",
			2576 => "00000000000000010010100010110101",
			2577 => "0000000011000000000101101100011000",
			2578 => "0000000011000000000101101100010000",
			2579 => "0000000011000000001100110000001000",
			2580 => "0000001101000000000110000100000100",
			2581 => "11111111110110100010100010110101",
			2582 => "11111110100010100010100010110101",
			2583 => "0000001100000000000100010100000100",
			2584 => "00000010010001110010100010110101",
			2585 => "11111111110100000010100010110101",
			2586 => "0000001111000000000101110100000100",
			2587 => "11111110101111110010100010110101",
			2588 => "11111101100100110010100010110101",
			2589 => "0000001000000000000010101000010000",
			2590 => "0000000100000000000000010100001000",
			2591 => "0000001000000000000111000100000100",
			2592 => "00000000000010110010100010110101",
			2593 => "00000000101010010010100010110101",
			2594 => "0000001010000000001010110000000100",
			2595 => "11111111000010100010100010110101",
			2596 => "00000000000111110010100010110101",
			2597 => "0000000010000000000010000000001000",
			2598 => "0000000110000000001010011000000100",
			2599 => "00000100100001010010100010110101",
			2600 => "00000000011100010010100010110101",
			2601 => "0000000100000000000010100100000100",
			2602 => "00000001001111110010100010110101",
			2603 => "11111111110001100010100010110101",
			2604 => "11111110011100010010100010110101",
			2605 => "0000001111000000000000110111100100",
			2606 => "0000001110000000001010000001101100",
			2607 => "0000001011000000000100010100110100",
			2608 => "0000000001000000001110100000011100",
			2609 => "0000001001000000001001111000010000",
			2610 => "0000001100000000000111111000001000",
			2611 => "0000000111000000000111111000000100",
			2612 => "00000000001001010010101110100011",
			2613 => "11111111010001000010101110100011",
			2614 => "0000000111000000001010000000000100",
			2615 => "11111101111101010010101110100011",
			2616 => "00000000101010010010101110100011",
			2617 => "0000001011000000000100010100001000",
			2618 => "0000001100000000000111111000000100",
			2619 => "11111111101001110010101110100011",
			2620 => "11111110001001110010101110100011",
			2621 => "00000001000000000010101110100011",
			2622 => "0000001100000000000111111000001100",
			2623 => "0000001001000000001001111000000100",
			2624 => "00000001010001100010101110100011",
			2625 => "0000000011000000001100001000000100",
			2626 => "11111110001000010010101110100011",
			2627 => "00000000000101000010101110100011",
			2628 => "0000000111000000001011000100001000",
			2629 => "0000001101000000000101101100000100",
			2630 => "00000010110001000010101110100011",
			2631 => "00000000111010010010101110100011",
			2632 => "11111111010110010010101110100011",
			2633 => "0000000110000000001100011000011000",
			2634 => "0000000010000000000010000000010000",
			2635 => "0000001001000000000010001100001000",
			2636 => "0000000001000000000110000000000100",
			2637 => "11111111100000000010101110100011",
			2638 => "00000011010011010010101110100011",
			2639 => "0000001110000000000000111000000100",
			2640 => "11111110110111100010101110100011",
			2641 => "11111111101111100010101110100011",
			2642 => "0000000010000000000010000000000100",
			2643 => "00000111101100100010101110100011",
			2644 => "00000000000000000010101110100011",
			2645 => "0000001111000000000100000100010000",
			2646 => "0000001111000000001000011000001000",
			2647 => "0000000010000000001111010000000100",
			2648 => "11111110010100110010101110100011",
			2649 => "00000001100011110010101110100011",
			2650 => "0000000111000000001100001000000100",
			2651 => "00000010001110100010101110100011",
			2652 => "11111110100100010010101110100011",
			2653 => "0000001101000000001110001100001000",
			2654 => "0000000101000000001101100000000100",
			2655 => "00000000111000100010101110100011",
			2656 => "11111110011011110010101110100011",
			2657 => "0000001001000000000110101000000100",
			2658 => "00000010011000010010101110100011",
			2659 => "11111110110111010010101110100011",
			2660 => "0000001101000000001100101100111100",
			2661 => "0000001011000000000000101000100000",
			2662 => "0000000011000000000101101100010000",
			2663 => "0000001111000000000101110100001000",
			2664 => "0000001100000000000100010100000100",
			2665 => "00000000001101000010101110100011",
			2666 => "00000010000100110010101110100011",
			2667 => "0000000111000000000100010100000100",
			2668 => "00000000011001110010101110100011",
			2669 => "11111110101110110010101110100011",
			2670 => "0000000100000000001010110100001000",
			2671 => "0000001111000000001010010100000100",
			2672 => "00000000110010010010101110100011",
			2673 => "11111110010001110010101110100011",
			2674 => "0000000100000000000000010100000100",
			2675 => "00000011000001000010101110100011",
			2676 => "00000001011001010010101110100011",
			2677 => "0000001010000000000001010000010000",
			2678 => "0000001010000000000110011000001000",
			2679 => "0000000111000000000100010100000100",
			2680 => "00000010011110110010101110100011",
			2681 => "00000000100001110010101110100011",
			2682 => "0000000010000000000100101000000100",
			2683 => "11111111000001000010101110100011",
			2684 => "00000001000101100010101110100011",
			2685 => "0000001111000000001011011100000100",
			2686 => "00000011000011100010101110100011",
			2687 => "0000001110000000000100010100000100",
			2688 => "11111111100010100010101110100011",
			2689 => "00000001011111000010101110100011",
			2690 => "0000001110000000001101100000100000",
			2691 => "0000001001000000000111100100010000",
			2692 => "0000000001000000001100110100001000",
			2693 => "0000001001000000000110101000000100",
			2694 => "00000000000111010010101110100011",
			2695 => "11111111000101010010101110100011",
			2696 => "0000001100000000000100000000000100",
			2697 => "00000000001100010010101110100011",
			2698 => "00000010100000100010101110100011",
			2699 => "0000000100000000000011001100001000",
			2700 => "0000000011000000001110001100000100",
			2701 => "11111110101101110010101110100011",
			2702 => "00000000101111010010101110100011",
			2703 => "0000000110000000001010011000000100",
			2704 => "11111110011110110010101110100011",
			2705 => "11111111111010110010101110100011",
			2706 => "0000001001000000001011101000010000",
			2707 => "0000001100000000000100010100001000",
			2708 => "0000001100000000000100010100000100",
			2709 => "00000000011110000010101110100011",
			2710 => "11111110101001110010101110100011",
			2711 => "0000001011000000000100000000000100",
			2712 => "00000001100000100010101110100011",
			2713 => "00000000100110110010101110100011",
			2714 => "0000001010000000001010110000001000",
			2715 => "0000000001000000001001111000000100",
			2716 => "11111111101100100010101110100011",
			2717 => "00000000110000110010101110100011",
			2718 => "11111101111100110010101110100011",
			2719 => "0000000111000000000100000001011100",
			2720 => "0000001010000000001100011100101100",
			2721 => "0000000100000000001010110100011000",
			2722 => "0000001100000000000100000000001100",
			2723 => "0000000110000000001101111100000100",
			2724 => "11111101111001100010101110100011",
			2725 => "0000000010000000000010000000000100",
			2726 => "00000000010110010010101110100011",
			2727 => "11111111010110010010101110100011",
			2728 => "0000001101000000001010111000001000",
			2729 => "0000001010000000000001010000000100",
			2730 => "11111101001110010010101110100011",
			2731 => "11111111000110010010101110100011",
			2732 => "00000000111001000010101110100011",
			2733 => "0000001101000000000101101100001000",
			2734 => "0000000111000000000111111000000100",
			2735 => "11111110110000000010101110100011",
			2736 => "00000010011001110010101110100011",
			2737 => "0000000010000000000011001000000100",
			2738 => "00000000110101100010101110100011",
			2739 => "0000001100000000000100000000000100",
			2740 => "11111110110111000010101110100011",
			2741 => "00000000100010100010101110100011",
			2742 => "0000001011000000001001110000100000",
			2743 => "0000000100000000000011010100010000",
			2744 => "0000000101000000000000001100001000",
			2745 => "0000000010000000000110010000000100",
			2746 => "00000001011100010010101110100011",
			2747 => "11111111010110010010101110100011",
			2748 => "0000000110000000001010011000000100",
			2749 => "00000011000000100010101110100011",
			2750 => "00000001100100110010101110100011",
			2751 => "0000000111000000001100001000001000",
			2752 => "0000001110000000001000111000000100",
			2753 => "11111110010101010010101110100011",
			2754 => "00000000101011110010101110100011",
			2755 => "0000001100000000000100010100000100",
			2756 => "00000000000000000010101110100011",
			2757 => "11111110010001110010101110100011",
			2758 => "0000001100000000000000101000000100",
			2759 => "00000001100000100010101110100011",
			2760 => "0000001110000000001100101100000100",
			2761 => "11111111010001010010101110100011",
			2762 => "0000000101000000001010111100000100",
			2763 => "11111101011001110010101110100011",
			2764 => "11111110101101100010101110100011",
			2765 => "0000000111000000001000111000011100",
			2766 => "0000001111000000000000110100000100",
			2767 => "11111110101001000010101110100011",
			2768 => "0000000001000000000010001100001100",
			2769 => "0000001011000000001000111000000100",
			2770 => "00000000010010000010101110100011",
			2771 => "0000000001000000000010001100000100",
			2772 => "00000001101000000010101110100011",
			2773 => "00000010110100100010101110100011",
			2774 => "0000000110000000001101011000001000",
			2775 => "0000000100000000000011110000000100",
			2776 => "00000001000010000010101110100011",
			2777 => "11111111100011100010101110100011",
			2778 => "00000001110101110010101110100011",
			2779 => "0000000011000000000100001000000100",
			2780 => "00000010100000110010101110100011",
			2781 => "0000001001000000000111100100001000",
			2782 => "0000001111000000001110101100000100",
			2783 => "11111110101011010010101110100011",
			2784 => "11111100111001100010101110100011",
			2785 => "0000001100000000000000101000001000",
			2786 => "0000000110000000001010011000000100",
			2787 => "00000000001010110010101110100011",
			2788 => "11111110110110010010101110100011",
			2789 => "0000000010000000000101110000000100",
			2790 => "11111110001111010010101110100011",
			2791 => "00000000000110000010101110100011",
			2792 => "0000000101000000001000000001110100",
			2793 => "0000000111000000001101100001011000",
			2794 => "0000000111000000001101100000111100",
			2795 => "0000000111000000000000101000100000",
			2796 => "0000000111000000000100010100010000",
			2797 => "0000000111000000000100010100001000",
			2798 => "0000000001000000001100110100000100",
			2799 => "00000000000101000010110100010101",
			2800 => "00000001110110100010110100010101",
			2801 => "0000001011000000000100010100000100",
			2802 => "11111110101010100010110100010101",
			2803 => "11111111101111100010110100010101",
			2804 => "0000000101000000000011011100001000",
			2805 => "0000000111000000001011000100000100",
			2806 => "00000010001100110010110100010101",
			2807 => "00000000110011000010110100010101",
			2808 => "0000000010000000000010000100000100",
			2809 => "00000000001111000010110100010101",
			2810 => "00000010111110010010110100010101",
			2811 => "0000000111000000000000101000001100",
			2812 => "0000000110000000000111101000000100",
			2813 => "00000001100011000010110100010101",
			2814 => "0000000101000000001110001100000100",
			2815 => "11111110100111110010110100010101",
			2816 => "11111111111100110010110100010101",
			2817 => "0000001010000000000111110100001000",
			2818 => "0000000010000000001001010000000100",
			2819 => "11111111100001100010110100010101",
			2820 => "11111101110010110010110100010101",
			2821 => "0000000111000000001100001000000100",
			2822 => "00000000010001000010110100010101",
			2823 => "11111111111110010010110100010101",
			2824 => "0000001110000000001010111000001100",
			2825 => "0000000111000000001101100000001000",
			2826 => "0000001000000000000110001000000100",
			2827 => "00000001011011010010110100010101",
			2828 => "00000100010001100010110100010101",
			2829 => "11111111000101010010110100010101",
			2830 => "0000000110000000001101011000000100",
			2831 => "11111110110100110010110100010101",
			2832 => "0000001100000000001000111100001000",
			2833 => "0000001011000000001100101100000100",
			2834 => "11111110101010110010110100010101",
			2835 => "00000000100011100010110100010101",
			2836 => "00000010011000100010110100010101",
			2837 => "0000001010000000000110011000010000",
			2838 => "0000001100000000001000111000000100",
			2839 => "11111110001010100010110100010101",
			2840 => "0000001100000000001001110000001000",
			2841 => "0000001010000000001100011000000100",
			2842 => "00000000000000000010110100010101",
			2843 => "00000010110001110010110100010101",
			2844 => "11111110111111110010110100010101",
			2845 => "0000001111000000001001010000000100",
			2846 => "11111110001110000010110100010101",
			2847 => "0000000011000000000000011100000100",
			2848 => "00000000100110110010110100010101",
			2849 => "11111110011100110010110100010101",
			2850 => "0000001110000000001001010100101100",
			2851 => "0000001010000000001100011100101000",
			2852 => "0000001000000000001111001000011000",
			2853 => "0000000101000000001000011000001100",
			2854 => "0000000010000000001100010000001000",
			2855 => "0000001010000000000001010000000100",
			2856 => "00000001001110000010110100010101",
			2857 => "11111110100001110010110100010101",
			2858 => "11111110010101110010110100010101",
			2859 => "0000000101000000001010001100001000",
			2860 => "0000000010000000001100100100000100",
			2861 => "00000000000000000010110100010101",
			2862 => "00000010100001100010110100010101",
			2863 => "00000000000000000010110100010101",
			2864 => "0000000010000000000111011000000100",
			2865 => "00000001001111010010110100010101",
			2866 => "0000001111000000000010000000001000",
			2867 => "0000000111000000001110001100000100",
			2868 => "00000011110101110010110100010101",
			2869 => "00000000000000000010110100010101",
			2870 => "00000000000000000010110100010101",
			2871 => "11111110100111010010110100010101",
			2872 => "0000000001000000001101101000001000",
			2873 => "0000000010000000000110010000000100",
			2874 => "00000000100001000010110100010101",
			2875 => "11111110010101100010110100010101",
			2876 => "0000001100000000001010111100010000",
			2877 => "0000000110000000001111000000001100",
			2878 => "0000000010000000000010000100000100",
			2879 => "11111111011011010010110100010101",
			2880 => "0000001100000000001100110000000100",
			2881 => "00000010000010110010110100010101",
			2882 => "00000000011011010010110100010101",
			2883 => "11111110111010100010110100010101",
			2884 => "11111110100111010010110100010101",
			2885 => "0000000111000000001101100001111000",
			2886 => "0000000001000000001100100000001000",
			2887 => "0000000110000000001101111100000100",
			2888 => "11111110010011000010111001111001",
			2889 => "00000001001010110010111001111001",
			2890 => "0000001000000000000111000101000000",
			2891 => "0000000110000000001101111100100000",
			2892 => "0000000010000000001010001000010000",
			2893 => "0000000011000000000100000000001000",
			2894 => "0000001011000000000111111000000100",
			2895 => "00000001100100010010111001111001",
			2896 => "11111111111100110010111001111001",
			2897 => "0000001010000000000111110100000100",
			2898 => "00000000001000100010111001111001",
			2899 => "00000001110011100010111001111001",
			2900 => "0000001000000000000110001000001000",
			2901 => "0000000011000000001110001100000100",
			2902 => "11111110000111000010111001111001",
			2903 => "11111111001010000010111001111001",
			2904 => "0000000111000000000100010100000100",
			2905 => "00000010001011100010111001111001",
			2906 => "11111110101010100010111001111001",
			2907 => "0000000010000000001001100000010000",
			2908 => "0000001000000000001111001000001000",
			2909 => "0000001100000000000100000000000100",
			2910 => "00000010100010100010111001111001",
			2911 => "00000001011100110010111001111001",
			2912 => "0000001010000000000001010000000100",
			2913 => "11111111111001010010111001111001",
			2914 => "00000001110110000010111001111001",
			2915 => "0000001110000000000001111100001000",
			2916 => "0000000010000000001110110100000100",
			2917 => "11111111001010100010111001111001",
			2918 => "11111101110111010010111001111001",
			2919 => "0000000101000000001010111000000100",
			2920 => "00000001101001010010111001111001",
			2921 => "11111111000100100010111001111001",
			2922 => "0000000111000000000111111000010100",
			2923 => "0000000010000000001101000100001000",
			2924 => "0000001011000000001110111100000100",
			2925 => "00000001011001010010111001111001",
			2926 => "11111111011010010010111001111001",
			2927 => "0000000001000000001110100000001000",
			2928 => "0000001000000000000010101000000100",
			2929 => "00000001110001010010111001111001",
			2930 => "00000100110100110010111001111001",
			2931 => "00000000100010110010111001111001",
			2932 => "0000001000000000000111000000010000",
			2933 => "0000000011000000000100010100001000",
			2934 => "0000000110000000001100011000000100",
			2935 => "11111110110011010010111001111001",
			2936 => "00000001100010110010111001111001",
			2937 => "0000000111000000001100001000000100",
			2938 => "00000001010101100010111001111001",
			2939 => "00000000010110010010111001111001",
			2940 => "0000000110000000000100110100000100",
			2941 => "00000010110011100010111001111001",
			2942 => "0000000001000000001110100000000100",
			2943 => "11111111101111100010111001111001",
			2944 => "11111110101011100010111001111001",
			2945 => "0000001100000000001100110000101100",
			2946 => "0000000011000000000001101000010000",
			2947 => "0000000011000000001001110100000100",
			2948 => "11111110001111000010111001111001",
			2949 => "0000000010000000000011001000001000",
			2950 => "0000000101000000001001110100000100",
			2951 => "00000001000111110010111001111001",
			2952 => "11111110100111100010111001111001",
			2953 => "11111110001111010010111001111001",
			2954 => "0000000110000000001011001100010000",
			2955 => "0000000110000000000001111000000100",
			2956 => "11111110011000000010111001111001",
			2957 => "0000001111000000001110101000000100",
			2958 => "00000100011001010010111001111001",
			2959 => "0000000010000000001100010000000100",
			2960 => "11111111101110110010111001111001",
			2961 => "00000010000111000010111001111001",
			2962 => "0000001101000000000111010000000100",
			2963 => "11111110010000010010111001111001",
			2964 => "0000000010000000000000010000000100",
			2965 => "00000101101000100010111001111001",
			2966 => "11111110010111100010111001111001",
			2967 => "0000000111000000001101111000001100",
			2968 => "0000000111000000001110001100000100",
			2969 => "11111110010111010010111001111001",
			2970 => "0000001100000000000110000100000100",
			2971 => "00000001100101100010111001111001",
			2972 => "11111110110110100010111001111001",
			2973 => "11111110010011010010111001111001",
			2974 => "0000001100000000000011011101101100",
			2975 => "0000000100000000000011111001101000",
			2976 => "0000000111000000001001110001000000",
			2977 => "0000001110000000001101100000100000",
			2978 => "0000001001000000001101101000010000",
			2979 => "0000000010000000001010001000001000",
			2980 => "0000001110000000000100010100000100",
			2981 => "00000000011010000010111110100101",
			2982 => "00000000111010110010111110100101",
			2983 => "0000001010000000000001010000000100",
			2984 => "11111111011011110010111110100101",
			2985 => "00000000011011010010111110100101",
			2986 => "0000000100000000000011001100001000",
			2987 => "0000000011000000001110001100000100",
			2988 => "11111110101001100010111110100101",
			2989 => "00000000101010110010111110100101",
			2990 => "0000001000000000000110001000000100",
			2991 => "11111101001010100010111110100101",
			2992 => "11111111010100100010111110100101",
			2993 => "0000001001000000001101101000010000",
			2994 => "0000000100000000001111100000001000",
			2995 => "0000001010000000000110011100000100",
			2996 => "00000001001100000010111110100101",
			2997 => "00000100000010100010111110100101",
			2998 => "0000001110000000001110001100000100",
			2999 => "11111110101010000010111110100101",
			3000 => "00000000110110010010111110100101",
			3001 => "0000001110000000000110000100001000",
			3002 => "0000000010000000000111111100000100",
			3003 => "00000000010000010010111110100101",
			3004 => "11111110100100010010111110100101",
			3005 => "0000000100000000001101001000000100",
			3006 => "00000001000010110010111110100101",
			3007 => "00000000001111000010111110100101",
			3008 => "0000000110000000001111000000100000",
			3009 => "0000000010000000000111011000010000",
			3010 => "0000001010000000001100011100001000",
			3011 => "0000000110000000000001111000000100",
			3012 => "11111110001110100010111110100101",
			3013 => "00000000001010100010111110100101",
			3014 => "0000001001000000001011101000000100",
			3015 => "00000000011011100010111110100101",
			3016 => "11111110010110110010111110100101",
			3017 => "0000000000000000001010000000001000",
			3018 => "0000000111000000001101100000000100",
			3019 => "11111110000100010010111110100101",
			3020 => "00000001100110010010111110100101",
			3021 => "0000001011000000000110000100000100",
			3022 => "00000100010001110010111110100101",
			3023 => "00000000110111110010111110100101",
			3024 => "0000001011000000000001111100000100",
			3025 => "11111110010110110010111110100101",
			3026 => "00000000100100110010111110100101",
			3027 => "11111110011000000010111110100101",
			3028 => "0000001100000000000110000100011000",
			3029 => "0000001011000000001000000000010100",
			3030 => "0000001001000000001101011100000100",
			3031 => "11111110001110000010111110100101",
			3032 => "0000001001000000001101011100000100",
			3033 => "00000010110100010010111110100101",
			3034 => "0000001011000000001010111100001000",
			3035 => "0000001101000000000111010000000100",
			3036 => "11111110111100010010111110100101",
			3037 => "00000010001100100010111110100101",
			3038 => "11111110010110010010111110100101",
			3039 => "00000001110100110010111110100101",
			3040 => "0000001100000000001010111100010000",
			3041 => "0000001000000000000110011100001100",
			3042 => "0000001000000000001100011100000100",
			3043 => "11111110011100000010111110100101",
			3044 => "0000001100000000000100001000000100",
			3045 => "00000000110000100010111110100101",
			3046 => "00000011000011110010111110100101",
			3047 => "11111110011000010010111110100101",
			3048 => "11111110010111110010111110100101",
			3049 => "0000001100000000000011011101111000",
			3050 => "0000000100000000000011111001110100",
			3051 => "0000001001000000001111001100111100",
			3052 => "0000000110000000001010011000100000",
			3053 => "0000001111000000000010110100010000",
			3054 => "0000001110000000000110000100001000",
			3055 => "0000001001000000001101101000000100",
			3056 => "00000000011111000011000100000001",
			3057 => "11111111010000110011000100000001",
			3058 => "0000001011000000000011011100000100",
			3059 => "00000001010101000011000100000001",
			3060 => "00000000000011010011000100000001",
			3061 => "0000000110000000001100011000001000",
			3062 => "0000001111000000001110101000000100",
			3063 => "11111111010010010011000100000001",
			3064 => "11111101101111110011000100000001",
			3065 => "0000000100000000001101001000000100",
			3066 => "00000001011011110011000100000001",
			3067 => "11111111111110000011000100000001",
			3068 => "0000000000000000001011000100010000",
			3069 => "0000001001000000001101101000001000",
			3070 => "0000000100000000001111100000000100",
			3071 => "00000010111100110011000100000001",
			3072 => "11111111010100110011000100000001",
			3073 => "0000000011000000000100011000000100",
			3074 => "00000000100010000011000100000001",
			3075 => "00000001110001100011000100000001",
			3076 => "0000000110000000001010011000000100",
			3077 => "00000011010011100011000100000001",
			3078 => "0000001110000000000000001100000100",
			3079 => "11111110110100110011000100000001",
			3080 => "00000001010000000011000100000001",
			3081 => "0000001110000000000111001000011100",
			3082 => "0000000000000000000011010000010000",
			3083 => "0000001111000000001010010100001000",
			3084 => "0000001011000000000110000100000100",
			3085 => "11111100111100110011000100000001",
			3086 => "11111110010110100011000100000001",
			3087 => "0000001011000000001100110000000100",
			3088 => "00000000000000000011000100000001",
			3089 => "00000010110001000011000100000001",
			3090 => "0000000011000000001001110100001000",
			3091 => "0000000111000000001101100000000100",
			3092 => "11111101010110110011000100000001",
			3093 => "11111110111110010011000100000001",
			3094 => "11111111111010000011000100000001",
			3095 => "0000001100000000000000101000001100",
			3096 => "0000000100000000001000000100000100",
			3097 => "00000000101010110011000100000001",
			3098 => "0000001011000000001101100000000100",
			3099 => "11111100100011110011000100000001",
			3100 => "11111110111000110011000100000001",
			3101 => "0000000111000000001000111000001000",
			3102 => "0000001001000000001001011000000100",
			3103 => "00000010010100010011000100000001",
			3104 => "11111111001000010011000100000001",
			3105 => "0000000100000000001000100000000100",
			3106 => "00000001110101000011000100000001",
			3107 => "00000000000001000011000100000001",
			3108 => "11111110011000110011000100000001",
			3109 => "0000001100000000000110000100100100",
			3110 => "0000001001000000001011111100010000",
			3111 => "0000000111000000000101101100000100",
			3112 => "11111110001101110011000100000001",
			3113 => "0000000111000000000101101100000100",
			3114 => "00000001001011010011000100000001",
			3115 => "0000001011000000001100101100000100",
			3116 => "00000000001001010011000100000001",
			3117 => "11111110010111110011000100000001",
			3118 => "0000000000000000000010101000001000",
			3119 => "0000001111000000001100100100000100",
			3120 => "11111110111100000011000100000001",
			3121 => "00000010010111110011000100000001",
			3122 => "0000001001000000000111101000001000",
			3123 => "0000001001000000001110010100000100",
			3124 => "11111111010000100011000100000001",
			3125 => "00000010001101110011000100000001",
			3126 => "11111110010111010011000100000001",
			3127 => "0000001100000000001010111100010000",
			3128 => "0000001000000000000110011100001100",
			3129 => "0000001000000000001100011100000100",
			3130 => "11111110011110100011000100000001",
			3131 => "0000001100000000000100001000000100",
			3132 => "00000000100111100011000100000001",
			3133 => "00000010010101000011000100000001",
			3134 => "11111110011001000011000100000001",
			3135 => "11111110011000010011000100000001",
			3136 => "0000001100000000001000111001111000",
			3137 => "0000001001000000000110000000000100",
			3138 => "11111110010100000011001001100101",
			3139 => "0000001110000000001100001000111000",
			3140 => "0000000111000000001100001000011100",
			3141 => "0000001110000000000011010000001100",
			3142 => "0000001000000000000101000100000100",
			3143 => "00000100011010010011001001100101",
			3144 => "0000001001000000001100110100000100",
			3145 => "00000001011101100011001001100101",
			3146 => "00000000000100010011001001100101",
			3147 => "0000001111000000000010001000001000",
			3148 => "0000001000000000000101000100000100",
			3149 => "11111110001110110011001001100101",
			3150 => "00000001100001110011001001100101",
			3151 => "0000001101000000001100101100000100",
			3152 => "00000000110110110011001001100101",
			3153 => "11111111011010110011001001100101",
			3154 => "0000000011000000001101100000010000",
			3155 => "0000001001000000000110101000001000",
			3156 => "0000000011000000001100001000000100",
			3157 => "11111110001110110011001001100101",
			3158 => "00000000001110010011001001100101",
			3159 => "0000001010000000001000010100000100",
			3160 => "11111111011100100011001001100101",
			3161 => "11111110001000010011001001100101",
			3162 => "0000001001000000000110101000000100",
			3163 => "00000011011011000011001001100101",
			3164 => "0000001111000000000000011100000100",
			3165 => "00000010010000000011001001100101",
			3166 => "11111111101110110011001001100101",
			3167 => "0000000010000000001010001000100000",
			3168 => "0000000110000000000001111000010000",
			3169 => "0000001011000000000100000000001000",
			3170 => "0000001101000000001110001100000100",
			3171 => "00000000000000110011001001100101",
			3172 => "00000010111111110011001001100101",
			3173 => "0000000110000000000111101000000100",
			3174 => "11111110010010110011001001100101",
			3175 => "11111111101001110011001001100101",
			3176 => "0000001001000000001101101000001000",
			3177 => "0000001111000000000010001000000100",
			3178 => "00000011001110000011001001100101",
			3179 => "00000010010000110011001001100101",
			3180 => "0000001000000000000111000100000100",
			3181 => "00000001111111010011001001100101",
			3182 => "11111110000111110011001001100101",
			3183 => "0000000011000000000001011000010000",
			3184 => "0000001110000000000110000100001000",
			3185 => "0000001011000000001100001000000100",
			3186 => "00000001100011000011001001100101",
			3187 => "00000000001010000011001001100101",
			3188 => "0000000111000000000100000000000100",
			3189 => "00000010010010010011001001100101",
			3190 => "00000001001011000011001001100101",
			3191 => "0000000101000000000001101000001000",
			3192 => "0000001101000000001000000000000100",
			3193 => "00000000010010000011001001100101",
			3194 => "11111110100101110011001001100101",
			3195 => "00000001010110110011001001100101",
			3196 => "0000001100000000001100110000101100",
			3197 => "0000001111000000001101000100010000",
			3198 => "0000000111000000001001110000000100",
			3199 => "00000000000000000011001001100101",
			3200 => "0000001111000000000010110100000100",
			3201 => "11111110010010100011001001100101",
			3202 => "0000001111000000000110100000000100",
			3203 => "00000000000000000011001001100101",
			3204 => "11111110010000000011001001100101",
			3205 => "0000000010000000001000001100010100",
			3206 => "0000001101000000000100000100001100",
			3207 => "0000000001000000000111100100001000",
			3208 => "0000001101000000000001101000000100",
			3209 => "00000000001000010011001001100101",
			3210 => "00000010011001100011001001100101",
			3211 => "11111110001110000011001001100101",
			3212 => "0000000011000000000110100000000100",
			3213 => "00000011101001000011001001100101",
			3214 => "00000000111001100011001001100101",
			3215 => "0000001010000000000001010000000100",
			3216 => "00000000110100100011001001100101",
			3217 => "11111110010110100011001001100101",
			3218 => "0000000111000000001101111000001100",
			3219 => "0000000111000000001110001100000100",
			3220 => "11111110011000010011001001100101",
			3221 => "0000001100000000000110000100000100",
			3222 => "00000001010111100011001001100101",
			3223 => "11111110111011110011001001100101",
			3224 => "11111110010100100011001001100101",
			3225 => "0000001100000000000110000101111000",
			3226 => "0000000100000000000011111001110100",
			3227 => "0000000010000000001110000100111100",
			3228 => "0000000110000000000111101000011100",
			3229 => "0000000101000000000101101100010000",
			3230 => "0000000011000000001000111100001000",
			3231 => "0000001000000000000001110000000100",
			3232 => "00000001101110010011001110001001",
			3233 => "11111111010101110011001110001001",
			3234 => "0000000111000000000100010100000100",
			3235 => "00000000001000000011001110001001",
			3236 => "00000011111110110011001110001001",
			3237 => "0000001111000000001010001100000100",
			3238 => "11111110010000100011001110001001",
			3239 => "0000001001000000001011101000000100",
			3240 => "11111111011110100011001110001001",
			3241 => "00000010111110100011001110001001",
			3242 => "0000001101000000001100110000010000",
			3243 => "0000000100000000001001001100001000",
			3244 => "0000001000000000001011010100000100",
			3245 => "00000000010111000011001110001001",
			3246 => "11111110111100010011001110001001",
			3247 => "0000001010000000000001010000000100",
			3248 => "00000011001001110011001110001001",
			3249 => "00000000001101110011001110001001",
			3250 => "0000001010000000001001000100001000",
			3251 => "0000000011000000001101100000000100",
			3252 => "11111111111010110011001110001001",
			3253 => "00000000111011110011001110001001",
			3254 => "0000000110000000001101111100000100",
			3255 => "00000010000110000011001110001001",
			3256 => "00000000110100110011001110001001",
			3257 => "0000001010000000001100011100011100",
			3258 => "0000000010000000001110000100001100",
			3259 => "0000000100000000001110100100000100",
			3260 => "11111101010011110011001110001001",
			3261 => "0000000100000000000011110000000100",
			3262 => "00000001110000100011001110001001",
			3263 => "11111110100011010011001110001001",
			3264 => "0000000100000000001110111000001000",
			3265 => "0000001010000000000001010000000100",
			3266 => "00000000000100110011001110001001",
			3267 => "00000000100100010011001110001001",
			3268 => "0000000001000000000110000000000100",
			3269 => "00000001010011110011001110001001",
			3270 => "11111111110100110011001110001001",
			3271 => "0000001111000000000111010000001100",
			3272 => "0000000010000000000101001000000100",
			3273 => "00000000000000000011001110001001",
			3274 => "0000000011000000000100010100000100",
			3275 => "00000001001101010011001110001001",
			3276 => "00000100101001000011001110001001",
			3277 => "0000001000000000000111000000001000",
			3278 => "0000000100000000000011011000000100",
			3279 => "00000000101011010011001110001001",
			3280 => "00000011110000100011001110001001",
			3281 => "0000000010000000000100101000000100",
			3282 => "11111110001011110011001110001001",
			3283 => "11111111101010010011001110001001",
			3284 => "11111110011010110011001110001001",
			3285 => "0000001100000000001010111100011000",
			3286 => "0000000011000000001100111000010000",
			3287 => "0000000111000000001101111000001100",
			3288 => "0000000110000000001011001100000100",
			3289 => "11111110101010000011001110001001",
			3290 => "0000000110000000001001100100000100",
			3291 => "00000001010011100011001110001001",
			3292 => "11111111111100100011001110001001",
			3293 => "11111110011011000011001110001001",
			3294 => "0000000100000000000011001100000100",
			3295 => "00000011000000010011001110001001",
			3296 => "00000000000000000011001110001001",
			3297 => "11111110011001100011001110001001",
			3298 => "0000000111000000000101101110000000",
			3299 => "0000001001000000001110100000001000",
			3300 => "0000000110000000001101111100000100",
			3301 => "11111110010101000011010100001101",
			3302 => "00000001010101000011010100001101",
			3303 => "0000000100000000001110111001000000",
			3304 => "0000000110000000001101111100100000",
			3305 => "0000000010000000000101110000010000",
			3306 => "0000001111000000001010011100001000",
			3307 => "0000001011000000000000101000000100",
			3308 => "00000000101010110011010100001101",
			3309 => "11111110111000100011010100001101",
			3310 => "0000000011000000000011011100000100",
			3311 => "00000000101001010011010100001101",
			3312 => "00000001011101000011010100001101",
			3313 => "0000000000000000001111000100001000",
			3314 => "0000000100000000001011110000000100",
			3315 => "00000000000000000011010100001101",
			3316 => "11111101111101100011010100001101",
			3317 => "0000000011000000001101111000000100",
			3318 => "11111111101010110011010100001101",
			3319 => "00000001011101100011010100001101",
			3320 => "0000001011000000000101101100010000",
			3321 => "0000000100000000000011001100001000",
			3322 => "0000001010000000000001010000000100",
			3323 => "00000010000011000011010100001101",
			3324 => "00000010111001010011010100001101",
			3325 => "0000001010000000000110011000000100",
			3326 => "11111111111101100011010100001101",
			3327 => "00000001101011100011010100001101",
			3328 => "0000000110000000001101011000001000",
			3329 => "0000000100000000000010010100000100",
			3330 => "00000011001110100011010100001101",
			3331 => "00000000101100010011010100001101",
			3332 => "0000001001000000000101011100000100",
			3333 => "11111111111010000011010100001101",
			3334 => "11111110101001010011010100001101",
			3335 => "0000001001000000000110101000011100",
			3336 => "0000000010000000000110100000010000",
			3337 => "0000000110000000001101111100001000",
			3338 => "0000000110000000000001111000000100",
			3339 => "11111110010110000011010100001101",
			3340 => "00000101011001000011010100001101",
			3341 => "0000000111000000000100010100000100",
			3342 => "11111110001100010011010100001101",
			3343 => "11111111100001000011010100001101",
			3344 => "0000001010000000000110011000000100",
			3345 => "11111110010110000011010100001101",
			3346 => "0000001100000000000000110000000100",
			3347 => "00000100001011110011010100001101",
			3348 => "00000001000100110011010100001101",
			3349 => "0000001110000000001011000100001100",
			3350 => "0000001000000000000010101000001000",
			3351 => "0000001111000000000110110100000100",
			3352 => "00000000010101110011010100001101",
			3353 => "11111110101101100011010100001101",
			3354 => "11111110001110100011010100001101",
			3355 => "0000000100000000001111100000001000",
			3356 => "0000001000000000000001110100000100",
			3357 => "00000000000000000011010100001101",
			3358 => "00000001100011000011010100001101",
			3359 => "0000000111000000001011000100000100",
			3360 => "00000001111000000011010100001101",
			3361 => "11111111100101000011010100001101",
			3362 => "0000001100000000000110000100101100",
			3363 => "0000001101000000000111010000011000",
			3364 => "0000001110000000001000000000000100",
			3365 => "11111110010011100011010100001101",
			3366 => "0000000100000000000110001100001100",
			3367 => "0000001111000000000111100000001000",
			3368 => "0000001110000000000110100100000100",
			3369 => "11111110101110100011010100001101",
			3370 => "00000000100101110011010100001101",
			3371 => "11111110001000010011010100001101",
			3372 => "0000001100000000000011011100000100",
			3373 => "00000010101111010011010100001101",
			3374 => "11111110011010010011010100001101",
			3375 => "0000000100000000001001001100010000",
			3376 => "0000000110000000001111000000001000",
			3377 => "0000000000000000001001101000000100",
			3378 => "11111110011011100011010100001101",
			3379 => "00000100001000110011010100001101",
			3380 => "0000001000000000001111001000000100",
			3381 => "11111110011000110011010100001101",
			3382 => "00000000110011100011010100001101",
			3383 => "11111110010101010011010100001101",
			3384 => "0000001100000000001010111100010100",
			3385 => "0000000111000000000110100100010000",
			3386 => "0000000111000000001101111000001100",
			3387 => "0000000111000000001110001100000100",
			3388 => "11111110011110000011010100001101",
			3389 => "0000001100000000000110000100000100",
			3390 => "00000000110100100011010100001101",
			3391 => "11111110111100010011010100001101",
			3392 => "11111110010110100011010100001101",
			3393 => "00000111010110100011010100001101",
			3394 => "11111110010100100011010100001101",
			3395 => "0000001000000000000111000010011000",
			3396 => "0000001010000000000110011101111000",
			3397 => "0000001010000000000001010000111100",
			3398 => "0000001000000000000110001000100000",
			3399 => "0000001001000000000110101000010000",
			3400 => "0000000111000000000111111000001000",
			3401 => "0000001000000000001011010100000100",
			3402 => "11111111101110000011011011011001",
			3403 => "11111101101101110011011011011001",
			3404 => "0000000100000000000101010100000100",
			3405 => "00000000001011000011011011011001",
			3406 => "00000001010011010011011011011001",
			3407 => "0000001001000000000110101000001000",
			3408 => "0000000110000000000001111000000100",
			3409 => "11111101111110110011011011011001",
			3410 => "11111111010111000011011011011001",
			3411 => "0000001001000000000110101000000100",
			3412 => "00000000101111000011011011011001",
			3413 => "11111111111001100011011011011001",
			3414 => "0000000100000000001110111000010000",
			3415 => "0000001010000000000001010000001000",
			3416 => "0000001100000000000111111000000100",
			3417 => "11111110100111100011011011011001",
			3418 => "00000000001100000011011011011001",
			3419 => "0000000111000000000100010100000100",
			3420 => "11111111010101110011011011011001",
			3421 => "11111101111101000011011011011001",
			3422 => "0000001000000000001111001000000100",
			3423 => "11111110001011010011011011011001",
			3424 => "0000000110000000000001111000000100",
			3425 => "11111110101001110011011011011001",
			3426 => "00000010000100010011011011011001",
			3427 => "0000000100000000000101010100100000",
			3428 => "0000001101000000001010111100010000",
			3429 => "0000000110000000001101111100001000",
			3430 => "0000001001000000000110101000000100",
			3431 => "11111111111000000011011011011001",
			3432 => "11111101111100000011011011011001",
			3433 => "0000001111000000000101110100000100",
			3434 => "00000001011101100011011011011001",
			3435 => "00000000100100110011011011011001",
			3436 => "0000001111000000001101000100001000",
			3437 => "0000001101000000001101010100000100",
			3438 => "11111110011001100011011011011001",
			3439 => "11111111110100110011011011011001",
			3440 => "0000001110000000000001111100000100",
			3441 => "00000010000010000011011011011001",
			3442 => "00000000010001000011011011011001",
			3443 => "0000001100000000000111111000001100",
			3444 => "0000001111000000000010110100001000",
			3445 => "0000001100000000000111111000000100",
			3446 => "00000000000101110011011011011001",
			3447 => "00000000111010000011011011011001",
			3448 => "00000010001011010011011011011001",
			3449 => "0000000000000000000000110000001000",
			3450 => "0000001001000000000111100100000100",
			3451 => "00000001001000100011011011011001",
			3452 => "11111110111101010011011011011001",
			3453 => "0000001101000000001010111100000100",
			3454 => "11111111110110010011011011011001",
			3455 => "00000000011010010011011011011001",
			3456 => "0000001001000000000110101000000100",
			3457 => "00000010001111010011011011011001",
			3458 => "0000001011000000001000111100001000",
			3459 => "0000001110000000000011011100000100",
			3460 => "11111110011100100011011011011001",
			3461 => "11111111101110000011011011011001",
			3462 => "0000001001000000001011101000001000",
			3463 => "0000001110000000001101100000000100",
			3464 => "00000000000000000011011011011001",
			3465 => "00000010010010010011011011011001",
			3466 => "0000001111000000001001010000000100",
			3467 => "11111110100000110011011011011001",
			3468 => "0000000001000000001001111000000100",
			3469 => "00000001110000110011011011011001",
			3470 => "11111110100001110011011011011001",
			3471 => "0000001100000000000111111000011100",
			3472 => "0000000000000000001000111100000100",
			3473 => "11111110101000000011011011011001",
			3474 => "0000001011000000000100010100010000",
			3475 => "0000001001000000001100110100001100",
			3476 => "0000001111000000000100001000000100",
			3477 => "11111111001101000011011011011001",
			3478 => "0000001100000000001010000000000100",
			3479 => "00000001010100000011011011011001",
			3480 => "00000000000000000011011011011001",
			3481 => "11111110111000100011011011011001",
			3482 => "0000001101000000000011011100000100",
			3483 => "11111111010111010011011011011001",
			3484 => "00000010111010110011011011011001",
			3485 => "0000000111000000001011000100010100",
			3486 => "0000000100000000000010010000001000",
			3487 => "0000001101000000001001110000000100",
			3488 => "11111111010010100011011011011001",
			3489 => "11111110001011100011011011011001",
			3490 => "0000000110000000000100110100001000",
			3491 => "0000000000000000001101111000000100",
			3492 => "00000001001101100011011011011001",
			3493 => "00000000000000000011011011011001",
			3494 => "11111111010110000011011011011001",
			3495 => "0000000001000000001110100000010000",
			3496 => "0000001010000000000101000100000100",
			3497 => "11111110100000000011011011011001",
			3498 => "0000001010000000000001010100000100",
			3499 => "00000001100111000011011011011001",
			3500 => "0000001001000000000010001100000100",
			3501 => "11111110110011010011011011011001",
			3502 => "00000000010101110011011011011001",
			3503 => "0000000000000000000000101000000100",
			3504 => "00000001000000110011011011011001",
			3505 => "0000001011000000001100001000000100",
			3506 => "00000000000000110011011011011001",
			3507 => "0000000100000000001111100000000100",
			3508 => "00000000000000000011011011011001",
			3509 => "11111110010111010011011011011001",
			3510 => "0000001100000000000110000101111100",
			3511 => "0000000100000000000011111001111000",
			3512 => "0000001100000000000000101001000000",
			3513 => "0000001100000000000100010100100000",
			3514 => "0000001100000000000100010100010000",
			3515 => "0000000111000000001011000100001000",
			3516 => "0000001011000000000100000000000100",
			3517 => "00000000101011000011100000011101",
			3518 => "00000010011000110011100000011101",
			3519 => "0000000111000000000000101000000100",
			3520 => "11111111110001100011100000011101",
			3521 => "00000000100110000011100000011101",
			3522 => "0000000111000000001100001000001000",
			3523 => "0000000111000000001100001000000100",
			3524 => "11111111010011000011100000011101",
			3525 => "00000010001110010011100000011101",
			3526 => "0000000111000000001100001000000100",
			3527 => "11111110001001000011100000011101",
			3528 => "11111111101110100011100000011101",
			3529 => "0000001100000000000100010100010000",
			3530 => "0000000111000000001100001000001000",
			3531 => "0000000111000000000000101000000100",
			3532 => "00000001111100000011100000011101",
			3533 => "11111111011100100011100000011101",
			3534 => "0000001011000000001100001000000100",
			3535 => "00000011110000110011100000011101",
			3536 => "00000001111011110011100000011101",
			3537 => "0000000100000000000100001100001000",
			3538 => "0000001100000000000100010100000100",
			3539 => "11111110111001000011100000011101",
			3540 => "00000000110101010011100000011101",
			3541 => "0000000001000000001110100000000100",
			3542 => "00000001001001110011100000011101",
			3543 => "11111110110101000011100000011101",
			3544 => "0000001100000000000000101000011000",
			3545 => "0000001101000000001010111100010000",
			3546 => "0000000110000000001100011000001000",
			3547 => "0000000010000000000111111100000100",
			3548 => "11111111001011000011100000011101",
			3549 => "11111101011010110011100000011101",
			3550 => "0000001110000000000110000100000100",
			3551 => "11111110111111110011100000011101",
			3552 => "00000001100001100011100000011101",
			3553 => "0000001101000000000111001000000100",
			3554 => "11111100111100100011100000011101",
			3555 => "11111110001011010011100000011101",
			3556 => "0000000110000000000100110100010000",
			3557 => "0000000100000000000110001100001000",
			3558 => "0000001010000000001000010100000100",
			3559 => "11111111101010010011100000011101",
			3560 => "00000001100011110011100000011101",
			3561 => "0000001110000000000101101100000100",
			3562 => "11111111001110010011100000011101",
			3563 => "11111101011111110011100000011101",
			3564 => "0000001010000000000110011000001000",
			3565 => "0000000100000000000011001100000100",
			3566 => "00000001000101110011100000011101",
			3567 => "11111111001000000011100000011101",
			3568 => "0000001001000000001111001100000100",
			3569 => "00000000011100100011100000011101",
			3570 => "11111111100100100011100000011101",
			3571 => "11111110011001000011100000011101",
			3572 => "0000001100000000001010111100100100",
			3573 => "0000000111000000001011000000011000",
			3574 => "0000000111000000000100011000010000",
			3575 => "0000000111000000001101111000001100",
			3576 => "0000000111000000001110001100000100",
			3577 => "11111110110000100011100000011101",
			3578 => "0000001100000000000110000100000100",
			3579 => "00000000010110100011100000011101",
			3580 => "11111111111101110011100000011101",
			3581 => "11111110011001100011100000011101",
			3582 => "0000001100000000000100001000000100",
			3583 => "00000011001100110011100000011101",
			3584 => "11111110100111100011100000011101",
			3585 => "0000000100000000000010010100000100",
			3586 => "11111110111001010011100000011101",
			3587 => "0000001010000000000001010000000100",
			3588 => "00000011110100110011100000011101",
			3589 => "11111111111010110011100000011101",
			3590 => "11111110011000100011100000011101",
			3591 => "0000001100000000000110000110101100",
			3592 => "0000001010000000001001000101101000",
			3593 => "0000000100000000001100001100101100",
			3594 => "0000000100000000001100001100100000",
			3595 => "0000000100000000001110000000010000",
			3596 => "0000001000000000001001101000001000",
			3597 => "0000001010000000000011101000000100",
			3598 => "11111111110101000011100110010001",
			3599 => "00000000101110100011100110010001",
			3600 => "0000000010000000001111010000000100",
			3601 => "00000000010101100011100110010001",
			3602 => "11111011111100110011100110010001",
			3603 => "0000000000000000001111000100001000",
			3604 => "0000000001000000001100110100000100",
			3605 => "11111111111110100011100110010001",
			3606 => "11111101111110100011100110010001",
			3607 => "0000001110000000001000111000000100",
			3608 => "11111111110100000011100110010001",
			3609 => "00000000101111110011100110010001",
			3610 => "0000001001000000000111100100001000",
			3611 => "0000001011000000000000101000000100",
			3612 => "00000011000000100011100110010001",
			3613 => "11111110100001000011100110010001",
			3614 => "00000010101010000011100110010001",
			3615 => "0000001111000000001011011100011100",
			3616 => "0000000001000000001110100000001100",
			3617 => "0000001110000000001110111100001000",
			3618 => "0000000111000000000000101000000100",
			3619 => "00000000110100000011100110010001",
			3620 => "11111110010011100011100110010001",
			3621 => "00000011011100110011100110010001",
			3622 => "0000001100000000000100010100001000",
			3623 => "0000001111000000000001011000000100",
			3624 => "11111111110110000011100110010001",
			3625 => "11111110000011100011100110010001",
			3626 => "0000001000000000001001101000000100",
			3627 => "00000000010010110011100110010001",
			3628 => "00000011001001010011100110010001",
			3629 => "0000001101000000001100101100010000",
			3630 => "0000001011000000000100010100001000",
			3631 => "0000000000000000000011111100000100",
			3632 => "11111110010001000011100110010001",
			3633 => "00000001101101110011100110010001",
			3634 => "0000001110000000000000101000000100",
			3635 => "11111101101110010011100110010001",
			3636 => "11111110100101110011100110010001",
			3637 => "0000001100000000000000101000001000",
			3638 => "0000001110000000001100101100000100",
			3639 => "00000000000011100011100110010001",
			3640 => "11111101101100110011100110010001",
			3641 => "0000001100000000000000101000000100",
			3642 => "11111110000010010011100110010001",
			3643 => "11111111101110110011100110010001",
			3644 => "0000000000000000001111000100010100",
			3645 => "0000001101000000000100011000000100",
			3646 => "11111011101110100011100110010001",
			3647 => "0000000010000000000010000000000100",
			3648 => "00000001101111110011100110010001",
			3649 => "0000001000000000001001101000001000",
			3650 => "0000001000000000001001101000000100",
			3651 => "11111110010110000011100110010001",
			3652 => "00000000101100110011100110010001",
			3653 => "11111110001111010011100110010001",
			3654 => "0000000100000000000011001100010000",
			3655 => "0000000000000000000000110000001100",
			3656 => "0000000001000000000110000000000100",
			3657 => "11111110001010110011100110010001",
			3658 => "0000001100000000001010000000000100",
			3659 => "11111110110101110011100110010001",
			3660 => "00000000101100110011100110010001",
			3661 => "11111101101101000011100110010001",
			3662 => "0000000111000000001100001000010000",
			3663 => "0000000111000000000000101000001000",
			3664 => "0000000111000000000000101000000100",
			3665 => "00000000011000000011100110010001",
			3666 => "11111111010110010011100110010001",
			3667 => "0000001111000000001011011100000100",
			3668 => "00000010011011000011100110010001",
			3669 => "00000000101010010011100110010001",
			3670 => "0000001000000000000110001000001000",
			3671 => "0000001111000000001001010100000100",
			3672 => "11111111010010100011100110010001",
			3673 => "11111110010100100011100110010001",
			3674 => "0000000111000000001100001000000100",
			3675 => "11111111100111110011100110010001",
			3676 => "00000000010010010011100110010001",
			3677 => "0000001100000000001010111100001100",
			3678 => "0000000000000000000111000100001000",
			3679 => "0000000000000000001111001000000100",
			3680 => "11111110101100010011100110010001",
			3681 => "00000010100011000011100110010001",
			3682 => "11111110011101000011100110010001",
			3683 => "11111110011001110011100110010001",
			3684 => "0000000011000000000100000010000000",
			3685 => "0000000100000000000011010100111000",
			3686 => "0000000000000000000100010100101000",
			3687 => "0000000011000000000100000000011000",
			3688 => "0000000010000000001111010000010000",
			3689 => "0000001111000000000100000100001000",
			3690 => "0000001000000000000111000100000100",
			3691 => "11111111100110000011101110000101",
			3692 => "00000000100011110011101110000101",
			3693 => "0000000101000000001001110000000100",
			3694 => "11111110111001000011101110000101",
			3695 => "00000001101111010011101110000101",
			3696 => "0000001101000000001001110000000100",
			3697 => "00000000111100000011101110000101",
			3698 => "11111110000101110011101110000101",
			3699 => "0000000111000000000111111000000100",
			3700 => "00000000011000010011101110000101",
			3701 => "0000001111000000000100000100001000",
			3702 => "0000001101000000000101101100000100",
			3703 => "00000000100000010011101110000101",
			3704 => "11111110101010000011101110000101",
			3705 => "11111110000101110011101110000101",
			3706 => "0000000110000000000100110100000100",
			3707 => "11111110001110000011101110000101",
			3708 => "0000001101000000001101100000000100",
			3709 => "00000001010001010011101110000101",
			3710 => "0000001101000000001100101100000100",
			3711 => "11111110100011100011101110000101",
			3712 => "00000000000000000011101110000101",
			3713 => "0000000100000000000011110100010100",
			3714 => "0000000001000000001110100000010000",
			3715 => "0000001010000000001100011100001100",
			3716 => "0000001000000000000001110100001000",
			3717 => "0000000110000000001101111100000100",
			3718 => "00000010101010100011101110000101",
			3719 => "00000000111011110011101110000101",
			3720 => "11111111001000010011101110000101",
			3721 => "00000010100001100011101110000101",
			3722 => "11111110100010100011101110000101",
			3723 => "0000000001000000000110000000011100",
			3724 => "0000001111000000001110110000010000",
			3725 => "0000001101000000000100000000001000",
			3726 => "0000001100000000001010000000000100",
			3727 => "11111111111100010011101110000101",
			3728 => "00000000110101110011101110000101",
			3729 => "0000000010000000001100100100000100",
			3730 => "11111110011010110011101110000101",
			3731 => "00000000000000000011101110000101",
			3732 => "0000001100000000000100010100001000",
			3733 => "0000001111000000000000011100000100",
			3734 => "00000001101010000011101110000101",
			3735 => "00000000000000000011101110000101",
			3736 => "11111110110000100011101110000101",
			3737 => "0000000010000000001100100100001100",
			3738 => "0000000011000000000111111000001000",
			3739 => "0000001010000000000101000100000100",
			3740 => "11111110100000110011101110000101",
			3741 => "00000000110110110011101110000101",
			3742 => "00000010100010010011101110000101",
			3743 => "0000001001000000000110101000001000",
			3744 => "0000000100000000000011011000000100",
			3745 => "11111111000101110011101110000101",
			3746 => "00000000001000100011101110000101",
			3747 => "00000010000000110011101110000101",
			3748 => "0000001001000000000010001100010100",
			3749 => "0000000110000000000001111000000100",
			3750 => "11111110001111100011101110000101",
			3751 => "0000000110000000001101111100000100",
			3752 => "00000010011111000011101110000101",
			3753 => "0000000110000000000100110100000100",
			3754 => "00000000000000000011101110000101",
			3755 => "0000000011000000001001110000000100",
			3756 => "00000000000010100011101110000101",
			3757 => "00000010001001110011101110000101",
			3758 => "0000001111000000000001011000101100",
			3759 => "0000001001000000000110101000010000",
			3760 => "0000000001000000001110100000001100",
			3761 => "0000000101000000000101101100001000",
			3762 => "0000000111000000001011000100000100",
			3763 => "00000000010111110011101110000101",
			3764 => "00000001111010110011101110000101",
			3765 => "11111110101111110011101110000101",
			3766 => "00000010101001010011101110000101",
			3767 => "0000001101000000001110001100010000",
			3768 => "0000001111000000000000011100001000",
			3769 => "0000001000000000001001101000000100",
			3770 => "11111110101000010011101110000101",
			3771 => "00000000000000000011101110000101",
			3772 => "0000000011000000000011011100000100",
			3773 => "00000001110101000011101110000101",
			3774 => "00000000010101010011101110000101",
			3775 => "0000001100000000000111111000000100",
			3776 => "11111110101001110011101110000101",
			3777 => "0000001101000000001101111000000100",
			3778 => "00000001100001110011101110000101",
			3779 => "00000000001100110011101110000101",
			3780 => "0000000110000000001101111100100000",
			3781 => "0000000011000000001110001100010000",
			3782 => "0000000101000000001100101100001000",
			3783 => "0000000100000000000010111000000100",
			3784 => "00000000010110100011101110000101",
			3785 => "11111111000100000011101110000101",
			3786 => "0000000100000000001110000000000100",
			3787 => "00000000000111100011101110000101",
			3788 => "11111110011011000011101110000101",
			3789 => "0000000011000000001010111100001000",
			3790 => "0000001100000000000100000000000100",
			3791 => "00000000111100110011101110000101",
			3792 => "11111110001010100011101110000101",
			3793 => "0000000001000000001001111000000100",
			3794 => "11111110110110000011101110000101",
			3795 => "00000000100100110011101110000101",
			3796 => "0000000010000000001100100100001100",
			3797 => "0000000101000000001110001100000100",
			3798 => "11111101010000100011101110000101",
			3799 => "0000001000000000001100000100000100",
			3800 => "11111110010110000011101110000101",
			3801 => "00000000101010000011101110000101",
			3802 => "0000001101000000000101101100001000",
			3803 => "0000000010000000000101001000000100",
			3804 => "00000010100001010011101110000101",
			3805 => "00000000010101100011101110000101",
			3806 => "0000000011000000000011011100000100",
			3807 => "11111111100000100011101110000101",
			3808 => "00000000000101010011101110000101",
			3809 => "0000000010000000000110010010010100",
			3810 => "0000000100000000000011011001010100",
			3811 => "0000000000000000001100001000110100",
			3812 => "0000000101000000001000111100010100",
			3813 => "0000000101000000001000111100010000",
			3814 => "0000000010000000001110000100001000",
			3815 => "0000000110000000000001111000000100",
			3816 => "00000000101010100011110111000001",
			3817 => "11111110100011100011110111000001",
			3818 => "0000000011000000000100010100000100",
			3819 => "00000001000100010011110111000001",
			3820 => "00000010110111100011110111000001",
			3821 => "00000011000110100011110111000001",
			3822 => "0000001011000000000111111000010000",
			3823 => "0000000100000000000000010100001000",
			3824 => "0000001101000000001101100000000100",
			3825 => "11111110011101000011110111000001",
			3826 => "00000000000000000011110111000001",
			3827 => "0000000111000000000111111000000100",
			3828 => "00000000111011110011110111000001",
			3829 => "11111110101111010011110111000001",
			3830 => "0000001001000000001001111000001000",
			3831 => "0000000011000000001100001000000100",
			3832 => "00000000001011110011110111000001",
			3833 => "00000001010010100011110111000001",
			3834 => "0000000110000000000100110100000100",
			3835 => "11111111111011100011110111000001",
			3836 => "00000000001010110011110111000001",
			3837 => "0000001110000000000000101000011000",
			3838 => "0000001011000000000111111000001100",
			3839 => "0000000101000000001000111100001000",
			3840 => "0000000101000000001000111100000100",
			3841 => "11111110010001110011110111000001",
			3842 => "11111111100001100011110111000001",
			3843 => "00000001001101010011110111000001",
			3844 => "0000001010000000000001010100001000",
			3845 => "0000000111000000000000101000000100",
			3846 => "11111110001100010011110111000001",
			3847 => "11111111000011110011110111000001",
			3848 => "00000000000000000011110111000001",
			3849 => "0000001110000000000100000000000100",
			3850 => "00000011000101100011110111000001",
			3851 => "11111110101010000011110111000001",
			3852 => "0000000100000000000001100100100100",
			3853 => "0000001010000000000110011100001100",
			3854 => "0000001011000000000111111000001000",
			3855 => "0000000111000000001010000000000100",
			3856 => "00000000000000000011110111000001",
			3857 => "00000011010000000011110111000001",
			3858 => "11111110100001110011110111000001",
			3859 => "0000001010000000000101000100001000",
			3860 => "0000001100000000000100010100000100",
			3861 => "00000001011011000011110111000001",
			3862 => "00000011010111110011110111000001",
			3863 => "0000000100000000000000100000001000",
			3864 => "0000001000000000001000110000000100",
			3865 => "11111110011001100011110111000001",
			3866 => "00000000111000000011110111000001",
			3867 => "0000000010000000000001000000000100",
			3868 => "00000010010110110011110111000001",
			3869 => "00000000101101010011110111000001",
			3870 => "0000000010000000001001010000001100",
			3871 => "0000000101000000001000111100001000",
			3872 => "0000001110000000000101000100000100",
			3873 => "11111110110111100011110111000001",
			3874 => "00000001011010000011110111000001",
			3875 => "11111110001011110011110111000001",
			3876 => "0000000010000000001010001000001100",
			3877 => "0000001110000000000010101000001000",
			3878 => "0000000110000000000100110100000100",
			3879 => "00000001000000110011110111000001",
			3880 => "11111110111000100011110111000001",
			3881 => "00000010000110110011110111000001",
			3882 => "11111110100000100011110111000001",
			3883 => "0000000110000000001010011001000000",
			3884 => "0000000101000000001101100000010100",
			3885 => "0000000100000000001011100000001000",
			3886 => "0000000000000000000011111100000100",
			3887 => "00000000000000000011110111000001",
			3888 => "00000010101101110011110111000001",
			3889 => "0000000000000000000000101000001000",
			3890 => "0000000111000000000111111000000100",
			3891 => "00000000000000000011110111000001",
			3892 => "00000000110011110011110111000001",
			3893 => "11111110011111100011110111000001",
			3894 => "0000000111000000001000111000011000",
			3895 => "0000001100000000000100000000010000",
			3896 => "0000000101000000001100101000001000",
			3897 => "0000001011000000001000111100000100",
			3898 => "11111111010001100011110111000001",
			3899 => "11111101101110100011110111000001",
			3900 => "0000000010000000001001100000000100",
			3901 => "00000001011100110011110111000001",
			3902 => "11111111000111110011110111000001",
			3903 => "0000000010000000001110110100000100",
			3904 => "11111101001011110011110111000001",
			3905 => "11111110100110010011110111000001",
			3906 => "0000000000000000000011111100001100",
			3907 => "0000000010000000001110110100000100",
			3908 => "11111101101101010011110111000001",
			3909 => "0000000110000000001010011000000100",
			3910 => "11111111010001110011110111000001",
			3911 => "00000001100101010011110111000001",
			3912 => "0000000100000000001111100000000100",
			3913 => "00000010000100110011110111000001",
			3914 => "11111110100101100011110111000001",
			3915 => "0000000110000000001010011000001100",
			3916 => "0000000111000000000101101100000100",
			3917 => "00000010100000100011110111000001",
			3918 => "0000001001000000001010011000000100",
			3919 => "11111110100101100011110111000001",
			3920 => "00000000000000000011110111000001",
			3921 => "0000001000000000001111001000100000",
			3922 => "0000000110000000001101011000010000",
			3923 => "0000000100000000000010110000001000",
			3924 => "0000000010000000000010000100000100",
			3925 => "00000000110110000011110111000001",
			3926 => "11111110011000000011110111000001",
			3927 => "0000000010000000000111011000000100",
			3928 => "11111101000011010011110111000001",
			3929 => "11111111010110010011110111000001",
			3930 => "0000000011000000000000011100001000",
			3931 => "0000001100000000000100000000000100",
			3932 => "11111111111001000011110111000001",
			3933 => "00000001111001000011110111000001",
			3934 => "0000000101000000001000011000000100",
			3935 => "11111110101101100011110111000001",
			3936 => "00000000000000000011110111000001",
			3937 => "0000000100000000001001001100010000",
			3938 => "0000000111000000001001110000001000",
			3939 => "0000001100000000000100000000000100",
			3940 => "00000000101101000011110111000001",
			3941 => "00000010001111010011110111000001",
			3942 => "0000001000000000000111000100000100",
			3943 => "00000010001001110011110111000001",
			3944 => "11111110100100110011110111000001",
			3945 => "0000000000000000001110111100001000",
			3946 => "0000000010000000001100010000000100",
			3947 => "11111110001000100011110111000001",
			3948 => "11111111100111110011110111000001",
			3949 => "0000000100000000000100001100000100",
			3950 => "00000000110011000011110111000001",
			3951 => "11111111110000010011110111000001",
			3952 => "0000001100000000001000111010111000",
			3953 => "0000001100000000000111111001101100",
			3954 => "0000001100000000000111111001000000",
			3955 => "0000001100000000000111111000100000",
			3956 => "0000000010000000001110010000010000",
			3957 => "0000000111000000000100010100001000",
			3958 => "0000000111000000000100010100000100",
			3959 => "11111111110001110011111110111101",
			3960 => "00000000111111000011111110111101",
			3961 => "0000000010000000001001010000000100",
			3962 => "11111111110001100011111110111101",
			3963 => "11111110110010110011111110111101",
			3964 => "0000000100000000001011100000001000",
			3965 => "0000001111000000001011110100000100",
			3966 => "00000011001111010011111110111101",
			3967 => "00000000110010100011111110111101",
			3968 => "0000000110000000000100110100000100",
			3969 => "00000000000000000011111110111101",
			3970 => "11111110000101010011111110111101",
			3971 => "0000001100000000000111111000010000",
			3972 => "0000001001000000000110101000001000",
			3973 => "0000001101000000001001110000000100",
			3974 => "11111111001001110011111110111101",
			3975 => "00000010001101110011111110111101",
			3976 => "0000001101000000001110001100000100",
			3977 => "11111111001111110011111110111101",
			3978 => "00000010010110100011111110111101",
			3979 => "0000000111000000000100010100001000",
			3980 => "0000000111000000000111111000000100",
			3981 => "00000000011000100011111110111101",
			3982 => "00000011000010110011111110111101",
			3983 => "0000000111000000000100010100000100",
			3984 => "11111101110001000011111110111101",
			3985 => "00000000001010010011111110111101",
			3986 => "0000001100000000000111111000010000",
			3987 => "0000000111000000000111111000000100",
			3988 => "00000001000101100011111110111101",
			3989 => "0000001001000000000111100100001000",
			3990 => "0000000011000000000101101100000100",
			3991 => "11111111000010000011111110111101",
			3992 => "11111101011101000011111110111101",
			3993 => "00000000011111010011111110111101",
			3994 => "0000000111000000000000101000010000",
			3995 => "0000000111000000000111111000001000",
			3996 => "0000000001000000000110000000000100",
			3997 => "00000000011011010011111110111101",
			3998 => "11111101110100110011111110111101",
			3999 => "0000000010000000000010110100000100",
			4000 => "11111110000110000011111110111101",
			4001 => "00000000011111100011111110111101",
			4002 => "0000000111000000000000101000000100",
			4003 => "11111101111011010011111110111101",
			4004 => "0000001011000000000000101000000100",
			4005 => "00000000101000010011111110111101",
			4006 => "11111111000110000011111110111101",
			4007 => "0000001100000000000100010100100000",
			4008 => "0000000000000000001000110000000100",
			4009 => "11111110101001000011111110111101",
			4010 => "0000000001000000001100110100010000",
			4011 => "0000000111000000000000101000001000",
			4012 => "0000001101000000001100110000000100",
			4013 => "11111111111110110011111110111101",
			4014 => "00000001010001100011111110111101",
			4015 => "0000000000000000000000111000000100",
			4016 => "11111101101010000011111110111101",
			4017 => "11111111111001010011111110111101",
			4018 => "0000001011000000001000111100001000",
			4019 => "0000000011000000000110000100000100",
			4020 => "00000010100111110011111110111101",
			4021 => "00000001110110100011111110111101",
			4022 => "00000000100010010011111110111101",
			4023 => "0000000001000000000110000000010000",
			4024 => "0000000011000000000011010000001000",
			4025 => "0000000010000000001110101000000100",
			4026 => "11111111001001100011111110111101",
			4027 => "00000010000100010011111110111101",
			4028 => "0000001101000000000101101100000100",
			4029 => "11111110001100110011111110111101",
			4030 => "11111111100010000011111110111101",
			4031 => "0000001101000000001101100000001100",
			4032 => "0000001100000000000100010100000100",
			4033 => "11111110001011110011111110111101",
			4034 => "0000000010000000001001010000000100",
			4035 => "00000001111101010011111110111101",
			4036 => "00000000001000010011111110111101",
			4037 => "0000000011000000001100110000001000",
			4038 => "0000001101000000001101111000000100",
			4039 => "11111111110111110011111110111101",
			4040 => "11111101111011110011111110111101",
			4041 => "0000001001000000000111100100000100",
			4042 => "00000000011010100011111110111101",
			4043 => "00000000000000100011111110111101",
			4044 => "0000001111000000001101000100001100",
			4045 => "0000000000000000000011010000001000",
			4046 => "0000001011000000001100101100000100",
			4047 => "00000000100110000011111110111101",
			4048 => "11111101111111000011111110111101",
			4049 => "11111110001001000011111110111101",
			4050 => "0000000001000000000110101000011100",
			4051 => "0000000101000000001001110100010000",
			4052 => "0000001010000000000110011100001100",
			4053 => "0000001010000000001010110000001000",
			4054 => "0000001010000000000001010000000100",
			4055 => "11111110001110100011111110111101",
			4056 => "00000001111110110011111110111101",
			4057 => "11111110010000010011111110111101",
			4058 => "00000010011011110011111110111101",
			4059 => "0000001011000000000001111100001000",
			4060 => "0000000011000000000001101000000100",
			4061 => "00000000000000000011111110111101",
			4062 => "00000010111101110011111110111101",
			4063 => "00000000000000000011111110111101",
			4064 => "0000000000000000000111000100010000",
			4065 => "0000001100000000001010111100001100",
			4066 => "0000000000000000001001101000000100",
			4067 => "00000000000000000011111110111101",
			4068 => "0000000001000000001110010100000100",
			4069 => "00000001101000000011111110111101",
			4070 => "00000000000000000011111110111101",
			4071 => "11111110110000100011111110111101",
			4072 => "0000000111000000001110001100000100",
			4073 => "11111110010010000011111110111101",
			4074 => "0000000111000000001101111000001000",
			4075 => "0000000010000000001011101100000100",
			4076 => "00000001001010010011111110111101",
			4077 => "00000000000000000011111110111101",
			4078 => "11111110100011110011111110111101",
			4079 => "0000001010000000000001010010010000",
			4080 => "0000001000000000001111001001110000",
			4081 => "0000000000000000000011010000111000",
			4082 => "0000000010000000000110010000100000",
			4083 => "0000001010000000001001000100010000",
			4084 => "0000000110000000001010011000001000",
			4085 => "0000000001000000001001111000000100",
			4086 => "11111111111101000100000111111001",
			4087 => "00000000101000000100000111111001",
			4088 => "0000000101000000000100011000000100",
			4089 => "11111101111101000100000111111001",
			4090 => "00000000000011000100000111111001",
			4091 => "0000000110000000001101111100001000",
			4092 => "0000001110000000000100010100000100",
			4093 => "11111111101001000100000111111001",
			4094 => "00000001111110100100000111111001",
			4095 => "0000000011000000001110001100000100",
			4096 => "11111110101101000100000111111001",
			4097 => "00000000011010000100000111111001",
			4098 => "0000001111000000000101001000001000",
			4099 => "0000000111000000000100000000000100",
			4100 => "11111111100000110100000111111001",
			4101 => "11111101010110100100000111111001",
			4102 => "0000001010000000000110011000001000",
			4103 => "0000001010000000000110011000000100",
			4104 => "11111111100010000100000111111001",
			4105 => "00000001011100100100000111111001",
			4106 => "0000000101000000001000011000000100",
			4107 => "11111110011110000100000111111001",
			4108 => "00000001000101010100000111111001",
			4109 => "0000001011000000001100001000011000",
			4110 => "0000001011000000001100001000010000",
			4111 => "0000000000000000000000111000001000",
			4112 => "0000001000000000000110001000000100",
			4113 => "00000000000010010100000111111001",
			4114 => "00000001010010100100000111111001",
			4115 => "0000001000000000001111001000000100",
			4116 => "11111111100110010100000111111001",
			4117 => "00000001000000110100000111111001",
			4118 => "0000001000000000000110001000000100",
			4119 => "00000000000000000100000111111001",
			4120 => "00000010110111100100000111111001",
			4121 => "0000001110000000000100000000010000",
			4122 => "0000001101000000001110001100001000",
			4123 => "0000000010000000000101110000000100",
			4124 => "11111111101101000100000111111001",
			4125 => "11111110010101010100000111111001",
			4126 => "0000000110000000000100110100000100",
			4127 => "11111101111110010100000111111001",
			4128 => "00000000111101100100000111111001",
			4129 => "0000001001000000001011101000001000",
			4130 => "0000001101000000001101111000000100",
			4131 => "11111111011000100100000111111001",
			4132 => "00000000001011010100000111111001",
			4133 => "0000001011000000000110000100000100",
			4134 => "11111110011000000100000111111001",
			4135 => "00000000001110000100000111111001",
			4136 => "0000001101000000001100110000010100",
			4137 => "0000000101000000000011011100010000",
			4138 => "0000000001000000000110000000001000",
			4139 => "0000000000000000000000101000000100",
			4140 => "00000010000001110100000111111001",
			4141 => "00000000000000000100000111111001",
			4142 => "0000000000000000001110111100000100",
			4143 => "11111111001010110100000111111001",
			4144 => "11111101111011000100000111111001",
			4145 => "00000000110111100100000111111001",
			4146 => "0000000111000000001100001000000100",
			4147 => "11111101100101010100000111111001",
			4148 => "0000001111000000000111110000000100",
			4149 => "11111111100011000100000111111001",
			4150 => "11111110010000000100000111111001",
			4151 => "0000000011000000001110111100110100",
			4152 => "0000001010000000000101000100011000",
			4153 => "0000001001000000001100110100010000",
			4154 => "0000001111000000000100011000000100",
			4155 => "11111110010110110100000111111001",
			4156 => "0000000101000000001000111100001000",
			4157 => "0000000011000000000011111100000100",
			4158 => "00000000000000000100000111111001",
			4159 => "00000001111111110100000111111001",
			4160 => "11111111101011100100000111111001",
			4161 => "0000001111000000001010111000000100",
			4162 => "00000000001000010100000111111001",
			4163 => "11111110001110110100000111111001",
			4164 => "0000000110000000001010011000011000",
			4165 => "0000000000000000001100110000001000",
			4166 => "0000001000000000001000110000000100",
			4167 => "00000000010010100100000111111001",
			4168 => "00000010001101010100000111111001",
			4169 => "0000000011000000000000110000001000",
			4170 => "0000000101000000001001110000000100",
			4171 => "00000000000111110100000111111001",
			4172 => "11111110010000100100000111111001",
			4173 => "0000000010000000000110010000000100",
			4174 => "00000001001110000100000111111001",
			4175 => "00000000000000000100000111111001",
			4176 => "11111110011011000100000111111001",
			4177 => "0000000010000000001111010000101000",
			4178 => "0000000000000000001011000100011000",
			4179 => "0000001110000000001101010000001000",
			4180 => "0000000010000000001100100100000100",
			4181 => "00000011100110010100000111111001",
			4182 => "00000000011111100100000111111001",
			4183 => "0000001000000000000001110100001000",
			4184 => "0000000001000000001110100000000100",
			4185 => "11111111110101100100000111111001",
			4186 => "00000000111110000100000111111001",
			4187 => "0000001111000000000111010000000100",
			4188 => "00000010110001100100000111111001",
			4189 => "11111111111001010100000111111001",
			4190 => "0000000011000000001011000100001000",
			4191 => "0000000001000000000110000000000100",
			4192 => "11111111110101110100000111111001",
			4193 => "11111110010010110100000111111001",
			4194 => "0000000001000000001110100000000100",
			4195 => "00000001011000000100000111111001",
			4196 => "11111110100110010100000111111001",
			4197 => "0000000010000000001001010000010100",
			4198 => "0000000110000000000100110100001000",
			4199 => "0000000010000000001111010000000100",
			4200 => "11111101101001110100000111111001",
			4201 => "11111111100000000100000111111001",
			4202 => "0000000001000000001110100000000100",
			4203 => "00000001010110110100000111111001",
			4204 => "0000000001000000001100110100000100",
			4205 => "11111110000011000100000111111001",
			4206 => "11111111111011110100000111111001",
			4207 => "0000001101000000001100110000010000",
			4208 => "0000001110000000000111111000001000",
			4209 => "0000000111000000000111111000000100",
			4210 => "00000000011001000100000111111001",
			4211 => "11111111100001110100000111111001",
			4212 => "0000000011000000001101100000000100",
			4213 => "11111101101000010100000111111001",
			4214 => "11111111011010110100000111111001",
			4215 => "0000001001000000000111100100001000",
			4216 => "0000000011000000000101101100000100",
			4217 => "00000000000101100100000111111001",
			4218 => "00000000101011100100000111111001",
			4219 => "0000000001000000001100110100000100",
			4220 => "11111111001001010100000111111001",
			4221 => "00000000000100000100000111111001",
			4222 => "0000001010000000000110011010101100",
			4223 => "0000001100000000000100010101010000",
			4224 => "0000000111000000001011000100100000",
			4225 => "0000000101000000001100101100011000",
			4226 => "0000000110000000001101111100001100",
			4227 => "0000000111000000001011000100001000",
			4228 => "0000000111000000001011000100000100",
			4229 => "00000000000110110100010000011101",
			4230 => "11111110100001100100010000011101",
			4231 => "00000010011010010100010000011101",
			4232 => "0000001011000000001100001000001000",
			4233 => "0000000100000000000010110000000100",
			4234 => "11111101011111010100010000011101",
			4235 => "11111111010000010100010000011101",
			4236 => "00000000000101100100010000011101",
			4237 => "0000000111000000001011000100000100",
			4238 => "00000000100110100100010000011101",
			4239 => "00000010011110100100010000011101",
			4240 => "0000001100000000000100010100100000",
			4241 => "0000000001000000001100110100010000",
			4242 => "0000000100000000000011001100001000",
			4243 => "0000000000000000000010111100000100",
			4244 => "11111111100010000100010000011101",
			4245 => "00000000101011010100010000011101",
			4246 => "0000000100000000000010111000000100",
			4247 => "11111101001111010100010000011101",
			4248 => "11111111001111010100010000011101",
			4249 => "0000001011000000001000111100001000",
			4250 => "0000000110000000000100110100000100",
			4251 => "11111110001010010100010000011101",
			4252 => "00000000010000010100010000011101",
			4253 => "0000000111000000001100001000000100",
			4254 => "11111111011001000100010000011101",
			4255 => "00000001011110100100010000011101",
			4256 => "0000000111000000001100001000001000",
			4257 => "0000000001000000001100110100000100",
			4258 => "11111110100111110100010000011101",
			4259 => "11111101000100010100010000011101",
			4260 => "0000001011000000000100000000000100",
			4261 => "00000000010011110100010000011101",
			4262 => "11111110001110110100010000011101",
			4263 => "0000001100000000000100010100100100",
			4264 => "0000000001000000001110100000010000",
			4265 => "0000001011000000001011000100001000",
			4266 => "0000001001000000001001111000000100",
			4267 => "11111111100010110100010000011101",
			4268 => "11111101111100010100010000011101",
			4269 => "0000000111000000000000101000000100",
			4270 => "00000010010011000100010000011101",
			4271 => "11111110001101110100010000011101",
			4272 => "0000001011000000001000111100001100",
			4273 => "0000000011000000001101111000001000",
			4274 => "0000000011000000001001110000000100",
			4275 => "00000010001111100100010000011101",
			4276 => "11111111111110100100010000011101",
			4277 => "00000010010001100100010000011101",
			4278 => "0000000111000000000100000000000100",
			4279 => "00000000100101010100010000011101",
			4280 => "11111110001001110100010000011101",
			4281 => "0000000010000000000110100000011000",
			4282 => "0000000011000000000100000000001000",
			4283 => "0000001101000000000110000100000100",
			4284 => "11111110010011000100010000011101",
			4285 => "00000000000000000100010000011101",
			4286 => "0000001010000000000011101000001000",
			4287 => "0000000011000000001010011100000100",
			4288 => "11111110001101100100010000011101",
			4289 => "00000000100000000100010000011101",
			4290 => "0000001100000000000000101000000100",
			4291 => "00000000111100110100010000011101",
			4292 => "00000010011000100100010000011101",
			4293 => "0000000010000000001100100100010000",
			4294 => "0000000010000000001110101000001000",
			4295 => "0000000010000000001110101000000100",
			4296 => "11111111100100100100010000011101",
			4297 => "00000001011010010100010000011101",
			4298 => "0000001010000000001000100100000100",
			4299 => "00000000000000000100010000011101",
			4300 => "11111101100001100100010000011101",
			4301 => "0000001101000000000000001100001000",
			4302 => "0000000001000000001100110100000100",
			4303 => "11111111110110100100010000011101",
			4304 => "00000001000001010100010000011101",
			4305 => "0000000101000000000000001100000100",
			4306 => "11111110100110010100010000011101",
			4307 => "00000000000101100100010000011101",
			4308 => "0000001010000000000110011000011000",
			4309 => "0000001100000000000100010100000100",
			4310 => "11111110101010100100010000011101",
			4311 => "0000001101000000001100101100000100",
			4312 => "00000011111001100100010000011101",
			4313 => "0000000100000000001101001000001100",
			4314 => "0000000110000000000100110100000100",
			4315 => "00000000011110010100010000011101",
			4316 => "0000000000000000001111000100000100",
			4317 => "00000000000000000100010000011101",
			4318 => "00000010011001010100010000011101",
			4319 => "11111110001001100100010000011101",
			4320 => "0000001100000000000000111000011000",
			4321 => "0000000010000000000110100000000100",
			4322 => "11111110110011010100010000011101",
			4323 => "0000000110000000000001111000000100",
			4324 => "11111111010100110100010000011101",
			4325 => "0000001100000000000000111000001000",
			4326 => "0000000001000000001110011100000100",
			4327 => "00000000000000000100010000011101",
			4328 => "00000000101101100100010000011101",
			4329 => "0000000000000000001101111000000100",
			4330 => "00000010011011010100010000011101",
			4331 => "00000000000000000100010000011101",
			4332 => "0000000011000000001011000100011100",
			4333 => "0000000100000000000100001100010000",
			4334 => "0000001100000000001010000000001000",
			4335 => "0000001100000000001010000000000100",
			4336 => "11111110101010110100010000011101",
			4337 => "00000001000011000100010000011101",
			4338 => "0000001010000000001010110000000100",
			4339 => "11111110100101110100010000011101",
			4340 => "11111111111100000100010000011101",
			4341 => "0000000000000000000100010100000100",
			4342 => "00000001111011100100010000011101",
			4343 => "0000000100000000001111100000000100",
			4344 => "11111110010011000100010000011101",
			4345 => "00000000001001010100010000011101",
			4346 => "0000001000000000001001101000001100",
			4347 => "0000000100000000001011110000001000",
			4348 => "0000000101000000001000000000000100",
			4349 => "00000000000000000100010000011101",
			4350 => "00000001010011100100010000011101",
			4351 => "11111101001110010100010000011101",
			4352 => "0000000010000000001110000100001000",
			4353 => "0000000010000000001110000100000100",
			4354 => "00000000011000010100010000011101",
			4355 => "00000010000110110100010000011101",
			4356 => "0000000100000000000101010100000100",
			4357 => "00000000010000110100010000011101",
			4358 => "00000000000011000100010000011101",
			4359 => "0000001011000000000110000110111100",
			4360 => "0000000100000000000100001101100000",
			4361 => "0000001110000000000111111000100100",
			4362 => "0000000100000000000110101100000100",
			4363 => "11100111111100100100011001100001",
			4364 => "0000000110000000001101111100010000",
			4365 => "0000000110000000000111101000001000",
			4366 => "0000001011000000000100010100000100",
			4367 => "11100000111110110100011001100001",
			4368 => "11011110011100110100011001100001",
			4369 => "0000000011000000000100010100000100",
			4370 => "11011111000100110100011001100001",
			4371 => "11100000101100000100011001100001",
			4372 => "0000000000000000000000111000001000",
			4373 => "0000001001000000001001111000000100",
			4374 => "11101010001010010100011001100001",
			4375 => "11100011010101000100011001100001",
			4376 => "0000000101000000000110000100000100",
			4377 => "11100001010010100100011001100001",
			4378 => "11011110010100110100011001100001",
			4379 => "0000000110000000000111101000011100",
			4380 => "0000001000000000000001010100010000",
			4381 => "0000001010000000000011101000001000",
			4382 => "0000000110000000001011111100000100",
			4383 => "11011110000011000100011001100001",
			4384 => "11011110111100010100011001100001",
			4385 => "0000000100000000000110111000000100",
			4386 => "11100011100111100100011001100001",
			4387 => "11011110101001110100011001100001",
			4388 => "0000001001000000000110101000001000",
			4389 => "0000000100000000001100001100000100",
			4390 => "11101000000010100100011001100001",
			4391 => "11100000001100100100011001100001",
			4392 => "11011110001010000100011001100001",
			4393 => "0000000100000000001101001000010000",
			4394 => "0000000110000000001101111100001000",
			4395 => "0000000010000000001100100100000100",
			4396 => "11100111011100000100011001100001",
			4397 => "11100011101100110100011001100001",
			4398 => "0000000111000000001001110000000100",
			4399 => "11101000000110100100011001100001",
			4400 => "11100010011000110100011001100001",
			4401 => "0000000111000000000000101000001000",
			4402 => "0000000110000000001100011000000100",
			4403 => "11100101010000110100011001100001",
			4404 => "11101001010011100100011001100001",
			4405 => "0000001110000000000110000100000100",
			4406 => "11100010010111100100011001100001",
			4407 => "11100100011110000100011001100001",
			4408 => "0000000110000000001101111100011100",
			4409 => "0000000100000000000011110100001100",
			4410 => "0000000000000000001010000000000100",
			4411 => "11011110001001010100011001100001",
			4412 => "0000000000000000000100010100000100",
			4413 => "11100101100111100100011001100001",
			4414 => "11100000011000100100011001100001",
			4415 => "0000000001000000000000011000000100",
			4416 => "11011110000001110100011001100001",
			4417 => "0000000100000000000011101100000100",
			4418 => "11011110001100000100011001100001",
			4419 => "0000001001000000000010001100000100",
			4420 => "11100000001100100100011001100001",
			4421 => "11011110001111000100011001100001",
			4422 => "0000001001000000001001111000100000",
			4423 => "0000000000000000001011000100010000",
			4424 => "0000000011000000001001110000001000",
			4425 => "0000000100000000001111100000000100",
			4426 => "11100001010101100100011001100001",
			4427 => "11100100011001100100011001100001",
			4428 => "0000000111000000001011000100000100",
			4429 => "11101000110111010100011001100001",
			4430 => "11100100001100110100011001100001",
			4431 => "0000000100000000001011100000001000",
			4432 => "0000000011000000001100001000000100",
			4433 => "11011110110001100100011001100001",
			4434 => "11100001000111000100011001100001",
			4435 => "0000000100000000000011111000000100",
			4436 => "11100010001101010100011001100001",
			4437 => "11011110000101110100011001100001",
			4438 => "0000001110000000000110000100010000",
			4439 => "0000000101000000000110000100001000",
			4440 => "0000000000000000000100010100000100",
			4441 => "11100010001111100100011001100001",
			4442 => "11011111100101000100011001100001",
			4443 => "0000000010000000001111010000000100",
			4444 => "11100010000010100100011001100001",
			4445 => "11011110111010010100011001100001",
			4446 => "0000000100000000000011010100001000",
			4447 => "0000001000000000000001110100000100",
			4448 => "11011111111000000100011001100001",
			4449 => "11100111110101000100011001100001",
			4450 => "0000001111000000001001010000000100",
			4451 => "11011111111110110100011001100001",
			4452 => "11100011001000110100011001100001",
			4453 => "0000000111000000000101101100111100",
			4454 => "0000000110000000001001100100101000",
			4455 => "0000000011000000000001101000010000",
			4456 => "0000000101000000001010111000000100",
			4457 => "11100001101110100100011001100001",
			4458 => "0000000011000000001000000000000100",
			4459 => "11011110000010100100011001100001",
			4460 => "0000000111000000001101100000000100",
			4461 => "11100001111100010100011001100001",
			4462 => "11011110001000010100011001100001",
			4463 => "0000001010000000001000010100001000",
			4464 => "0000000110000000001101111100000100",
			4465 => "11100011010000000100011001100001",
			4466 => "11101001000011000100011001100001",
			4467 => "0000001001000000000101011100001000",
			4468 => "0000001011000000001101111000000100",
			4469 => "11100001010101010100011001100001",
			4470 => "11100101101110110100011001100001",
			4471 => "0000000000000000000010111100000100",
			4472 => "11011110001111000100011001100001",
			4473 => "11011111100011100100011001100001",
			4474 => "0000000110000000001001100100010000",
			4475 => "0000000111000000001001110000000100",
			4476 => "11100001100101100100011001100001",
			4477 => "0000001111000000001001011100000100",
			4478 => "11011110000100110100011001100001",
			4479 => "0000000001000000000111100100000100",
			4480 => "11011110001111000100011001100001",
			4481 => "11100000100111000100011001100001",
			4482 => "11011110000010100100011001100001",
			4483 => "0000000111000000001101111000011100",
			4484 => "0000001110000000001001001000001100",
			4485 => "0000001011000000001110001100001000",
			4486 => "0000000101000000000011100000000100",
			4487 => "11011110001100110100011001100001",
			4488 => "11011111011011000100011001100001",
			4489 => "11011110000010000100011001100001",
			4490 => "0000000010000000000111010100001100",
			4491 => "0000000000000000001011010100000100",
			4492 => "11011110000100010100011001100001",
			4493 => "0000001011000000000100001000000100",
			4494 => "11011111100110010100011001100001",
			4495 => "11101000001110110100011001100001",
			4496 => "11011110000011100100011001100001",
			4497 => "0000001000000000000110011100001100",
			4498 => "0000001010000000000010101100000100",
			4499 => "11011110000001110100011001100001",
			4500 => "0000001000000000001100011100000100",
			4501 => "11011110001011100100011001100001",
			4502 => "11011110011010000100011001100001",
			4503 => "11011110000001110100011001100001",
			4504 => "0000001000000000001001101010101000",
			4505 => "0000001000000000001001101001100100",
			4506 => "0000001101000000000101101100101100",
			4507 => "0000000111000000000100010100011100",
			4508 => "0000001100000000000111111000010000",
			4509 => "0000000011000000001011000100001000",
			4510 => "0000000111000000001110111100000100",
			4511 => "00000000000000000100100010110101",
			4512 => "00000010110111110100100010110101",
			4513 => "0000000011000000001000111000000100",
			4514 => "11111111010001100100100010110101",
			4515 => "00000001111000010100100010110101",
			4516 => "0000001101000000001100110000001000",
			4517 => "0000001001000000000010001100000100",
			4518 => "00000000000000000100100010110101",
			4519 => "11111110001001100100100010110101",
			4520 => "00000000011101010100100010110101",
			4521 => "0000000010000000001101000100001100",
			4522 => "0000000011000000000100010100000100",
			4523 => "00000000000010110100100010110101",
			4524 => "0000001110000000000000110000000100",
			4525 => "00000011011111100100100010110101",
			4526 => "00000001001101110100100010110101",
			4527 => "11111111011101010100100010110101",
			4528 => "0000001110000000001000111100011000",
			4529 => "0000000111000000000100010100001000",
			4530 => "0000000001000000001110100000000100",
			4531 => "11111111010110010100100010110101",
			4532 => "00000010110110110100100010110101",
			4533 => "0000001011000000000000101000001000",
			4534 => "0000000000000000000010111100000100",
			4535 => "11111110000110010100100010110101",
			4536 => "11111111100000010100100010110101",
			4537 => "0000001011000000001100001000000100",
			4538 => "00000000100101100100100010110101",
			4539 => "11111111011011010100100010110101",
			4540 => "0000000111000000000000101000010000",
			4541 => "0000000010000000000101001000001000",
			4542 => "0000000101000000001100101100000100",
			4543 => "00000000000000000100100010110101",
			4544 => "00000001011100100100100010110101",
			4545 => "0000000100000000000110001100000100",
			4546 => "00000010000001000100100010110101",
			4547 => "00000011000110010100100010110101",
			4548 => "0000000100000000000110001100001000",
			4549 => "0000000000000000001111000100000100",
			4550 => "11111111110100010100100010110101",
			4551 => "00000000110010000100100010110101",
			4552 => "0000001101000000000001111100000100",
			4553 => "11111111101001100100100010110101",
			4554 => "11111101001101100100100010110101",
			4555 => "0000000010000000000101110000100100",
			4556 => "0000001010000000001000010100010000",
			4557 => "0000000000000000000011111100001100",
			4558 => "0000001010000000001000010100000100",
			4559 => "00000000000000000100100010110101",
			4560 => "0000001011000000001100001000000100",
			4561 => "11111101110000110100100010110101",
			4562 => "11111111000111000100100010110101",
			4563 => "00000000010111010100100010110101",
			4564 => "0000000000000000001111000100000100",
			4565 => "11111101011000010100100010110101",
			4566 => "0000000011000000000110000100001000",
			4567 => "0000000010000000000111100000000100",
			4568 => "00000000100010100100100010110101",
			4569 => "11111110111000010100100010110101",
			4570 => "0000001100000000000000101000000100",
			4571 => "00000010000001000100100010110101",
			4572 => "00000000000100100100100010110101",
			4573 => "0000000001000000001001111000010000",
			4574 => "0000001110000000001010111100001100",
			4575 => "0000001110000000001101111000001000",
			4576 => "0000000010000000001100010100000100",
			4577 => "11111110011011100100100010110101",
			4578 => "00000001111101000100100010110101",
			4579 => "00000001111011110100100010110101",
			4580 => "11111100011010010100100010110101",
			4581 => "0000001010000000000110011000001100",
			4582 => "0000000010000000000010000100001000",
			4583 => "0000001110000000001010111000000100",
			4584 => "11111110111110100100100010110101",
			4585 => "00000001011000000100100010110101",
			4586 => "11111101110010010100100010110101",
			4587 => "11111101011111000100100010110101",
			4588 => "0000001000000000001011010100101100",
			4589 => "0000000010000000001110010000011100",
			4590 => "0000001100000000001010000000000100",
			4591 => "00000010110101100100100010110101",
			4592 => "0000001010000000001001000100001000",
			4593 => "0000001010000000001001000100000100",
			4594 => "00000000000010100100100010110101",
			4595 => "11111110001111000100100010110101",
			4596 => "0000000101000000001100101100001000",
			4597 => "0000000001000000001100110100000100",
			4598 => "00000001001011010100100010110101",
			4599 => "11111110101110000100100010110101",
			4600 => "0000001101000000000100001000000100",
			4601 => "00000010001101110100100010110101",
			4602 => "00000001000101110100100010110101",
			4603 => "0000000010000000001110110100001000",
			4604 => "0000000001000000001001111000000100",
			4605 => "11111111111101000100100010110101",
			4606 => "11111100110010110100100010110101",
			4607 => "0000000111000000000110000100000100",
			4608 => "00000001111101110100100010110101",
			4609 => "11111111110000010100100010110101",
			4610 => "0000001000000000001011010100011000",
			4611 => "0000000000000000000011010000010100",
			4612 => "0000000100000000000010111000001100",
			4613 => "0000001110000000000000101000000100",
			4614 => "00000001000110100100100010110101",
			4615 => "0000001110000000001110001100000100",
			4616 => "11111101111011000100100010110101",
			4617 => "00000000000100100100100010110101",
			4618 => "0000000000000000000011111100000100",
			4619 => "00000000000000000100100010110101",
			4620 => "00000011111100110100100010110101",
			4621 => "11111101110010010100100010110101",
			4622 => "0000000000000000000000111000100000",
			4623 => "0000001000000000001011010100010000",
			4624 => "0000001010000000000110011000001000",
			4625 => "0000000001000000001100110100000100",
			4626 => "11111111101011110100100010110101",
			4627 => "11111101001010000100100010110101",
			4628 => "0000000100000000000011001100000100",
			4629 => "00000001010110100100100010110101",
			4630 => "11111111001111110100100010110101",
			4631 => "0000000010000000001001011100001000",
			4632 => "0000000100000000000110001100000100",
			4633 => "11111111101001010100100010110101",
			4634 => "00000001000100100100100010110101",
			4635 => "0000000100000000000010111000000100",
			4636 => "00000000100000000100100010110101",
			4637 => "11111111000010110100100010110101",
			4638 => "0000000101000000000110000100010000",
			4639 => "0000000001000000001100110100001000",
			4640 => "0000001001000000000111100100000100",
			4641 => "00000000001011110100100010110101",
			4642 => "11111110100000100100100010110101",
			4643 => "0000001100000000000100010100000100",
			4644 => "00000001111001100100100010110101",
			4645 => "00000000000000000100100010110101",
			4646 => "0000000100000000000100001100001000",
			4647 => "0000001110000000001000111000000100",
			4648 => "11111111101111110100100010110101",
			4649 => "00000000001100100100100010110101",
			4650 => "0000001000000000001111001000000100",
			4651 => "00000100010110100100100010110101",
			4652 => "11111111010111100100100010110101",
			4653 => "0000001100000000000110000111001100",
			4654 => "0000001010000000000001010001100000",
			4655 => "0000000010000000001110101000101100",
			4656 => "0000000010000000001110101000100000",
			4657 => "0000001010000000000011101000010000",
			4658 => "0000001011000000001011000100001000",
			4659 => "0000001111000000000110100100000100",
			4660 => "00000010010110000100101001101001",
			4661 => "11111110111001110100101001101001",
			4662 => "0000001111000000000100010000000100",
			4663 => "11111110100010000100101001101001",
			4664 => "00000000100000100100101001101001",
			4665 => "0000000010000000000000110100001000",
			4666 => "0000001000000000000001010100000100",
			4667 => "00000010000100000100101001101001",
			4668 => "11111111000100000100101001101001",
			4669 => "0000001111000000000110100100000100",
			4670 => "00000001110111000100101001101001",
			4671 => "00000000100100000100101001101001",
			4672 => "0000000101000000001101100000000100",
			4673 => "11111111100101110100101001101001",
			4674 => "0000001101000000000110000100000100",
			4675 => "00000011110111100100101001101001",
			4676 => "00000001110110100100101001101001",
			4677 => "0000000101000000000100011000011100",
			4678 => "0000000010000000001110010000010000",
			4679 => "0000001110000000001100001000001000",
			4680 => "0000001001000000000110101000000100",
			4681 => "00000000000011110100101001101001",
			4682 => "11111111011011000100101001101001",
			4683 => "0000001000000000001001101000000100",
			4684 => "11111111111010100100101001101001",
			4685 => "00000000100010000100101001101001",
			4686 => "0000001100000000001000111000001000",
			4687 => "0000000000000000000000111000000100",
			4688 => "11111111001011110100101001101001",
			4689 => "11111111110101110100101001101001",
			4690 => "00000001111110100100101001101001",
			4691 => "0000001110000000000001101000001100",
			4692 => "0000001100000000001001110000001000",
			4693 => "0000000011000000001000011000000100",
			4694 => "00000001010101000100101001101001",
			4695 => "00000100000000010100101001101001",
			4696 => "00000000010111110100101001101001",
			4697 => "0000000001000000000110101000000100",
			4698 => "11111110001110110100101001101001",
			4699 => "0000000000000000000001110100000100",
			4700 => "00000010000001110100101001101001",
			4701 => "00000000001101100100101001101001",
			4702 => "0000000100000000001001001101000000",
			4703 => "0000001001000000001011101000100000",
			4704 => "0000000010000000001110010000010000",
			4705 => "0000001001000000000110101000001000",
			4706 => "0000000000000000001110111100000100",
			4707 => "00000010100110010100101001101001",
			4708 => "00000000100110000100101001101001",
			4709 => "0000000000000000000000111000000100",
			4710 => "00000010000101010100101001101001",
			4711 => "11111111101100010100101001101001",
			4712 => "0000001011000000001001110000001000",
			4713 => "0000001001000000001101101000000100",
			4714 => "00000001011000100100101001101001",
			4715 => "11111111101011110100101001101001",
			4716 => "0000001000000000001111001000000100",
			4717 => "00000000011110010100101001101001",
			4718 => "00000010100010000100101001101001",
			4719 => "0000000010000000001100010000010000",
			4720 => "0000000000000000000000111000001000",
			4721 => "0000001101000000000011100000000100",
			4722 => "00000001011110000100101001101001",
			4723 => "11111111001000010100101001101001",
			4724 => "0000000011000000001001001000000100",
			4725 => "11111110000110110100101001101001",
			4726 => "11111111110101110100101001101001",
			4727 => "0000001011000000000110000100001000",
			4728 => "0000000101000000000111001000000100",
			4729 => "00000000100110100100101001101001",
			4730 => "00000010100111010100101001101001",
			4731 => "0000001010000000001010110000000100",
			4732 => "00000010110001000100101001101001",
			4733 => "11111111001000000100101001101001",
			4734 => "0000000011000000000011111100001100",
			4735 => "0000000000000000000011011100000100",
			4736 => "11111110001000010100101001101001",
			4737 => "0000000100000000000011111000000100",
			4738 => "00000000101010110100101001101001",
			4739 => "11111110011101100100101001101001",
			4740 => "0000001111000000000100000100010000",
			4741 => "0000000011000000001000111100001000",
			4742 => "0000001001000000001001111000000100",
			4743 => "00000000101100000100101001101001",
			4744 => "11111110010000010100101001101001",
			4745 => "0000000001000000001100110100000100",
			4746 => "00000101001001010100101001101001",
			4747 => "00000011000011100100101001101001",
			4748 => "0000001100000000001110111100001000",
			4749 => "0000001100000000001010000000000100",
			4750 => "00000000000100110100101001101001",
			4751 => "00000010000100000100101001101001",
			4752 => "0000000011000000001100001000000100",
			4753 => "11111110110100010100101001101001",
			4754 => "00000000000111100100101001101001",
			4755 => "0000001100000000001010111100001100",
			4756 => "0000000000000000000111000100001000",
			4757 => "0000000000000000001111001000000100",
			4758 => "11111110101111000100101001101001",
			4759 => "00000010010100010100101001101001",
			4760 => "11111110011101110100101001101001",
			4761 => "11111110011010000100101001101001",
			4762 => "0000001111000000000010001010000100",
			4763 => "0000000011000000000110000101011000",
			4764 => "0000001101000000001101111000110100",
			4765 => "0000000101000000001110001100100000",
			4766 => "0000001011000000000100000000010000",
			4767 => "0000000001000000001100110100001000",
			4768 => "0000000101000000001100101100000100",
			4769 => "00000000000100110100110011000101",
			4770 => "11111111000001110100110011000101",
			4771 => "0000001001000000000111100100000100",
			4772 => "00000000111010100100110011000101",
			4773 => "11111110110000000100110011000101",
			4774 => "0000000100000000000101000000001000",
			4775 => "0000000001000000001110100000000100",
			4776 => "11111110110100000100110011000101",
			4777 => "00000001010101100100110011000101",
			4778 => "0000000001000000001110100000000100",
			4779 => "00000000000000000100110011000101",
			4780 => "11111110100001010100110011000101",
			4781 => "0000000100000000001000000100000100",
			4782 => "11111101111101010100110011000101",
			4783 => "0000000100000000001010110100001000",
			4784 => "0000000100000000000011001100000100",
			4785 => "00000000100110100100110011000101",
			4786 => "00000010011110000100110011000101",
			4787 => "0000000100000000001110111000000100",
			4788 => "11111110010110000100110011000101",
			4789 => "00000000111010000100110011000101",
			4790 => "0000001111000000001011011100011100",
			4791 => "0000001101000000001100101000010000",
			4792 => "0000000011000000001100110000001000",
			4793 => "0000000111000000001100001000000100",
			4794 => "00000000001010110100110011000101",
			4795 => "11111110010010110100110011000101",
			4796 => "0000000110000000001101111100000100",
			4797 => "11111111100111110100110011000101",
			4798 => "00000001100011000100110011000101",
			4799 => "0000001011000000001001110000000100",
			4800 => "11111110010010000100110011000101",
			4801 => "0000000110000000000100110100000100",
			4802 => "11111111111100000100110011000101",
			4803 => "00000000111100010100110011000101",
			4804 => "0000000001000000001110100000000100",
			4805 => "00000000000000000100110011000101",
			4806 => "11111101101011010100110011000101",
			4807 => "0000000111000000001100001000010000",
			4808 => "0000000111000000000100010100000100",
			4809 => "11111110101100000100110011000101",
			4810 => "0000000110000000000001111000000100",
			4811 => "00000000011101100100110011000101",
			4812 => "0000001110000000001000111100000100",
			4813 => "00000010111011100100110011000101",
			4814 => "00000001101010000100110011000101",
			4815 => "0000001001000000000111100100001100",
			4816 => "0000001111000000000101100100000100",
			4817 => "11111110100010000100110011000101",
			4818 => "0000000011000000001100101100000100",
			4819 => "00000010010111110100110011000101",
			4820 => "00000001000010110100110011000101",
			4821 => "0000001011000000001100001000000100",
			4822 => "11111101110111010100110011000101",
			4823 => "0000000011000000000110000100000100",
			4824 => "00000010011011010100110011000101",
			4825 => "0000000110000000001101111100000100",
			4826 => "00000000010110010100110011000101",
			4827 => "11111110111010100100110011000101",
			4828 => "0000000011000000001100101100110100",
			4829 => "0000000011000000001100101100101000",
			4830 => "0000000101000000001101111000100000",
			4831 => "0000000101000000001100101100010000",
			4832 => "0000001011000000000100000000001000",
			4833 => "0000001101000000001110001100000100",
			4834 => "11111111111000110100110011000101",
			4835 => "11111110100100110100110011000101",
			4836 => "0000000111000000001100001000000100",
			4837 => "11111111111011010100110011000101",
			4838 => "00000010110101010100110011000101",
			4839 => "0000000001000000001100110100001000",
			4840 => "0000001110000000000000101000000100",
			4841 => "11111101111000100100110011000101",
			4842 => "11111111000111100100110011000101",
			4843 => "0000000111000000000100000000000100",
			4844 => "00000001110001000100110011000101",
			4845 => "11111110010110000100110011000101",
			4846 => "0000000111000000000100000000000100",
			4847 => "00000010110110100100110011000101",
			4848 => "11111111011111000100110011000101",
			4849 => "0000001001000000000111100100001000",
			4850 => "0000001101000000000110000100000100",
			4851 => "00000000000000000100110011000101",
			4852 => "11111101111011010100110011000101",
			4853 => "11111111111110010100110011000101",
			4854 => "0000000100000000000101010100111000",
			4855 => "0000000001000000001100110100100000",
			4856 => "0000000000000000000011111100010000",
			4857 => "0000000110000000000001111000001000",
			4858 => "0000001101000000001101111000000100",
			4859 => "00000001100001010100110011000101",
			4860 => "11111111011101010100110011000101",
			4861 => "0000000011000000001101111000000100",
			4862 => "00000000010010000100110011000101",
			4863 => "11111111010010010100110011000101",
			4864 => "0000000001000000001100110100001000",
			4865 => "0000001011000000000000101000000100",
			4866 => "00000001101011100100110011000101",
			4867 => "11111111100011100100110011000101",
			4868 => "0000001011000000001100001000000100",
			4869 => "00000000001010100100110011000101",
			4870 => "00000001001001010100110011000101",
			4871 => "0000001011000000000100000000001100",
			4872 => "0000000011000000001010111000001000",
			4873 => "0000001101000000001101111000000100",
			4874 => "11111111101001100100110011000101",
			4875 => "11111101111001100100110011000101",
			4876 => "00000001000011110100110011000101",
			4877 => "0000001101000000001101111000000100",
			4878 => "00000010101110000100110011000101",
			4879 => "0000000000000000001110111100000100",
			4880 => "00000000000011010100110011000101",
			4881 => "11111110100000110100110011000101",
			4882 => "0000001000000000000111000100100000",
			4883 => "0000001011000000001000111100010000",
			4884 => "0000000001000000001100110100001000",
			4885 => "0000001101000000000101101100000100",
			4886 => "00000001010010100100110011000101",
			4887 => "11111110001001100100110011000101",
			4888 => "0000001101000000001101111000000100",
			4889 => "00000001000111110100110011000101",
			4890 => "11111111110110000100110011000101",
			4891 => "0000001010000000000001010000001000",
			4892 => "0000001000000000001011010100000100",
			4893 => "11111111110010110100110011000101",
			4894 => "00000001000010010100110011000101",
			4895 => "0000000000000000000000110000000100",
			4896 => "11111110001011100100110011000101",
			4897 => "11111111000111010100110011000101",
			4898 => "0000000100000000000100001100010000",
			4899 => "0000000110000000001101011000001000",
			4900 => "0000000111000000001000111100000100",
			4901 => "00000000001010000100110011000101",
			4902 => "00000000111101110100110011000101",
			4903 => "0000001111000000001101000100000100",
			4904 => "11111110010100100100110011000101",
			4905 => "11111111111001100100110011000101",
			4906 => "0000001010000000000110011100001000",
			4907 => "0000000101000000000110000100000100",
			4908 => "00000000100101010100110011000101",
			4909 => "11111110111010110100110011000101",
			4910 => "0000001111000000000001001000000100",
			4911 => "00000001100011110100110011000101",
			4912 => "00000000000110000100110011000101",
			4913 => "0000001010000000000110011010101100",
			4914 => "0000001000000000001001101001011000",
			4915 => "0000001000000000001100000100110000",
			4916 => "0000000100000000001000011100010100",
			4917 => "0000000000000000000010011000010000",
			4918 => "0000000100000000001000110100001000",
			4919 => "0000000100000000001110000000000100",
			4920 => "00000000001111100100111100101001",
			4921 => "11111111100100010100111100101001",
			4922 => "0000001011000000001000111100000100",
			4923 => "00000001111111000100111100101001",
			4924 => "11111111101011100100111100101001",
			4925 => "11111110001110100100111100101001",
			4926 => "0000001010000000001000010100010000",
			4927 => "0000001010000000001000100100001000",
			4928 => "0000001110000000000100000000000100",
			4929 => "11111111000110000100111100101001",
			4930 => "00000000100111100100111100101001",
			4931 => "0000000100000000000010110000000100",
			4932 => "11111110001001100100111100101001",
			4933 => "00000000100101000100111100101001",
			4934 => "0000001010000000001000010100001000",
			4935 => "0000000000000000001101010000000100",
			4936 => "00000000000000000100111100101001",
			4937 => "00000010000000000100111100101001",
			4938 => "11111110010011010100111100101001",
			4939 => "0000000100000000000110111000001000",
			4940 => "0000001101000000001110110000000100",
			4941 => "11111101111011010100111100101001",
			4942 => "00000000000000000100111100101001",
			4943 => "0000000100000000000011110000010000",
			4944 => "0000000000000000000010111100001000",
			4945 => "0000000000000000000010111100000100",
			4946 => "00000000111100010100111100101001",
			4947 => "11111111001110000100111100101001",
			4948 => "0000001110000000000100010100000100",
			4949 => "00000000011100010100111100101001",
			4950 => "00000010011010110100111100101001",
			4951 => "0000000111000000001011000100001000",
			4952 => "0000000011000000001000111000000100",
			4953 => "11111111000100010100111100101001",
			4954 => "00000010001001010100111100101001",
			4955 => "0000001011000000001100001000000100",
			4956 => "00000000001110110100111100101001",
			4957 => "11111110101011000100111100101001",
			4958 => "0000001010000000001001000100100000",
			4959 => "0000001100000000000111111000001100",
			4960 => "0000000000000000000011111100000100",
			4961 => "11111110001100010100111100101001",
			4962 => "0000000101000000000011011100000100",
			4963 => "11111111000011000100111100101001",
			4964 => "00000001101111100100111100101001",
			4965 => "0000000111000000001100001000010000",
			4966 => "0000001001000000000110101000001000",
			4967 => "0000001001000000001001111000000100",
			4968 => "11111110001100000100111100101001",
			4969 => "00000000000000000100111100101001",
			4970 => "0000001100000000000100010100000100",
			4971 => "11111110010010010100111100101001",
			4972 => "11111101000110110100111100101001",
			4973 => "11111111111010000100111100101001",
			4974 => "0000001101000000000000001100011000",
			4975 => "0000000000000000000011010000001100",
			4976 => "0000000100000000001000110100000100",
			4977 => "11111110010000010100111100101001",
			4978 => "0000000100000000000101000000000100",
			4979 => "00000001110110010100111100101001",
			4980 => "00000000010010000100111100101001",
			4981 => "0000000100000000001000001000000100",
			4982 => "11111101100110110100111100101001",
			4983 => "0000001100000000000100010100000100",
			4984 => "11111111100000010100111100101001",
			4985 => "00000001010101000100111100101001",
			4986 => "0000000101000000000000001100001100",
			4987 => "0000000111000000001011000100000100",
			4988 => "00000000010011110100111100101001",
			4989 => "0000000111000000001100001000000100",
			4990 => "11111100001011010100111100101001",
			4991 => "11111110011111000100111100101001",
			4992 => "0000000101000000001101010100001000",
			4993 => "0000000001000000000010001100000100",
			4994 => "11111111111011010100111100101001",
			4995 => "00000001001110010100111100101001",
			4996 => "0000000100000000000011110000000100",
			4997 => "00000000000011100100111100101001",
			4998 => "11111101110110000100111100101001",
			4999 => "0000000100000000001000001001001100",
			5000 => "0000000000000000000010111100011000",
			5001 => "0000000010000000000100101000000100",
			5002 => "11111101100011100100111100101001",
			5003 => "0000000100000000000011110000010000",
			5004 => "0000000100000000001110100100001000",
			5005 => "0000000011000000001001110100000100",
			5006 => "11111110010011100100111100101001",
			5007 => "00000000000000000100111100101001",
			5008 => "0000001001000000000000111100000100",
			5009 => "00000001110000100100111100101001",
			5010 => "11111110100100010100111100101001",
			5011 => "11111101011000100100111100101001",
			5012 => "0000000000000000000000111000011100",
			5013 => "0000001101000000001010111000010000",
			5014 => "0000001010000000000001010000001000",
			5015 => "0000000100000000000010110000000100",
			5016 => "00000001000010010100111100101001",
			5017 => "11111111110001110100111100101001",
			5018 => "0000000100000000000110001100000100",
			5019 => "00000001000001000100111100101001",
			5020 => "00000001111110000100111100101001",
			5021 => "0000000101000000001101010100000100",
			5022 => "11111110100111010100111100101001",
			5023 => "0000001100000000001000111100000100",
			5024 => "00000001010100010100111100101001",
			5025 => "11111111110010100100111100101001",
			5026 => "0000000010000000000100101000001000",
			5027 => "0000001010000000000001010000000100",
			5028 => "11111101100000000100111100101001",
			5029 => "11111111011100110100111100101001",
			5030 => "0000000111000000001000111000001000",
			5031 => "0000001000000000001111001000000100",
			5032 => "00000001110100000100111100101001",
			5033 => "00000000000000000100111100101001",
			5034 => "0000000000000000000000111000000100",
			5035 => "11111111100101100100111100101001",
			5036 => "11111110001110010100111100101001",
			5037 => "0000000000000000000011111100001000",
			5038 => "0000001000000000001011010100000100",
			5039 => "11111110101100010100111100101001",
			5040 => "11111101101101110100111100101001",
			5041 => "0000001011000000001100101100100000",
			5042 => "0000001001000000001101101000010000",
			5043 => "0000001011000000000011011100001000",
			5044 => "0000001110000000000110000100000100",
			5045 => "00000000000011000100111100101001",
			5046 => "00000000100011110100111100101001",
			5047 => "0000000011000000000111001000000100",
			5048 => "00000010001111100100111100101001",
			5049 => "11111111111011010100111100101001",
			5050 => "0000001110000000001100101100001000",
			5051 => "0000000000000000000000110000000100",
			5052 => "11111111110010010100111100101001",
			5053 => "11111110101000110100111100101001",
			5054 => "0000001100000000000000101000000100",
			5055 => "11111111010010000100111100101001",
			5056 => "00000000001101000100111100101001",
			5057 => "0000000010000000001000001100010000",
			5058 => "0000001100000000000011011100001000",
			5059 => "0000001110000000000111001000000100",
			5060 => "00000011100011000100111100101001",
			5061 => "00000001000111100100111100101001",
			5062 => "0000001001000000001001011000000100",
			5063 => "11111111000110100100111100101001",
			5064 => "00000001010111100100111100101001",
			5065 => "11111110100100000100111100101001",
			5066 => "0000001001000000001101101011000100",
			5067 => "0000000111000000001100001001011000",
			5068 => "0000000111000000001100001001000000",
			5069 => "0000000111000000000000101000100000",
			5070 => "0000000111000000000000101000010000",
			5071 => "0000000111000000000000101000001000",
			5072 => "0000001100000000000000101000000100",
			5073 => "00000000000101010101000101100101",
			5074 => "00000001100001110101000101100101",
			5075 => "0000001000000000001010101100000100",
			5076 => "11111111010001000101000101100101",
			5077 => "00000001101011010101000101100101",
			5078 => "0000001001000000000110101000001000",
			5079 => "0000001011000000000000101000000100",
			5080 => "11111110001010010101000101100101",
			5081 => "00000000110110000101000101100101",
			5082 => "0000001110000000001110111100000100",
			5083 => "11111111100010100101000101100101",
			5084 => "11111101110001110101000101100101",
			5085 => "0000001001000000000111100100010000",
			5086 => "0000000001000000001100110100001000",
			5087 => "0000001011000000000000101000000100",
			5088 => "00000001001000000101000101100101",
			5089 => "00000000000010100101000101100101",
			5090 => "0000000010000000001001010000000100",
			5091 => "00000010000011010101000101100101",
			5092 => "00000000101001000101000101100101",
			5093 => "0000000111000000001100001000001000",
			5094 => "0000001000000000001001101000000100",
			5095 => "11111111100110000101000101100101",
			5096 => "00000000101000010101000101100101",
			5097 => "0000000000000000000011010000000100",
			5098 => "00000000101011100101000101100101",
			5099 => "11111111000111010101000101100101",
			5100 => "0000000001000000000010001100010100",
			5101 => "0000001111000000001101000100010000",
			5102 => "0000000110000000001100011000001000",
			5103 => "0000001100000000000100010100000100",
			5104 => "11111110011010110101000101100101",
			5105 => "11111111011101000101000101100101",
			5106 => "0000001100000000000100010100000100",
			5107 => "00000011010101100101000101100101",
			5108 => "11111111101011010101000101100101",
			5109 => "11111101001100010101000101100101",
			5110 => "11111100110111100101000101100101",
			5111 => "0000001110000000001000111000110000",
			5112 => "0000001011000000000100000000011000",
			5113 => "0000000111000000000100000000010000",
			5114 => "0000001110000000001010000000001000",
			5115 => "0000000010000000001100100100000100",
			5116 => "00000001101001100101000101100101",
			5117 => "11111110111011100101000101100101",
			5118 => "0000001111000000000101110100000100",
			5119 => "00000010110010110101000101100101",
			5120 => "00000000011001010101000101100101",
			5121 => "0000000110000000001100011000000100",
			5122 => "11111101001110100101000101100101",
			5123 => "11111111111010010101000101100101",
			5124 => "0000000011000000001100110000001000",
			5125 => "0000001000000000001001101000000100",
			5126 => "00000000000000000101000101100101",
			5127 => "11111110001101100101000101100101",
			5128 => "0000001111000000000001011000001000",
			5129 => "0000000011000000000110000100000100",
			5130 => "00000010100101010101000101100101",
			5131 => "00000000100101010101000101100101",
			5132 => "0000001001000000000111100100000100",
			5133 => "00000000000110110101000101100101",
			5134 => "11111110111110100101000101100101",
			5135 => "0000001001000000000111100100100000",
			5136 => "0000001000000000000111000100010000",
			5137 => "0000000111000000000100000000001000",
			5138 => "0000001110000000000011011100000100",
			5139 => "00000010010001100101000101100101",
			5140 => "00000000110100010101000101100101",
			5141 => "0000000111000000000100000000000100",
			5142 => "11111110010110010101000101100101",
			5143 => "00000001001100100101000101100101",
			5144 => "0000000100000000000100001100001000",
			5145 => "0000001100000000000000101000000100",
			5146 => "00000001111111010101000101100101",
			5147 => "00000011100010110101000101100101",
			5148 => "0000000011000000001010111100000100",
			5149 => "11111111010100000101000101100101",
			5150 => "00000010101100010101000101100101",
			5151 => "0000001100000000000100010100010000",
			5152 => "0000000110000000001100011000001000",
			5153 => "0000001111000000000101110100000100",
			5154 => "00000011000010110101000101100101",
			5155 => "00000000100111100101000101100101",
			5156 => "0000001111000000001110101100000100",
			5157 => "00000000111000010101000101100101",
			5158 => "00000011000010100101000101100101",
			5159 => "0000001100000000001011000100000100",
			5160 => "11111101100110000101000101100101",
			5161 => "0000000001000000001100110100000100",
			5162 => "11111111101001100101000101100101",
			5163 => "00000000101001100101000101100101",
			5164 => "0000001111000000000110110100010000",
			5165 => "0000001000000000001010110000001100",
			5166 => "0000000011000000001000000000000100",
			5167 => "11111110010011000101000101100101",
			5168 => "0000001110000000000111001000000100",
			5169 => "00000000000000000101000101100101",
			5170 => "11111111101101000101000101100101",
			5171 => "00000011011110100101000101100101",
			5172 => "0000000011000000000001111100010100",
			5173 => "0000000001000000000010001100000100",
			5174 => "11111111111001110101000101100101",
			5175 => "0000000010000000001001010000000100",
			5176 => "11111111100110010101000101100101",
			5177 => "0000000100000000001000001000000100",
			5178 => "11111100010101000101000101100101",
			5179 => "0000000111000000001000111000000100",
			5180 => "11111101110101110101000101100101",
			5181 => "11111110111010010101000101100101",
			5182 => "0000001100000000000100010100011000",
			5183 => "0000001100000000000100010100001000",
			5184 => "0000000010000000000110010000000100",
			5185 => "00000001110000100101000101100101",
			5186 => "11111111000000000101000101100101",
			5187 => "0000000111000000000100000000001000",
			5188 => "0000000111000000001100001000000100",
			5189 => "11111110101001010101000101100101",
			5190 => "00000001000111010101000101100101",
			5191 => "0000001011000000000011011100000100",
			5192 => "11111101000110010101000101100101",
			5193 => "11111111110000100101000101100101",
			5194 => "0000000111000000000100000000010000",
			5195 => "0000001110000000001100101000001000",
			5196 => "0000000011000000001010111000000100",
			5197 => "00000000010100010101000101100101",
			5198 => "11111110010011010101000101100101",
			5199 => "0000000110000000001100011000000100",
			5200 => "00000000010111100101000101100101",
			5201 => "00000001110111110101000101100101",
			5202 => "0000000110000000001101111100001000",
			5203 => "0000000010000000001001010000000100",
			5204 => "00000000000110000101000101100101",
			5205 => "11111110000000000101000101100101",
			5206 => "0000000100000000000011110000000100",
			5207 => "00000000010101010101000101100101",
			5208 => "11111111110010000101000101100101",
			5209 => "0000001100000000000110000111010000",
			5210 => "0000001010000000000001010001101100",
			5211 => "0000000010000000001110101000110000",
			5212 => "0000000010000000001101000100011100",
			5213 => "0000001010000000000011101000001100",
			5214 => "0000001011000000000100010100000100",
			5215 => "00000010010011110101001100100001",
			5216 => "0000000110000000000111101000000100",
			5217 => "11111110010101100101001100100001",
			5218 => "11111111111111010101001100100001",
			5219 => "0000000010000000000000110100001000",
			5220 => "0000001000000000000001010100000100",
			5221 => "00000010010010110101001100100001",
			5222 => "11111110111110010101001100100001",
			5223 => "0000000100000000001001001100000100",
			5224 => "00000000101011100101001100100001",
			5225 => "00000010111100010101001100100001",
			5226 => "0000001100000000000000101000010000",
			5227 => "0000001000000000001011010100001000",
			5228 => "0000000100000000001000001000000100",
			5229 => "00000010010011000101001100100001",
			5230 => "00000101010010000101001100100001",
			5231 => "0000000100000000000101010100000100",
			5232 => "11111111000110000101001100100001",
			5233 => "00000100001011010101001100100001",
			5234 => "11111111011011010101001100100001",
			5235 => "0000000110000000001100011000100000",
			5236 => "0000000010000000000011001000010000",
			5237 => "0000001010000000000001010000001000",
			5238 => "0000000110000000001101111100000100",
			5239 => "11111111101100100101001100100001",
			5240 => "00000000001100100101001100100001",
			5241 => "0000001100000000000100010100000100",
			5242 => "11111101101111100101001100100001",
			5243 => "11111111111001000101001100100001",
			5244 => "0000000001000000001100110100001000",
			5245 => "0000000001000000001100110100000100",
			5246 => "11111111000101010101001100100001",
			5247 => "00000000111101110101001100100001",
			5248 => "0000000010000000000011001000000100",
			5249 => "00000000001100110101001100100001",
			5250 => "11111110000001110101001100100001",
			5251 => "0000001001000000001101101000001100",
			5252 => "0000001000000000001111001000001000",
			5253 => "0000000100000000000101010100000100",
			5254 => "00000001110110110101001100100001",
			5255 => "00000000101010010101001100100001",
			5256 => "11111111010101000101001100100001",
			5257 => "0000000100000000001010110100001000",
			5258 => "0000000000000000001111000100000100",
			5259 => "11111111100101100101001100100001",
			5260 => "00000000100011110101001100100001",
			5261 => "0000001011000000001100101100000100",
			5262 => "11111110111000000101001100100001",
			5263 => "00000010110101110101001100100001",
			5264 => "0000000100000000001001001101000000",
			5265 => "0000001001000000001011101000100000",
			5266 => "0000000010000000001110010000010000",
			5267 => "0000001001000000000111100100001000",
			5268 => "0000001000000000000111000100000100",
			5269 => "00000001110001000101001100100001",
			5270 => "11111111100110000101001100100001",
			5271 => "0000000000000000000000110000000100",
			5272 => "00000001010011000101001100100001",
			5273 => "11111110111001110101001100100001",
			5274 => "0000001100000000000000101000001000",
			5275 => "0000001100000000000000101000000100",
			5276 => "00000001010010100101001100100001",
			5277 => "11111111010110000101001100100001",
			5278 => "0000000101000000001100101000000100",
			5279 => "00000001001010100101001100100001",
			5280 => "00000010111111100101001100100001",
			5281 => "0000000010000000001100000000010000",
			5282 => "0000000000000000000000111000001000",
			5283 => "0000001101000000000011100000000100",
			5284 => "00000001101010100101001100100001",
			5285 => "11111111001011110101001100100001",
			5286 => "0000001110000000001101010100000100",
			5287 => "11111101110110010101001100100001",
			5288 => "11111111101110100101001100100001",
			5289 => "0000001110000000000010001000001000",
			5290 => "0000000100000000000011001100000100",
			5291 => "00000101100011100101001100100001",
			5292 => "00000001101011000101001100100001",
			5293 => "0000000111000000000110000100000100",
			5294 => "11111110011100100101001100100001",
			5295 => "00000001110110000101001100100001",
			5296 => "0000001010000000001100000100100000",
			5297 => "0000001000000000001111001000010000",
			5298 => "0000000111000000001100001000001000",
			5299 => "0000001001000000001001111000000100",
			5300 => "11111110101010000101001100100001",
			5301 => "00000010011011110101001100100001",
			5302 => "0000001000000000001111001000000100",
			5303 => "00000000001100110101001100100001",
			5304 => "11111101110110010101001100100001",
			5305 => "0000000000000000001010000000001000",
			5306 => "0000001000000000000111000100000100",
			5307 => "11111101111000110101001100100001",
			5308 => "00000000000001010101001100100001",
			5309 => "0000001110000000001111000100000100",
			5310 => "11111111101100110101001100100001",
			5311 => "00000000011000100101001100100001",
			5312 => "11111110011001010101001100100001",
			5313 => "0000001100000000001010111100001100",
			5314 => "0000000000000000000111000100001000",
			5315 => "0000000000000000001111001000000100",
			5316 => "11111110101001100101001100100001",
			5317 => "00000010110001110101001100100001",
			5318 => "11111110011100010101001100100001",
			5319 => "11111110011001100101001100100001",
			5320 => "0000001111000000000000110111010000",
			5321 => "0000000011000000001001110001101000",
			5322 => "0000001001000000001001111000110000",
			5323 => "0000000001000000001110100000011100",
			5324 => "0000001101000000000110000100010000",
			5325 => "0000000011000000001000111000001000",
			5326 => "0000001111000000000110110100000100",
			5327 => "00000000000011000101010111001101",
			5328 => "11111111001101110101010111001101",
			5329 => "0000001100000000000000110000000100",
			5330 => "11111110000010110101010111001101",
			5331 => "00000001100000110101010111001101",
			5332 => "0000000001000000000110000000001000",
			5333 => "0000001110000000000011111100000100",
			5334 => "11111110110011000101010111001101",
			5335 => "00000001100000100101010111001101",
			5336 => "11111110010001000101010111001101",
			5337 => "0000000010000000000100101000001100",
			5338 => "0000001110000000001110111100001000",
			5339 => "0000001000000000000111000100000100",
			5340 => "00000000000000000101010111001101",
			5341 => "00000001010110100101010111001101",
			5342 => "00000010100011000101010111001101",
			5343 => "0000000011000000000100000000000100",
			5344 => "00000000001011010101010111001101",
			5345 => "11111110001001100101010111001101",
			5346 => "0000000001000000001110100000011000",
			5347 => "0000000111000000000100010100001000",
			5348 => "0000000101000000001101100000000100",
			5349 => "11111110101001010101010111001101",
			5350 => "00000010001111110101010111001101",
			5351 => "0000001100000000000100010100001000",
			5352 => "0000000110000000001110010100000100",
			5353 => "00000000010011110101010111001101",
			5354 => "11111110011011100101010111001101",
			5355 => "0000000111000000000000101000000100",
			5356 => "00000000100101110101010111001101",
			5357 => "11111110001011010101010111001101",
			5358 => "0000001100000000000111111000010000",
			5359 => "0000001100000000000111111000001000",
			5360 => "0000001111000000000101100100000100",
			5361 => "00000000000110100101010111001101",
			5362 => "11111110001101100101010111001101",
			5363 => "0000000011000000001000111100000100",
			5364 => "11111111001111010101010111001101",
			5365 => "11111110000011100101010111001101",
			5366 => "0000000101000000000110000100001000",
			5367 => "0000001000000000000111000100000100",
			5368 => "00000001000000010101010111001101",
			5369 => "11111111100100000101010111001101",
			5370 => "0000000111000000001100001000000100",
			5371 => "11111110000111000101010111001101",
			5372 => "00000000000000000101010111001101",
			5373 => "0000000111000000000100010100101100",
			5374 => "0000000001000000001110100000011100",
			5375 => "0000000100000000001000001000001100",
			5376 => "0000000100000000001100001100001000",
			5377 => "0000001100000000001010000000000100",
			5378 => "00000001001101110101010111001101",
			5379 => "11111111010110110101010111001101",
			5380 => "11111101001011000101010111001101",
			5381 => "0000000010000000001110010000001000",
			5382 => "0000001010000000001010110000000100",
			5383 => "00000000111000100101010111001101",
			5384 => "00000010110000000101010111001101",
			5385 => "0000001000000000000001110100000100",
			5386 => "11111110100000000101010111001101",
			5387 => "00000000011111110101010111001101",
			5388 => "0000000010000000000010011100001100",
			5389 => "0000001101000000001100101100000100",
			5390 => "11111111000100000101010111001101",
			5391 => "0000000101000000001100101100000100",
			5392 => "00000001111101000101010111001101",
			5393 => "00000000101111100101010111001101",
			5394 => "00000010010011000101010111001101",
			5395 => "0000000111000000001000111000100000",
			5396 => "0000001100000000000100000000010000",
			5397 => "0000001100000000000100000000001000",
			5398 => "0000001100000000000000101000000100",
			5399 => "00000000000010110101010111001101",
			5400 => "00000000011011100101010111001101",
			5401 => "0000001010000000001010110000000100",
			5402 => "11111110001001000101010111001101",
			5403 => "00000000100100000101010111001101",
			5404 => "0000000101000000000000001100001000",
			5405 => "0000001101000000000000001100000100",
			5406 => "00000001000001100101010111001101",
			5407 => "00000010110010110101010111001101",
			5408 => "0000001110000000001101100000000100",
			5409 => "11111111011000100101010111001101",
			5410 => "00000001010010100101010111001101",
			5411 => "0000001000000000001111001000010000",
			5412 => "0000000101000000001010111100001000",
			5413 => "0000001110000000000110000100000100",
			5414 => "11111111101110110101010111001101",
			5415 => "00000010001011110101010111001101",
			5416 => "0000001100000000000000101000000100",
			5417 => "11111101111101110101010111001101",
			5418 => "11111111110010110101010111001101",
			5419 => "0000001001000000001101101000001000",
			5420 => "0000000101000000001100101000000100",
			5421 => "11111110101001000101010111001101",
			5422 => "00000000011001010101010111001101",
			5423 => "11111110001010000101010111001101",
			5424 => "0000001110000000000100001001010000",
			5425 => "0000001111000000001101000100110000",
			5426 => "0000001111000000000010110100011100",
			5427 => "0000000010000000001001011100001100",
			5428 => "0000000010000000000111111100001000",
			5429 => "0000000110000000000100110100000100",
			5430 => "11111111010010010101010111001101",
			5431 => "00000000101101000101010111001101",
			5432 => "11111101000011010101010111001101",
			5433 => "0000000111000000001100001000001000",
			5434 => "0000000011000000001110001100000100",
			5435 => "11111111010110000101010111001101",
			5436 => "00000000110100000101010111001101",
			5437 => "0000000111000000000100000000000100",
			5438 => "11111111001010010101010111001101",
			5439 => "00000000001111100101010111001101",
			5440 => "0000000111000000001001110000010000",
			5441 => "0000000110000000001010011000001000",
			5442 => "0000001001000000001101101000000100",
			5443 => "11111111100100110101010111001101",
			5444 => "11111110010011000101010111001101",
			5445 => "0000000010000000000110010000000100",
			5446 => "00000000110001010101010111001101",
			5447 => "11111111001000110101010111001101",
			5448 => "11111101101010110101010111001101",
			5449 => "0000000010000000000110010000000100",
			5450 => "00000010001010010101010111001101",
			5451 => "0000001001000000001101101000001100",
			5452 => "0000000100000000001011100000001000",
			5453 => "0000000001000000000010001100000100",
			5454 => "00000000100011110101010111001101",
			5455 => "00000010000100010101010111001101",
			5456 => "11111110100000010101010111001101",
			5457 => "0000001100000000000100000000001000",
			5458 => "0000000100000000000000010100000100",
			5459 => "11111101100010000101010111001101",
			5460 => "11111111010111110101010111001101",
			5461 => "0000000111000000001001110000000100",
			5462 => "00000000100100100101010111001101",
			5463 => "11111110011010010101010111001101",
			5464 => "0000001110000000000001111100011100",
			5465 => "0000001100000000000100000000010100",
			5466 => "0000000101000000001010111100010000",
			5467 => "0000000011000000001110110000001000",
			5468 => "0000000011000000000111001000000100",
			5469 => "00000000111110000101010111001101",
			5470 => "11111110011100000101010111001101",
			5471 => "0000000010000000000010000100000100",
			5472 => "00000001111111000101010111001101",
			5473 => "00000000100101110101010111001101",
			5474 => "11111101111111000101010111001101",
			5475 => "0000001001000000001111001100000100",
			5476 => "00000010100010000101010111001101",
			5477 => "11111111010000100101010111001101",
			5478 => "0000000111000000000000101000000100",
			5479 => "00000001101101110101010111001101",
			5480 => "0000000001000000001100110100001000",
			5481 => "0000000100000000001001001100000100",
			5482 => "11111111000111010101010111001101",
			5483 => "11111101101001100101010111001101",
			5484 => "0000001111000000001001011100001000",
			5485 => "0000001111000000001110101000000100",
			5486 => "00000000010010110101010111001101",
			5487 => "11111111101100010101010111001101",
			5488 => "0000001111000000000010000000000100",
			5489 => "00000000111110100101010111001101",
			5490 => "11111111100100100101010111001101",
			5491 => "0000001100000000000100001011010100",
			5492 => "0000001111000000001010010101011000",
			5493 => "0000001101000000000111001001000000",
			5494 => "0000001110000000000111111000100000",
			5495 => "0000000111000000001100001000010000",
			5496 => "0000000001000000001100110100001000",
			5497 => "0000000101000000000101101100000100",
			5498 => "00000000001000110101011101111011",
			5499 => "11111111011111000101011101111011",
			5500 => "0000001011000000001100001000000100",
			5501 => "00000011010100110101011101111011",
			5502 => "00000000010000100101011101111011",
			5503 => "0000000101000000000110000100001000",
			5504 => "0000001010000000000110011100000100",
			5505 => "11111110000110000101011101111011",
			5506 => "00000000100001110101011101111011",
			5507 => "0000001001000000000110101000000100",
			5508 => "00000001010010010101011101111011",
			5509 => "11111110100110110101011101111011",
			5510 => "0000000100000000001111100000010000",
			5511 => "0000001001000000000110101000001000",
			5512 => "0000001101000000000101101100000100",
			5513 => "00000000000100000101011101111011",
			5514 => "00000001011100010101011101111011",
			5515 => "0000000001000000001110100000000100",
			5516 => "11111110101010100101011101111011",
			5517 => "00000000010000110101011101111011",
			5518 => "0000000010000000001001011100001000",
			5519 => "0000001010000000000110011100000100",
			5520 => "00000100000001010101011101111011",
			5521 => "11111110101001000101011101111011",
			5522 => "0000001111000000000111110000000100",
			5523 => "11111111100001110101011101111011",
			5524 => "00000010100000110101011101111011",
			5525 => "0000000001000000000010001100001000",
			5526 => "0000001101000000000011100000000100",
			5527 => "11111100000001010101011101111011",
			5528 => "11111110101011110101011101111011",
			5529 => "0000000100000000001000001000001100",
			5530 => "0000001010000000001000010100001000",
			5531 => "0000000100000000001000101000000100",
			5532 => "11111111111100010101011101111011",
			5533 => "11111101001101110101011101111011",
			5534 => "00000001101010100101011101111011",
			5535 => "11111101110110100101011101111011",
			5536 => "0000000110000000001100011000111100",
			5537 => "0000001110000000001101100000100000",
			5538 => "0000001001000000000110101000010000",
			5539 => "0000001010000000000110011000001000",
			5540 => "0000001110000000001001110000000100",
			5541 => "11111101101101100101011101111011",
			5542 => "00000000000000000101011101111011",
			5543 => "0000000010000000001100010100000100",
			5544 => "00000000111011110101011101111011",
			5545 => "11111111010010110101011101111011",
			5546 => "0000000001000000001100110100001000",
			5547 => "0000000010000000001110010000000100",
			5548 => "11111100001011100101011101111011",
			5549 => "11111101111001000101011101111011",
			5550 => "0000001001000000001101101000000100",
			5551 => "00000000000001100101011101111011",
			5552 => "11111110011110010101011101111011",
			5553 => "0000000010000000000110010000010000",
			5554 => "0000001101000000000000001100001000",
			5555 => "0000001100000000001010000000000100",
			5556 => "11111010101110110101011101111011",
			5557 => "00000000111100110101011101111011",
			5558 => "0000000110000000001100011000000100",
			5559 => "11111111111100110101011101111011",
			5560 => "11111101011100010101011101111011",
			5561 => "0000001100000000000100010100000100",
			5562 => "00000000000010110101011101111011",
			5563 => "0000000000000000000010111100000100",
			5564 => "11111111110111000101011101111011",
			5565 => "11111110000011110101011101111011",
			5566 => "0000001001000000001101101000100000",
			5567 => "0000000100000000001111100000010000",
			5568 => "0000001010000000001100011100001000",
			5569 => "0000001101000000001101010100000100",
			5570 => "00000000001100010101011101111011",
			5571 => "00000010010000000101011101111011",
			5572 => "0000001011000000001000111100000100",
			5573 => "00000000111101110101011101111011",
			5574 => "00000010010101000101011101111011",
			5575 => "0000001001000000000110101000001000",
			5576 => "0000000010000000001001100000000100",
			5577 => "11111111010001010101011101111011",
			5578 => "00000001101101010101011101111011",
			5579 => "0000000110000000001101011000000100",
			5580 => "11111110101101000101011101111011",
			5581 => "00000000001101000101011101111011",
			5582 => "0000000010000000000111011000010000",
			5583 => "0000000000000000001110111100001000",
			5584 => "0000001100000000000100010100000100",
			5585 => "11111111000011100101011101111011",
			5586 => "00000000001001010101011101111011",
			5587 => "0000001011000000001000111000000100",
			5588 => "00000000101100000101011101111011",
			5589 => "11111111000010010101011101111011",
			5590 => "0000000010000000000111011000001000",
			5591 => "0000001110000000000100011000000100",
			5592 => "00000011001001010101011101111011",
			5593 => "00000001011000100101011101111011",
			5594 => "0000000100000000001011100000000100",
			5595 => "00000000101011100101011101111011",
			5596 => "11111110011101110101011101111011",
			5597 => "11111110011101110101011101111011",
			5598 => "0000000111000000001101111001110100",
			5599 => "0000000100000000000001001101101000",
			5600 => "0000000000000000000100010100110000",
			5601 => "0000000110000000000001000100010000",
			5602 => "0000000011000000000000111000000100",
			5603 => "00000010100100010101100010000101",
			5604 => "0000000011000000000111111000001000",
			5605 => "0000000011000000001110111100000100",
			5606 => "11111110110011100101100010000101",
			5607 => "00000000011100010101100010000101",
			5608 => "11111110010111010101100010000101",
			5609 => "0000000111000000001100001000010000",
			5610 => "0000000011000000001101100000001000",
			5611 => "0000000111000000000111111000000100",
			5612 => "00000010101010000101100010000101",
			5613 => "00000000100111010101100010000101",
			5614 => "0000000010000000000100101000000100",
			5615 => "00000001101011000101100010000101",
			5616 => "00000000111011110101100010000101",
			5617 => "0000000111000000001100001000001000",
			5618 => "0000001101000000001100101000000100",
			5619 => "11111111011000010101100010000101",
			5620 => "11111101011011110101100010000101",
			5621 => "0000000110000000000001111000000100",
			5622 => "11111110100001100101100010000101",
			5623 => "00000000110011000101100010000101",
			5624 => "0000000110000000001010011000100000",
			5625 => "0000001010000000000110011100010000",
			5626 => "0000000101000000001000111100001000",
			5627 => "0000000010000000000001000000000100",
			5628 => "11111111110000100101100010000101",
			5629 => "00000010111001110101100010000101",
			5630 => "0000001111000000000101100100000100",
			5631 => "11111111000101010101100010000101",
			5632 => "00000000001100010101100010000101",
			5633 => "0000000100000000000001101100001000",
			5634 => "0000001000000000000111000000000100",
			5635 => "00000001101110010101100010000101",
			5636 => "11111110110010100101100010000101",
			5637 => "0000000110000000001100011000000100",
			5638 => "00000011010100010101100010000101",
			5639 => "00000000001001110101100010000101",
			5640 => "0000000010000000001100010000001100",
			5641 => "0000001000000000000010101000000100",
			5642 => "00000000001111010101100010000101",
			5643 => "0000001101000000001110110000000100",
			5644 => "11111110011101010101100010000101",
			5645 => "00000000000000000101100010000101",
			5646 => "0000001011000000001101100000001000",
			5647 => "0000000001000000000010001100000100",
			5648 => "00000000001010100101100010000101",
			5649 => "00000100100101010101100010000101",
			5650 => "11111110010010110101100010000101",
			5651 => "0000000100000000001011100100001000",
			5652 => "0000000110000000001011111100000100",
			5653 => "11111110101110110101100010000101",
			5654 => "00000000001010010101100010000101",
			5655 => "11111110010110100101100010000101",
			5656 => "0000001010000000000111110100010000",
			5657 => "0000000010000000001100111000001100",
			5658 => "0000000111000000001100101000001000",
			5659 => "0000001000000000000000001000000100",
			5660 => "11111110101000110101100010000101",
			5661 => "00000001100101100101100010000101",
			5662 => "11111110010111000101100010000101",
			5663 => "00000101010010100101100010000101",
			5664 => "11111110010110100101100010000101",
			5665 => "0000000010000000001110101001010100",
			5666 => "0000000001000000001001111001001100",
			5667 => "0000001110000000001000111100111000",
			5668 => "0000000101000000001110001100100000",
			5669 => "0000001110000000000000110000010000",
			5670 => "0000001101000000000101101100001000",
			5671 => "0000001111000000001010001100000100",
			5672 => "00000000011010000101101000000001",
			5673 => "11111110101110100101101000000001",
			5674 => "0000000011000000001000111100000100",
			5675 => "11111111101101010101101000000001",
			5676 => "11111110001011000101101000000001",
			5677 => "0000001000000000001001101000001000",
			5678 => "0000000110000000000001111000000100",
			5679 => "00000000110101010101101000000001",
			5680 => "11111110111111100101101000000001",
			5681 => "0000000111000000000000101000000100",
			5682 => "00000010101001000101101000000001",
			5683 => "00000001001010110101101000000001",
			5684 => "0000001111000000001111011100001100",
			5685 => "0000000100000000001010110100001000",
			5686 => "0000000010000000000000110100000100",
			5687 => "11111110111110000101101000000001",
			5688 => "00000001010011000101101000000001",
			5689 => "11111110010110110101101000000001",
			5690 => "0000000101000000001110001100000100",
			5691 => "11111101011101110101101000000001",
			5692 => "0000001101000000001101111000000100",
			5693 => "00000000100010010101101000000001",
			5694 => "11111110101011000101101000000001",
			5695 => "0000001010000000000011101000001100",
			5696 => "0000000100000000000110111100001000",
			5697 => "0000000001000000001100110100000100",
			5698 => "00000000000000000101101000000001",
			5699 => "00000000111111110101101000000001",
			5700 => "11111110100010110101101000000001",
			5701 => "0000001111000000000010001000000100",
			5702 => "00000001111100010101101000000001",
			5703 => "00000000110110010101101000000001",
			5704 => "0000001111000000001001010100000100",
			5705 => "11111101101110010101101000000001",
			5706 => "00000000000000000101101000000001",
			5707 => "0000000010000000001110101000010100",
			5708 => "0000000111000000000000101000001100",
			5709 => "0000001110000000000000110000001000",
			5710 => "0000000111000000001110111100000100",
			5711 => "00000001001100010101101000000001",
			5712 => "11111110001100110101101000000001",
			5713 => "00000000100001110101101000000001",
			5714 => "0000000101000000000011100000000100",
			5715 => "11111101111011110101101000000001",
			5716 => "00000000000000000101101000000001",
			5717 => "0000000011000000000100010100101000",
			5718 => "0000000100000000001011100000001100",
			5719 => "0000000110000000000001111000001000",
			5720 => "0000000001000000000110000000000100",
			5721 => "00000001011010110101101000000001",
			5722 => "11111110100010000101101000000001",
			5723 => "11111110010100100101101000000001",
			5724 => "0000000111000000000100010100010000",
			5725 => "0000000010000000000101110000001000",
			5726 => "0000000011000000001110111100000100",
			5727 => "00000000011000110101101000000001",
			5728 => "00000010001000010101101000000001",
			5729 => "0000001111000000001111011100000100",
			5730 => "00000000000110110101101000000001",
			5731 => "11111110011001100101101000000001",
			5732 => "0000000010000000000101110000000100",
			5733 => "11111110010100010101101000000001",
			5734 => "0000001110000000000111000000000100",
			5735 => "00000000000000000101101000000001",
			5736 => "00000000111011100101101000000001",
			5737 => "0000001101000000000011011100010100",
			5738 => "0000000111000000000100010100010000",
			5739 => "0000001111000000000100010000001000",
			5740 => "0000000100000000001010110100000100",
			5741 => "11111111111000100101101000000001",
			5742 => "00000001100101010101101000000001",
			5743 => "0000000010000000000011001000000100",
			5744 => "11111110001101000101101000000001",
			5745 => "00000000101110100101101000000001",
			5746 => "11111110100101100101101000000001",
			5747 => "0000001111000000001010011100001100",
			5748 => "0000001111000000001010011100001000",
			5749 => "0000001101000000000110000100000100",
			5750 => "11111110010010110101101000000001",
			5751 => "00000001110001110101101000000001",
			5752 => "00000010111110000101101000000001",
			5753 => "0000000011000000000011011100001000",
			5754 => "0000001111000000000110110100000100",
			5755 => "11111111111011100101101000000001",
			5756 => "11111111010001000101101000000001",
			5757 => "0000001001000000000110101000000100",
			5758 => "00000000011010110101101000000001",
			5759 => "11111111111100100101101000000001",
			5760 => "0000001100000000000011011101101000",
			5761 => "0000000100000000000011111001100100",
			5762 => "0000000111000000001001110001000000",
			5763 => "0000001110000000001000111000100000",
			5764 => "0000001111000000000010001000010000",
			5765 => "0000001101000000000000001100001000",
			5766 => "0000000011000000001101100000000100",
			5767 => "00000000011111000101101100100101",
			5768 => "00000001001111000101101100100101",
			5769 => "0000000001000000000010001100000100",
			5770 => "11111110110110000101101100100101",
			5771 => "00000010101010100101101100100101",
			5772 => "0000001010000000001001000100001000",
			5773 => "0000000101000000001101111000000100",
			5774 => "11111110100100010101101100100101",
			5775 => "00000000110011010101101100100101",
			5776 => "0000000000000000000011111100000100",
			5777 => "00000010000001100101101100100101",
			5778 => "00000000000111000101101100100101",
			5779 => "0000001001000000001101101000010000",
			5780 => "0000000111000000001100001000001000",
			5781 => "0000000111000000001100001000000100",
			5782 => "00000000110110000101101100100101",
			5783 => "11111111101100000101101100100101",
			5784 => "0000000100000000001111100000000100",
			5785 => "00000001100000010101101100100101",
			5786 => "11111111110010110101101100100101",
			5787 => "0000001110000000000110000100001000",
			5788 => "0000000001000000000010001100000100",
			5789 => "11111110001001110101101100100101",
			5790 => "11111111101111000101101100100101",
			5791 => "0000000100000000001101001000000100",
			5792 => "00000000111011100101101100100101",
			5793 => "00000000001101010101101100100101",
			5794 => "0000000101000000001100101000000100",
			5795 => "00000001110100110101101100100101",
			5796 => "0000000011000000000100011000010000",
			5797 => "0000000101000000000111001000001000",
			5798 => "0000001111000000001110101100000100",
			5799 => "11111101110100110101101100100101",
			5800 => "11111111101011000101101100100101",
			5801 => "0000000011000000000111001000000100",
			5802 => "00000010110000100101101100100101",
			5803 => "11111110100000010101101100100101",
			5804 => "0000000110000000001011001100001000",
			5805 => "0000001111000000001001010000000100",
			5806 => "00000000000000010101101100100101",
			5807 => "00000001011010010101101100100101",
			5808 => "0000001010000000000110011000000100",
			5809 => "00000001100111100101101100100101",
			5810 => "11111110111111110101101100100101",
			5811 => "11111110011000010101101100100101",
			5812 => "0000001100000000000110000100011000",
			5813 => "0000001011000000001000000000010100",
			5814 => "0000001001000000001101011100000100",
			5815 => "11111110001111110101101100100101",
			5816 => "0000001001000000001101011100000100",
			5817 => "00000010010011100101101100100101",
			5818 => "0000001011000000001010111100001000",
			5819 => "0000001101000000000111010000000100",
			5820 => "11111111000001000101101100100101",
			5821 => "00000001111101100101101100100101",
			5822 => "11111110010111010101101100100101",
			5823 => "00000001100110000101101100100101",
			5824 => "0000001100000000001010111100010000",
			5825 => "0000001010000000000111110100001100",
			5826 => "0000001010000000000111110100000100",
			5827 => "11111110011101010101101100100101",
			5828 => "0000001100000000000000001100000100",
			5829 => "11111111101010000101101100100101",
			5830 => "00000010010010110101101100100101",
			5831 => "11111110011000110101101100100101",
			5832 => "11111110011000000101101100100101",
			5833 => "0000001110000000001000000010001100",
			5834 => "0000001001000000001111001101010100",
			5835 => "0000001011000000000101101101000000",
			5836 => "0000000001000000001110100000100000",
			5837 => "0000001001000000000010001100010000",
			5838 => "0000000011000000001100001000001000",
			5839 => "0000001111000000000001011000000100",
			5840 => "00000000000101110101110011101001",
			5841 => "11111111000111000101110011101001",
			5842 => "0000000101000000001100110000000100",
			5843 => "00000001010011010101110011101001",
			5844 => "11111110100010100101110011101001",
			5845 => "0000000101000000001100110000001000",
			5846 => "0000001010000000001010110000000100",
			5847 => "11111110110101000101110011101001",
			5848 => "11111111100110110101110011101001",
			5849 => "0000001110000000000000110000000100",
			5850 => "11111111000111010101110011101001",
			5851 => "00000001010011110101110011101001",
			5852 => "0000001111000000001111011100010000",
			5853 => "0000001111000000001010011100001000",
			5854 => "0000001011000000001011000100000100",
			5855 => "00000001011011100101110011101001",
			5856 => "11111111111000000101110011101001",
			5857 => "0000001011000000000000101000000100",
			5858 => "00000000011000100101110011101001",
			5859 => "00000001101110010101110011101001",
			5860 => "0000000101000000000011011100001000",
			5861 => "0000001100000000000111111000000100",
			5862 => "11111111111101000101110011101001",
			5863 => "00000001101011010101110011101001",
			5864 => "0000001011000000001011000100000100",
			5865 => "11111111010010100101110011101001",
			5866 => "00000000000001010101110011101001",
			5867 => "0000000101000000001110110000001100",
			5868 => "0000000101000000000111001000000100",
			5869 => "00000000001111100101110011101001",
			5870 => "0000000011000000000011100000000100",
			5871 => "11111111111100100101110011101001",
			5872 => "00000011001100110101110011101001",
			5873 => "0000001001000000001111001100000100",
			5874 => "11111110100100100101110011101001",
			5875 => "00000001010011110101110011101001",
			5876 => "0000000000000000000000110000100000",
			5877 => "0000000001000000001001111000000100",
			5878 => "11111110000000100101110011101001",
			5879 => "0000000111000000001000111000001100",
			5880 => "0000001010000000000110011000001000",
			5881 => "0000000011000000001001001000000100",
			5882 => "11111101011101100101110011101001",
			5883 => "11111111111011100101110011101001",
			5884 => "00000000011011010101110011101001",
			5885 => "0000001001000000001101011100001000",
			5886 => "0000001100000000001001110000000100",
			5887 => "00000001100100000101110011101001",
			5888 => "11111110010100000101110011101001",
			5889 => "0000001010000000000001010000000100",
			5890 => "00000000010110110101110011101001",
			5891 => "11111110111110100101110011101001",
			5892 => "0000001001000000001001011000010000",
			5893 => "0000000110000000001001100100000100",
			5894 => "11111110001101010101110011101001",
			5895 => "0000000101000000000100011000000100",
			5896 => "11111110111011000101110011101001",
			5897 => "0000000001000000001001111000000100",
			5898 => "00000001100010000101110011101001",
			5899 => "00000000000000000101110011101001",
			5900 => "0000001011000000000000001100000100",
			5901 => "00000001100011100101110011101001",
			5902 => "00000000000000000101110011101001",
			5903 => "0000000110000000001001100101000100",
			5904 => "0000001010000000001100011100110000",
			5905 => "0000001100000000000100000000011000",
			5906 => "0000000110000000001011001100001100",
			5907 => "0000000011000000000110100100000100",
			5908 => "11111111101001000101110011101001",
			5909 => "0000001100000000000000101000000100",
			5910 => "00000000101110000101110011101001",
			5911 => "00000001111001010101110011101001",
			5912 => "0000000001000000000111100100001000",
			5913 => "0000000000000000000011111100000100",
			5914 => "11111111001111110101110011101001",
			5915 => "11111101101101010101110011101001",
			5916 => "00000001011010100101110011101001",
			5917 => "0000000001000000001001111000001000",
			5918 => "0000000001000000001001111000000100",
			5919 => "11111111010011110101110011101001",
			5920 => "11111110000010100101110011101001",
			5921 => "0000000110000000001001100100001000",
			5922 => "0000001110000000001010001100000100",
			5923 => "00000000101010010101110011101001",
			5924 => "11111111100110100101110011101001",
			5925 => "0000000101000000001000000000000100",
			5926 => "00000000001010100101110011101001",
			5927 => "00000010101001110101110011101001",
			5928 => "0000001111000000000100101000001000",
			5929 => "0000001100000000000100000000000100",
			5930 => "00000001010101000101110011101001",
			5931 => "11111110010000000101110011101001",
			5932 => "0000001111000000000010000000001000",
			5933 => "0000001100000000000011011100000100",
			5934 => "00000010101000000101110011101001",
			5935 => "11111111101011100101110011101001",
			5936 => "11111110101101100101110011101001",
			5937 => "0000000001000000000110101000001000",
			5938 => "0000001011000000000110000100000100",
			5939 => "00000001000010110101110011101001",
			5940 => "11111110101001100101110011101001",
			5941 => "0000000110000000000100111100000100",
			5942 => "11111110010110100101110011101001",
			5943 => "0000001111000000000010000000000100",
			5944 => "00000001011011000101110011101001",
			5945 => "11111110101011010101110011101001",
			5946 => "0000000111000000001101100010011000",
			5947 => "0000000010000000001110101001001000",
			5948 => "0000000001000000000110000000011100",
			5949 => "0000000101000000000011011100011000",
			5950 => "0000000101000000001001110000001100",
			5951 => "0000000101000000001000111000001000",
			5952 => "0000000011000000000011111100000100",
			5953 => "11111111010010110101111010010101",
			5954 => "00000001010110000101111010010101",
			5955 => "11111110010000110101111010010101",
			5956 => "0000000011000000000000111000000100",
			5957 => "11111110100110100101111010010101",
			5958 => "0000000000000000000000111000000100",
			5959 => "00000000100010010101111010010101",
			5960 => "00000011001011000101111010010101",
			5961 => "11111110010010110101111010010101",
			5962 => "0000001001000000000010001100010000",
			5963 => "0000000111000000000100010100001000",
			5964 => "0000000011000000001110111100000100",
			5965 => "11111111010000100101111010010101",
			5966 => "00000011000100000101111010010101",
			5967 => "0000000101000000000011011100000100",
			5968 => "00000011100101000101111010010101",
			5969 => "00000110101000100101111010010101",
			5970 => "0000000110000000000111101000010000",
			5971 => "0000001110000000000000110000001000",
			5972 => "0000000100000000000110111000000100",
			5973 => "00000001101011100101111010010101",
			5974 => "11111110001111000101111010010101",
			5975 => "0000001010000000000111110100000100",
			5976 => "11111111000110010101111010010101",
			5977 => "00000001110000000101111010010101",
			5978 => "0000000011000000001110111100000100",
			5979 => "11111110010110100101111010010101",
			5980 => "0000000111000000000000101000000100",
			5981 => "00000001010011100101111010010101",
			5982 => "00000000011110110101111010010101",
			5983 => "0000001111000000001001011100111000",
			5984 => "0000001001000000001101011100100000",
			5985 => "0000001010000000001000010100010000",
			5986 => "0000000100000000001110000000001000",
			5987 => "0000000010000000001001010000000100",
			5988 => "00000000101111000101111010010101",
			5989 => "11111111001010000101111010010101",
			5990 => "0000001011000000001100001000000100",
			5991 => "00000000000110000101111010010101",
			5992 => "11111110100000010101111010010101",
			5993 => "0000000100000000001110100100001000",
			5994 => "0000000000000000001111000100000100",
			5995 => "00000000001000010101111010010101",
			5996 => "00000001011000100101111010010101",
			5997 => "0000001010000000000110011000000100",
			5998 => "11111111111000000101111010010101",
			5999 => "00000000010000000101111010010101",
			6000 => "0000000000000000000011111100001100",
			6001 => "0000001111000000001110101100000100",
			6002 => "11111110000011100101111010010101",
			6003 => "0000000110000000001101011000000100",
			6004 => "00000001001110010101111010010101",
			6005 => "11111111100000000101111010010101",
			6006 => "0000001010000000000001010000000100",
			6007 => "11111100101011110101111010010101",
			6008 => "0000001110000000001011000000000100",
			6009 => "11111101111000100101111010010101",
			6010 => "11111111010101000101111010010101",
			6011 => "0000000011000000001001010100010100",
			6012 => "0000001001000000001011111100010000",
			6013 => "0000001000000000000111000100001000",
			6014 => "0000000100000000000010110000000100",
			6015 => "00000001001001100101111010010101",
			6016 => "11111110001000110101111010010101",
			6017 => "0000000100000000000100001100000100",
			6018 => "00000011010010100101111010010101",
			6019 => "11111111100111000101111010010101",
			6020 => "00000110001101010101111010010101",
			6021 => "11111110100011000101111010010101",
			6022 => "0000000011000000001010011100010000",
			6023 => "0000001111000000000010011100001100",
			6024 => "0000001011000000001100101100000100",
			6025 => "11111101110100100101111010010101",
			6026 => "0000001011000000001100101100000100",
			6027 => "00000000000000000101111010010101",
			6028 => "11111110011000010101111010010101",
			6029 => "00000010010001010101111010010101",
			6030 => "0000001001000000000101011100011000",
			6031 => "0000000001000000001001111000000100",
			6032 => "11111110011110110101111010010101",
			6033 => "0000000010000000000010000100001000",
			6034 => "0000000010000000000110010000000100",
			6035 => "00000001111101000101111010010101",
			6036 => "11111110010010010101111010010101",
			6037 => "0000001111000000001110010000001000",
			6038 => "0000000110000000001001100100000100",
			6039 => "00000011001101000101111010010101",
			6040 => "11111111010001110101111010010101",
			6041 => "11111110101011000101111010010101",
			6042 => "0000000111000000000110100100010100",
			6043 => "0000000101000000000001000000010000",
			6044 => "0000001011000000000100001000001000",
			6045 => "0000000100000000001100111000000100",
			6046 => "00000000110001110101111010010101",
			6047 => "11111110001001110101111010010101",
			6048 => "0000000111000000000110000100000100",
			6049 => "00000010010011100101111010010101",
			6050 => "11111111001111000101111010010101",
			6051 => "00000010010010010101111010010101",
			6052 => "11111110011010100101111010010101",
			6053 => "0000001100000000000110000101111000",
			6054 => "0000000100000000000011111001110100",
			6055 => "0000001100000000000000101000111100",
			6056 => "0000001100000000000100010100011100",
			6057 => "0000001100000000000100010100010000",
			6058 => "0000001010000000000001010000001000",
			6059 => "0000000010000000000101110000000100",
			6060 => "00000000011100000101111111010001",
			6061 => "11111111100111000101111111010001",
			6062 => "0000000100000000001001001100000100",
			6063 => "00000001010111000101111111010001",
			6064 => "00000000011100010101111111010001",
			6065 => "0000000100000000000001101100001000",
			6066 => "0000000100000000000011000000000100",
			6067 => "11111100011101010101111111010001",
			6068 => "11111111101111010101111111010001",
			6069 => "00000011010101010101111111010001",
			6070 => "0000001100000000000100010100010000",
			6071 => "0000000011000000000011011100001000",
			6072 => "0000001101000000000110000100000100",
			6073 => "00000001101101010101111111010001",
			6074 => "11111110101110110101111111010001",
			6075 => "0000001101000000001101111000000100",
			6076 => "00000010010000110101111111010001",
			6077 => "00000001000100000101111111010001",
			6078 => "0000000100000000000100001100001000",
			6079 => "0000001000000000000001110100000100",
			6080 => "00000000100100000101111111010001",
			6081 => "00000010110010100101111111010001",
			6082 => "0000000001000000001110100000000100",
			6083 => "00000000111011100101111111010001",
			6084 => "11111110111000010101111111010001",
			6085 => "0000001100000000000000101000011000",
			6086 => "0000001101000000001010111100010000",
			6087 => "0000001000000000001011010100001000",
			6088 => "0000000010000000001100100100000100",
			6089 => "00000000000000000101111111010001",
			6090 => "11111101100000100101111111010001",
			6091 => "0000000101000000001100101000000100",
			6092 => "11111111001000010101111111010001",
			6093 => "00000001110110110101111111010001",
			6094 => "0000001101000000000111001000000100",
			6095 => "11111101001011000101111111010001",
			6096 => "11111110010110110101111111010001",
			6097 => "0000001110000000001001110000010000",
			6098 => "0000001111000000000111010000001000",
			6099 => "0000001110000000000000111000000100",
			6100 => "11111111001111010101111111010001",
			6101 => "00000010010010110101111111010001",
			6102 => "0000000101000000000101101100000100",
			6103 => "00000001001111010101111111010001",
			6104 => "11111111010111000101111111010001",
			6105 => "0000001001000000001101101000001000",
			6106 => "0000001100000000001000111100000100",
			6107 => "00000001011010110101111111010001",
			6108 => "11111110000000110101111111010001",
			6109 => "0000000100000000001001001100000100",
			6110 => "00000000010110010101111111010001",
			6111 => "11111111101110100101111111010001",
			6112 => "11111110011001110101111111010001",
			6113 => "0000001100000000001010111100100100",
			6114 => "0000000111000000001011000000011000",
			6115 => "0000000111000000000100011000010000",
			6116 => "0000000111000000001101111000001100",
			6117 => "0000000111000000001110001100000100",
			6118 => "11111110110101010101111111010001",
			6119 => "0000001100000000000110000100000100",
			6120 => "00000000011010110101111111010001",
			6121 => "00000000000000000101111111010001",
			6122 => "11111110011010010101111111010001",
			6123 => "0000001100000000000100001000000100",
			6124 => "00000010010110000101111111010001",
			6125 => "11111110101101000101111111010001",
			6126 => "0000000111000000001000000000000100",
			6127 => "00000110001000110101111111010001",
			6128 => "0000000100000000001011110000000100",
			6129 => "11111111001011100101111111010001",
			6130 => "00000001011010110101111111010001",
			6131 => "11111110011001000101111111010001",
			6132 => "0000001100000000001000111010011100",
			6133 => "0000000100000000000100001101011100",
			6134 => "0000000011000000000100000000101100",
			6135 => "0000001011000000000100010100010100",
			6136 => "0000000100000000001110000000000100",
			6137 => "00000110001111000110000101110101",
			6138 => "0000000011000000001010000000001000",
			6139 => "0000001011000000000100010100000100",
			6140 => "11111110001100000110000101110101",
			6141 => "00000000000000000110000101110101",
			6142 => "0000001001000000001100110100000100",
			6143 => "00000101101101110110000101110101",
			6144 => "00000000110010000110000101110101",
			6145 => "0000001110000000000000111000001100",
			6146 => "0000001100000000001010000000000100",
			6147 => "00000010001000000110000101110101",
			6148 => "0000000000000000001010000000000100",
			6149 => "11111111011010010110000101110101",
			6150 => "11111110011000000110000101110101",
			6151 => "0000001010000000001000010100000100",
			6152 => "11111110001110000110000101110101",
			6153 => "0000001111000000001111011100000100",
			6154 => "00000101100101100110000101110101",
			6155 => "00000000011010110110000101110101",
			6156 => "0000000011000000000001011000011100",
			6157 => "0000001010000000000111110100001100",
			6158 => "0000000110000000001101111100001000",
			6159 => "0000000110000000001011111100000100",
			6160 => "11111110010100110110000101110101",
			6161 => "00000000001100110110000101110101",
			6162 => "00000100010111010110000101110101",
			6163 => "0000000100000000000110001100001000",
			6164 => "0000000011000000001101100000000100",
			6165 => "00000001001000000110000101110101",
			6166 => "00000011010001110110000101110101",
			6167 => "0000001000000000001001101000000100",
			6168 => "11111111101001110110000101110101",
			6169 => "00000010001010110110000101110101",
			6170 => "0000000000000000001000101100000100",
			6171 => "00000011111111000110000101110101",
			6172 => "0000000000000000000000110000001000",
			6173 => "0000001011000000000000001100000100",
			6174 => "11111110100110010110000101110101",
			6175 => "00000001011001010110000101110101",
			6176 => "0000000001000000000111100100000100",
			6177 => "00000010110111100110000101110101",
			6178 => "11111110011010110110000101110101",
			6179 => "0000001001000000000110000000000100",
			6180 => "11111110010001100110000101110101",
			6181 => "0000000010000000001100010100011100",
			6182 => "0000001011000000000111111000001100",
			6183 => "0000000110000000000001111000000100",
			6184 => "11111110011000100110000101110101",
			6185 => "0000000010000000001101000100000100",
			6186 => "00000000001110100110000101110101",
			6187 => "00000100011110100110000101110101",
			6188 => "0000000000000000001011000100001000",
			6189 => "0000001000000000001010101100000100",
			6190 => "00000000101110100110000101110101",
			6191 => "00000100111000100110000101110101",
			6192 => "0000000100000000000011011000000100",
			6193 => "11111111011000010110000101110101",
			6194 => "00000001000111010110000101110101",
			6195 => "0000000100000000000011101100010000",
			6196 => "0000001010000000001100011100001000",
			6197 => "0000001100000000000111111000000100",
			6198 => "00000010000010010110000101110101",
			6199 => "11111110111101100110000101110101",
			6200 => "0000001001000000001101011100000100",
			6201 => "00000001110101100110000101110101",
			6202 => "11111110001110010110000101110101",
			6203 => "0000001110000000001110001100001000",
			6204 => "0000001010000000001011010100000100",
			6205 => "11111110011100010110000101110101",
			6206 => "00000000000000000110000101110101",
			6207 => "0000000011000000000011100000000100",
			6208 => "00000010110101010110000101110101",
			6209 => "11111110011111100110000101110101",
			6210 => "0000001100000000001100110000101100",
			6211 => "0000001111000000001101000100001100",
			6212 => "0000000011000000000111001000001000",
			6213 => "0000000101000000001010111000000100",
			6214 => "00000000101001000110000101110101",
			6215 => "11111110011010110110000101110101",
			6216 => "11111110010101110110000101110101",
			6217 => "0000000010000000001000001100011000",
			6218 => "0000001011000000000100001000010000",
			6219 => "0000000001000000000110101000001000",
			6220 => "0000001011000000001101111000000100",
			6221 => "00000000000010110110000101110101",
			6222 => "00000011111111000110000101110101",
			6223 => "0000001011000000001101111000000100",
			6224 => "11111111101011000110000101110101",
			6225 => "11111110001100110110000101110101",
			6226 => "0000000101000000001010001100000100",
			6227 => "00000011110010000110000101110101",
			6228 => "00000000101011010110000101110101",
			6229 => "0000001010000000000001010000000100",
			6230 => "00000001000011110110000101110101",
			6231 => "11111110010101000110000101110101",
			6232 => "0000001100000000000100001000001000",
			6233 => "0000001100000000000000001100000100",
			6234 => "11111110010111000110000101110101",
			6235 => "11111111011101100110000101110101",
			6236 => "11111110010001010110000101110101",
			6237 => "0000000111000000000110000110001000",
			6238 => "0000000001000000000000011000001000",
			6239 => "0000000110000000000100110100000100",
			6240 => "11111110010101110110001011011001",
			6241 => "00000001001000010110001011011001",
			6242 => "0000001001000000001001111001000000",
			6243 => "0000000011000000000100000000100000",
			6244 => "0000001001000000001001111000010000",
			6245 => "0000000011000000000100010100001000",
			6246 => "0000001010000000000111110100000100",
			6247 => "00000011000110000110001011011001",
			6248 => "11111111111100110110001011011001",
			6249 => "0000001001000000000010001100000100",
			6250 => "00000001101011110110001011011001",
			6251 => "00000000010101010110001011011001",
			6252 => "0000000001000000001110100000001000",
			6253 => "0000000101000000000011011100000100",
			6254 => "11111111010111000110001011011001",
			6255 => "11111110000110110110001011011001",
			6256 => "0000000001000000001110100000000100",
			6257 => "00000011011111110110001011011001",
			6258 => "11111111110111010110001011011001",
			6259 => "0000001111000000000110110100010000",
			6260 => "0000001000000000001100000100001000",
			6261 => "0000001011000000001011000100000100",
			6262 => "11111110010101000110001011011001",
			6263 => "00000000000011010110001011011001",
			6264 => "0000001010000000001010110000000100",
			6265 => "00000010100011010110001011011001",
			6266 => "00000101100001010110001011011001",
			6267 => "0000000011000000001000111000001000",
			6268 => "0000001001000000000010001100000100",
			6269 => "00000001111111100110001011011001",
			6270 => "11111110110100000110001011011001",
			6271 => "0000000111000000000100010100000100",
			6272 => "00000001111101000110001011011001",
			6273 => "00000000001011110110001011011001",
			6274 => "0000001110000000001000111100100000",
			6275 => "0000001001000000000110101000010000",
			6276 => "0000000011000000000011011100001000",
			6277 => "0000001111000000000110110100000100",
			6278 => "00000000001100110110001011011001",
			6279 => "11111110101101000110001011011001",
			6280 => "0000001011000000000100000000000100",
			6281 => "00000000101001110110001011011001",
			6282 => "00000011000110110110001011011001",
			6283 => "0000001111000000001010010100001000",
			6284 => "0000000101000000000110000100000100",
			6285 => "00000001001100000110001011011001",
			6286 => "11111111101010000110001011011001",
			6287 => "0000000100000000000011010100000100",
			6288 => "11111101101111010110001011011001",
			6289 => "11111111011100010110001011011001",
			6290 => "0000001001000000001101101000010000",
			6291 => "0000000010000000000010000000001000",
			6292 => "0000001010000000001100011100000100",
			6293 => "00000000111010000110001011011001",
			6294 => "00000010011010010110001011011001",
			6295 => "0000001000000000000001110100000100",
			6296 => "11111111000010010110001011011001",
			6297 => "00000000100101100110001011011001",
			6298 => "0000001110000000001101111000001000",
			6299 => "0000000010000000000100101000000100",
			6300 => "00000000001110100110001011011001",
			6301 => "11111111100010010110001011011001",
			6302 => "0000001001000000001111001100000100",
			6303 => "00000000110110110110001011011001",
			6304 => "00000000000001100110001011011001",
			6305 => "0000000111000000001100101000011000",
			6306 => "0000001011000000000001111100000100",
			6307 => "11111110010100100110001011011001",
			6308 => "0000000010000000000111010100010000",
			6309 => "0000000010000000000010000000000100",
			6310 => "11111110100100110110001011011001",
			6311 => "0000000100000000001000110100000100",
			6312 => "00000000010110010110001011011001",
			6313 => "0000000011000000000001001000000100",
			6314 => "00000000110100110110001011011001",
			6315 => "00000011010101100110001011011001",
			6316 => "11111110011101010110001011011001",
			6317 => "0000001010000000000111110100010000",
			6318 => "0000000010000000000001011100001100",
			6319 => "0000000111000000000001111100001000",
			6320 => "0000001111000000000001011000000100",
			6321 => "11111111110001000110001011011001",
			6322 => "00000000101110110110001011011001",
			6323 => "11111110011010000110001011011001",
			6324 => "00000011100010010110001011011001",
			6325 => "11111110011001010110001011011001",
			6326 => "0000000000000000001100001010100100",
			6327 => "0000000010000000000010110101000000",
			6328 => "0000000010000000000001001000011100",
			6329 => "0000000000000000001000110000010100",
			6330 => "0000001011000000001011000100000100",
			6331 => "00000001111010000110010010110101",
			6332 => "0000001100000000001011000100001000",
			6333 => "0000000000000000001011010100000100",
			6334 => "00000000000000000110010010110101",
			6335 => "11111110110010110110010010110101",
			6336 => "0000000110000000001011111100000100",
			6337 => "00000000000000000110010010110101",
			6338 => "00000001011111110110010010110101",
			6339 => "0000001100000000001010000000000100",
			6340 => "00000000000000000110010010110101",
			6341 => "11111110010111100110010010110101",
			6342 => "0000001011000000000100010100010000",
			6343 => "0000001101000000000011011100001100",
			6344 => "0000001111000000001001110100001000",
			6345 => "0000001111000000001011000000000100",
			6346 => "00000001100110010110010010110101",
			6347 => "11111110100011110110010010110101",
			6348 => "00000001101101010110010010110101",
			6349 => "11111110010110100110010010110101",
			6350 => "0000000000000000001110111100010000",
			6351 => "0000001010000000001000010100001000",
			6352 => "0000000000000000001000110000000100",
			6353 => "00000000001000000110010010110101",
			6354 => "00000001111001110110010010110101",
			6355 => "0000001010000000001001000100000100",
			6356 => "11111101111010000110010010110101",
			6357 => "00000000011110110110010010110101",
			6358 => "00000010100111000110010010110101",
			6359 => "0000001010000000001100011100110100",
			6360 => "0000000101000000001001110100100000",
			6361 => "0000000010000000001001100000010000",
			6362 => "0000001111000000000110100000001000",
			6363 => "0000001111000000000010110100000100",
			6364 => "11111111111110000110010010110101",
			6365 => "11111111011101010110010010110101",
			6366 => "0000001110000000000001111100000100",
			6367 => "00000001010000000110010010110101",
			6368 => "00000000000010110110010010110101",
			6369 => "0000000101000000001010111100001000",
			6370 => "0000000101000000000101101100000100",
			6371 => "00000001101001000110010010110101",
			6372 => "11111111000011010110010010110101",
			6373 => "0000001001000000001101011100000100",
			6374 => "00000000101010110110010010110101",
			6375 => "11111110110110100110010010110101",
			6376 => "0000001001000000000101011100000100",
			6377 => "00000001111000010110010010110101",
			6378 => "0000001011000000001110001100001000",
			6379 => "0000000111000000001001110000000100",
			6380 => "00000000000000000110010010110101",
			6381 => "00000010000001010110010010110101",
			6382 => "0000001001000000001011111100000100",
			6383 => "11111110110100000110010010110101",
			6384 => "00000000101000100110010010110101",
			6385 => "0000000101000000001100110000010100",
			6386 => "0000000110000000001100011000001000",
			6387 => "0000000000000000001011000100000100",
			6388 => "00000001001010100110010010110101",
			6389 => "11111110011001110110010010110101",
			6390 => "0000000101000000000011011100000100",
			6391 => "00000000000001110110010010110101",
			6392 => "0000001001000000001001111000000100",
			6393 => "00000010111011010110010010110101",
			6394 => "00000000101100010110010010110101",
			6395 => "0000001100000000000100010100001100",
			6396 => "0000000100000000001111100000001000",
			6397 => "0000001110000000001100001000000100",
			6398 => "11111110110100010110010010110101",
			6399 => "00000001000101100110010010110101",
			6400 => "11111110001111010110010010110101",
			6401 => "0000001001000000000111100100001000",
			6402 => "0000000011000000001101111000000100",
			6403 => "00000000010100100110010010110101",
			6404 => "00000001111101010110010010110101",
			6405 => "0000000110000000001101011000000100",
			6406 => "11111111100000100110010010110101",
			6407 => "00000000010110100110010010110101",
			6408 => "0000000010000000000010000000101100",
			6409 => "0000001110000000000000101000101000",
			6410 => "0000001100000000000100010100011000",
			6411 => "0000000011000000000100000000010000",
			6412 => "0000000011000000001011000100001000",
			6413 => "0000001010000000000110011100000100",
			6414 => "11111110011001100110010010110101",
			6415 => "00000000000010100110010010110101",
			6416 => "0000001010000000000110011100000100",
			6417 => "00000010100010010110010010110101",
			6418 => "00000000011010110110010010110101",
			6419 => "0000001010000000000101000100000100",
			6420 => "11111110010100000110010010110101",
			6421 => "00000000000000000110010010110101",
			6422 => "0000000010000000001010001000000100",
			6423 => "11111110010011110110010010110101",
			6424 => "0000000010000000001010001000001000",
			6425 => "0000000110000000001010011000000100",
			6426 => "00000000000000000110010010110101",
			6427 => "00000001100000000110010010110101",
			6428 => "11111110100101110110010010110101",
			6429 => "00000001010101000110010010110101",
			6430 => "0000000101000000001110001100000100",
			6431 => "11111110010001110110010010110101",
			6432 => "0000001001000000000110101000001100",
			6433 => "0000000010000000000010000100000100",
			6434 => "00000000000000000110010010110101",
			6435 => "0000000000000000000001101000000100",
			6436 => "00000001110001000110010010110101",
			6437 => "00000000000000000110010010110101",
			6438 => "0000001100000000001001110000001000",
			6439 => "0000001110000000001001001000000100",
			6440 => "11111110011011010110010010110101",
			6441 => "00000000100001010110010010110101",
			6442 => "0000000011000000001010111000000100",
			6443 => "00000001011111010110010010110101",
			6444 => "00000000000000000110010010110101",
			6445 => "0000001001000000000110101010001000",
			6446 => "0000001001000000000110101001100000",
			6447 => "0000000000000000000000110000100100",
			6448 => "0000001001000000000110101000010100",
			6449 => "0000001111000000001010010100010000",
			6450 => "0000000100000000001010110100001000",
			6451 => "0000000000000000000000111000000100",
			6452 => "00000000011100010110011010100001",
			6453 => "11111111011111010110011010100001",
			6454 => "0000001111000000000101110100000100",
			6455 => "00000001010110010110011010100001",
			6456 => "11111110010011100110011010100001",
			6457 => "11111101111010110110011010100001",
			6458 => "0000000000000000000000111000001100",
			6459 => "0000000010000000001001010000001000",
			6460 => "0000000110000000000001111000000100",
			6461 => "11111110001100000110011010100001",
			6462 => "00000000001111100110011010100001",
			6463 => "11111101011011010110011010100001",
			6464 => "00000000100101100110011010100001",
			6465 => "0000000011000000001100110000100000",
			6466 => "0000001111000000000110110100010000",
			6467 => "0000000011000000000100000000001000",
			6468 => "0000001000000000001111001000000100",
			6469 => "11111111001100110110011010100001",
			6470 => "11111111111101110110011010100001",
			6471 => "0000001111000000000000011100000100",
			6472 => "00000001111000010110011010100001",
			6473 => "00000000001001000110011010100001",
			6474 => "0000000111000000001011000100001000",
			6475 => "0000000010000000000100101000000100",
			6476 => "11111110011111000110011010100001",
			6477 => "11111111111000110110011010100001",
			6478 => "0000001100000000000111111000000100",
			6479 => "11111111011000100110011010100001",
			6480 => "11111110010110000110011010100001",
			6481 => "0000001100000000000100010100001100",
			6482 => "0000001010000000001100011100001000",
			6483 => "0000001001000000001001111000000100",
			6484 => "00000001010111010110011010100001",
			6485 => "11111111111000100110011010100001",
			6486 => "11111110011001010110011010100001",
			6487 => "0000000001000000001110100000001000",
			6488 => "0000001100000000000000101000000100",
			6489 => "00000000110001010110011010100001",
			6490 => "11111101110111000110011010100001",
			6491 => "0000001100000000000100010100000100",
			6492 => "00000010100001000110011010100001",
			6493 => "00000000111111000110011010100001",
			6494 => "0000000110000000001100011000011100",
			6495 => "0000000010000000001110000100001000",
			6496 => "0000001000000000001100000100000100",
			6497 => "00000001001101000110011010100001",
			6498 => "11111110101011000110011010100001",
			6499 => "0000000011000000001101100000001000",
			6500 => "0000000000000000001010000000000100",
			6501 => "00000001111100000110011010100001",
			6502 => "00000011000101010110011010100001",
			6503 => "0000001101000000001100101100001000",
			6504 => "0000000011000000000101101100000100",
			6505 => "00000010010011010110011010100001",
			6506 => "00000000011010000110011010100001",
			6507 => "00000000001110000110011010100001",
			6508 => "0000000010000000000101110000000100",
			6509 => "00000001011011000110011010100001",
			6510 => "0000000010000000000011001000000100",
			6511 => "11111101111101000110011010100001",
			6512 => "00000000110110000110011010100001",
			6513 => "0000000001000000001110100000001100",
			6514 => "0000001100000000000111111000000100",
			6515 => "11111111100001100110011010100001",
			6516 => "0000000000000000000000110000000100",
			6517 => "11111101000111100110011010100001",
			6518 => "11111110010010100110011010100001",
			6519 => "0000000011000000000101101100111000",
			6520 => "0000001100000000000000101000011100",
			6521 => "0000000000000000001010000000010000",
			6522 => "0000000100000000001000000100001000",
			6523 => "0000000100000000001011110000000100",
			6524 => "00000000000000000110011010100001",
			6525 => "11111101011001010110011010100001",
			6526 => "0000000001000000001100110100000100",
			6527 => "11111111111011010110011010100001",
			6528 => "00000000110100110110011010100001",
			6529 => "0000001101000000000110000100000100",
			6530 => "00000000011110000110011010100001",
			6531 => "0000000111000000000100000000000100",
			6532 => "11111110110011010110011010100001",
			6533 => "00000000101011100110011010100001",
			6534 => "0000001111000000000101100100001100",
			6535 => "0000001100000000000000101000000100",
			6536 => "11111101111110010110011010100001",
			6537 => "0000001100000000000100000000000100",
			6538 => "00000000010011100110011010100001",
			6539 => "11111110001100110110011010100001",
			6540 => "0000001111000000000101110100001000",
			6541 => "0000000011000000000101101100000100",
			6542 => "11111110011111100110011010100001",
			6543 => "11111101010100010110011010100001",
			6544 => "0000000110000000001100011000000100",
			6545 => "00000000001110110110011010100001",
			6546 => "11111110101010110110011010100001",
			6547 => "0000000011000000000110000100010000",
			6548 => "0000000010000000000100101000001000",
			6549 => "0000000010000000000101001000000100",
			6550 => "00000010001011100110011010100001",
			6551 => "11111110100010100110011010100001",
			6552 => "0000001010000000001010110000000100",
			6553 => "00000010111000010110011010100001",
			6554 => "00000000001100010110011010100001",
			6555 => "0000000011000000000110000100001100",
			6556 => "0000000100000000001010110100000100",
			6557 => "11111101100101100110011010100001",
			6558 => "0000001110000000001011000100000100",
			6559 => "11111110001010100110011010100001",
			6560 => "00000000001000010110011010100001",
			6561 => "0000001100000000000111111000001000",
			6562 => "0000001111000000000111110000000100",
			6563 => "00000000001100010110011010100001",
			6564 => "11111110110000110110011010100001",
			6565 => "0000000001000000001110100000000100",
			6566 => "00000000111010000110011010100001",
			6567 => "00000000000000000110011010100001",
			6568 => "0000001100000000000011011101110000",
			6569 => "0000000100000000001011100101101100",
			6570 => "0000000000000000000100010100111100",
			6571 => "0000000111000000001011000100011100",
			6572 => "0000000101000000001100110000010000",
			6573 => "0000001100000000000111111000001000",
			6574 => "0000001001000000001110100000000100",
			6575 => "11111110011010110110100000001101",
			6576 => "00000001010111000110100000001101",
			6577 => "0000000100000000001111100000000100",
			6578 => "00000000010010110110100000001101",
			6579 => "00000011001000010110100000001101",
			6580 => "0000000010000000000000110100000100",
			6581 => "11111110010010110110100000001101",
			6582 => "0000001001000000001001111000000100",
			6583 => "00000011001100000110100000001101",
			6584 => "00000001011010110110100000001101",
			6585 => "0000000110000000000111101000010000",
			6586 => "0000001011000000000100000000001000",
			6587 => "0000000100000000001000011100000100",
			6588 => "00000001011100110110100000001101",
			6589 => "11111110011100010110100000001101",
			6590 => "0000001001000000000001000100000100",
			6591 => "11111110011111000110100000001101",
			6592 => "00000010110110110110100000001101",
			6593 => "0000000100000000000011001100001000",
			6594 => "0000000110000000001101111100000100",
			6595 => "00000000011111000110100000001101",
			6596 => "00000001001100100110100000001101",
			6597 => "0000001010000000000110011000000100",
			6598 => "11111111101111000110100000001101",
			6599 => "00000000101001010110100000001101",
			6600 => "0000000110000000001010011000010100",
			6601 => "0000000110000000001010011000010000",
			6602 => "0000000000000000001000111100001000",
			6603 => "0000000011000000000100010100000100",
			6604 => "11111111011011010110100000001101",
			6605 => "00000000010101100110100000001101",
			6606 => "0000001111000000000111010000000100",
			6607 => "00000010011111010110100000001101",
			6608 => "00000000000000000110100000001101",
			6609 => "00000100001111110110100000001101",
			6610 => "0000000010000000001100010000010000",
			6611 => "0000000000000000001011000100001000",
			6612 => "0000000001000000001100110100000100",
			6613 => "00000001111000110110100000001101",
			6614 => "11111110001110110110100000001101",
			6615 => "0000001101000000001010111000000100",
			6616 => "11111110011110000110100000001101",
			6617 => "00000000001000100110100000001101",
			6618 => "0000000100000000000011101100000100",
			6619 => "00000011000000010110100000001101",
			6620 => "0000001111000000000001000000000100",
			6621 => "11111110010110010110100000001101",
			6622 => "00000000001100000110100000001101",
			6623 => "11111110010111000110100000001101",
			6624 => "0000001100000000000110000100101000",
			6625 => "0000000011000000000110100100000100",
			6626 => "11111110010000000110100000001101",
			6627 => "0000000010000000000111011000010100",
			6628 => "0000000100000000000010110000010000",
			6629 => "0000001001000000001011111100001000",
			6630 => "0000001100000000001100110000000100",
			6631 => "11111110001111000110100000001101",
			6632 => "00000000000000000110100000001101",
			6633 => "0000001011000000001010111100000100",
			6634 => "00000001101111100110100000001101",
			6635 => "11111110011011000110100000001101",
			6636 => "00000010111110000110100000001101",
			6637 => "0000001101000000001001010100001100",
			6638 => "0000000110000000001001100100000100",
			6639 => "11111110010000100110100000001101",
			6640 => "0000000001000000000111100100000100",
			6641 => "00000000011111010110100000001101",
			6642 => "11111110100000100110100000001101",
			6643 => "00000001001111100110100000001101",
			6644 => "0000001100000000001010111100011100",
			6645 => "0000000111000000000110100100011000",
			6646 => "0000000111000000001101111000001100",
			6647 => "0000000000000000000011010000001000",
			6648 => "0000000111000000001110001100000100",
			6649 => "11111110111011110110100000001101",
			6650 => "00000001010101000110100000001101",
			6651 => "11111110011110100110100000001101",
			6652 => "0000000111000000000100011000000100",
			6653 => "11111110010111100110100000001101",
			6654 => "0000000111000000000100011000000100",
			6655 => "00000000110111010110100000001101",
			6656 => "11111110011100100110100000001101",
			6657 => "00000010010011100110100000001101",
			6658 => "11111110010111000110100000001101",
			6659 => "0000001100000000000110000110101100",
			6660 => "0000001001000000000110101001100100",
			6661 => "0000001100000000000100010100111100",
			6662 => "0000000010000000001110101000011100",
			6663 => "0000001110000000000000110000010000",
			6664 => "0000000111000000000000101000001000",
			6665 => "0000000011000000000010111100000100",
			6666 => "11111111010001010110100101111001",
			6667 => "00000000101010010110100101111001",
			6668 => "0000001010000000000001010000000100",
			6669 => "11111110001110000110100101111001",
			6670 => "00000001011001100110100101111001",
			6671 => "0000000000000000000011111100001000",
			6672 => "0000001011000000000000101000000100",
			6673 => "11111111101001010110100101111001",
			6674 => "00000001101100100110100101111001",
			6675 => "00000011011111110110100101111001",
			6676 => "0000001010000000000110011000010000",
			6677 => "0000000010000000000101110000001000",
			6678 => "0000001000000000001011010100000100",
			6679 => "00000000010000110110100101111001",
			6680 => "11111111000011000110100101111001",
			6681 => "0000000000000000000000111000000100",
			6682 => "11111101110100010110100101111001",
			6683 => "00000001010100010110100101111001",
			6684 => "0000000100000000000010111000001000",
			6685 => "0000000010000000000101110000000100",
			6686 => "00000010100001000110100101111001",
			6687 => "00000000001001010110100101111001",
			6688 => "0000001101000000001110001100000100",
			6689 => "00000000001010000110100101111001",
			6690 => "00000010011101000110100101111001",
			6691 => "0000000001000000001100110100100000",
			6692 => "0000001110000000001110111100010000",
			6693 => "0000001101000000000101101100001000",
			6694 => "0000001011000000001011000100000100",
			6695 => "00000000001111100110100101111001",
			6696 => "00000011011101110110100101111001",
			6697 => "0000000010000000001001010000000100",
			6698 => "00000000001100110110100101111001",
			6699 => "11111110101011110110100101111001",
			6700 => "0000000010000000001110010000001000",
			6701 => "0000001010000000000110011100000100",
			6702 => "00000001100011100110100101111001",
			6703 => "00000101100110110110100101111001",
			6704 => "0000000111000000000000101000000100",
			6705 => "00000000110110000110100101111001",
			6706 => "11111110000010000110100101111001",
			6707 => "0000001100000000000000101000000100",
			6708 => "00000001011000100110100101111001",
			6709 => "00000101000100000110100101111001",
			6710 => "0000000001000000001110100000001100",
			6711 => "0000000010000000000011001000001000",
			6712 => "0000000111000000001011000100000100",
			6713 => "11111110010110110110100101111001",
			6714 => "11111100101101000110100101111001",
			6715 => "11111111011000100110100101111001",
			6716 => "0000000011000000001101111000011100",
			6717 => "0000001001000000001101101000010000",
			6718 => "0000000111000000001100001000001000",
			6719 => "0000000111000000001011000100000100",
			6720 => "00000000010100010110100101111001",
			6721 => "11111111101010100110100101111001",
			6722 => "0000000011000000000011011100000100",
			6723 => "11111110001010110110100101111001",
			6724 => "00000000101111100110100101111001",
			6725 => "0000001110000000001100110000001000",
			6726 => "0000001011000000000100000000000100",
			6727 => "11111101111100100110100101111001",
			6728 => "11111111110000100110100101111001",
			6729 => "11111011101111100110100101111001",
			6730 => "0000001001000000000111100100010000",
			6731 => "0000001100000000000000101000001000",
			6732 => "0000000010000000000110010000000100",
			6733 => "00000001010100100110100101111001",
			6734 => "11111111011100010110100101111001",
			6735 => "0000000001000000001100110100000100",
			6736 => "00000001110001010110100101111001",
			6737 => "00000100010100110110100101111001",
			6738 => "0000000011000000000000001100001000",
			6739 => "0000001001000000001101101000000100",
			6740 => "00000001011001000110100101111001",
			6741 => "11111101111010010110100101111001",
			6742 => "0000001110000000001101100000000100",
			6743 => "11111111011010010110100101111001",
			6744 => "00000000001011100110100101111001",
			6745 => "0000001100000000001010111100001000",
			6746 => "0000000101000000001110101000000100",
			6747 => "11111110011100010110100101111001",
			6748 => "00000010001111100110100101111001",
			6749 => "11111110011010100110100101111001",
			6750 => "0000001100000000000110000110111100",
			6751 => "0000001001000000001101101001011100",
			6752 => "0000000111000000000000101000110100",
			6753 => "0000000111000000000000101000011000",
			6754 => "0000001100000000000000101000010000",
			6755 => "0000000010000000000001000000001000",
			6756 => "0000000000000000000100010100000100",
			6757 => "00000000100110010110101100000101",
			6758 => "11111111011100100110101100000101",
			6759 => "0000001010000000001001000100000100",
			6760 => "11111110110110100110101100000101",
			6761 => "00000000000101000110101100000101",
			6762 => "0000000100000000001110111000000100",
			6763 => "11111111110001110110101100000101",
			6764 => "00000011001100000110101100000101",
			6765 => "0000001010000000001010110000010000",
			6766 => "0000001100000000000100010100001000",
			6767 => "0000001111000000001011011100000100",
			6768 => "11111110111111110110101100000101",
			6769 => "11111101110111110110101100000101",
			6770 => "0000000010000000001100100100000100",
			6771 => "11111101110010010110101100000101",
			6772 => "00000000110010000110101100000101",
			6773 => "0000001100000000000111111000000100",
			6774 => "11111110010000100110101100000101",
			6775 => "0000000101000000000110000100000100",
			6776 => "00000001011001010110101100000101",
			6777 => "11111111101001100110101100000101",
			6778 => "0000001010000000000111110100001100",
			6779 => "0000000001000000001100110100001000",
			6780 => "0000000111000000001100001000000100",
			6781 => "11111110111100100110101100000101",
			6782 => "11111101111100000110101100000101",
			6783 => "00000001010001000110101100000101",
			6784 => "0000000100000000000011001100010000",
			6785 => "0000001100000000000111111000001000",
			6786 => "0000001110000000000100000000000100",
			6787 => "11111110111011110110101100000101",
			6788 => "00000000111010000110101100000101",
			6789 => "0000001001000000000111100100000100",
			6790 => "00000001101001100110101100000101",
			6791 => "00000000101110010110101100000101",
			6792 => "0000001101000000001101100000000100",
			6793 => "00000100011000000110101100000101",
			6794 => "0000001110000000001100001000000100",
			6795 => "11111111111000000110101100000101",
			6796 => "00000000100000010110101100000101",
			6797 => "0000001110000000000110000100110000",
			6798 => "0000000001000000001100110100010000",
			6799 => "0000000100000000001100001100000100",
			6800 => "11111100110011010110101100000101",
			6801 => "0000000010000000000100101000000100",
			6802 => "00000001000100110110101100000101",
			6803 => "0000000100000000001010110100000100",
			6804 => "11111100111011010110101100000101",
			6805 => "11111110110011110110101100000101",
			6806 => "0000001101000000001101010100010000",
			6807 => "0000001111000000000001001000001000",
			6808 => "0000001110000000001101100000000100",
			6809 => "11111111101000010110101100000101",
			6810 => "00000000101111000110101100000101",
			6811 => "0000001000000000000110001000000100",
			6812 => "11111110001001100110101100000101",
			6813 => "11111111111101110110101100000101",
			6814 => "0000001100000000001000111000001000",
			6815 => "0000001111000000001110101100000100",
			6816 => "11111110000101010110101100000101",
			6817 => "00000000000000000110101100000101",
			6818 => "0000001000000000000111000100000100",
			6819 => "11111110111010000110101100000101",
			6820 => "00000100000100100110101100000101",
			6821 => "0000001001000000001101101000011000",
			6822 => "0000000010000000001001100000001100",
			6823 => "0000001111000000000110100000001000",
			6824 => "0000001100000000000000101000000100",
			6825 => "00000001111011100110101100000101",
			6826 => "00000000011101000110101100000101",
			6827 => "00000010101111000110101100000101",
			6828 => "0000001000000000000001110100000100",
			6829 => "11111110001110010110101100000101",
			6830 => "0000001011000000001000111000000100",
			6831 => "11111111101011100110101100000101",
			6832 => "00000001111011010110101100000101",
			6833 => "0000001111000000001011110100001100",
			6834 => "0000001100000000000000101000000100",
			6835 => "00000000111100000110101100000101",
			6836 => "0000001111000000000101110100000100",
			6837 => "11111110111100010110101100000101",
			6838 => "11111011001010000110101100000101",
			6839 => "0000001111000000000111110000000100",
			6840 => "00000001111111100110101100000101",
			6841 => "0000001110000000001101111000000100",
			6842 => "11111111100010110110101100000101",
			6843 => "00000000001010000110101100000101",
			6844 => "0000001010000000000111110100001000",
			6845 => "0000000010000000000001011100000100",
			6846 => "11111110100001000110101100000101",
			6847 => "00000001101111100110101100000101",
			6848 => "11111110011011100110101100000101",
			6849 => "0000001100000000000110000111000000",
			6850 => "0000001111000000001011011101010000",
			6851 => "0000000011000000001100110000101000",
			6852 => "0000001001000000000110101000011000",
			6853 => "0000000001000000001100110100010000",
			6854 => "0000001001000000000110101000001000",
			6855 => "0000000011000000000100000000000100",
			6856 => "00000000000110000110110010011001",
			6857 => "00000000110100100110110010011001",
			6858 => "0000001101000000001100101100000100",
			6859 => "00000000100010110110110010011001",
			6860 => "11111111001111110110110010011001",
			6861 => "0000001100000000000100010100000100",
			6862 => "00000011110000100110110010011001",
			6863 => "00000000011110000110110010011001",
			6864 => "0000001110000000000111111000000100",
			6865 => "11111101111101010110110010011001",
			6866 => "0000000010000000001110000100001000",
			6867 => "0000001101000000001101111000000100",
			6868 => "00000001011111010110110010011001",
			6869 => "11111110100110110110110010011001",
			6870 => "11111101100111100110110010011001",
			6871 => "0000001101000000000001111100011100",
			6872 => "0000000100000000000010111000001100",
			6873 => "0000001000000000001011010100001000",
			6874 => "0000001111000000000111010000000100",
			6875 => "00000010000110110110110010011001",
			6876 => "00000000101101010110110010011001",
			6877 => "11111101000010010110110010011001",
			6878 => "0000000010000000001111010000001000",
			6879 => "0000001111000000000101100100000100",
			6880 => "00000011100111110110110010011001",
			6881 => "00000010000001010110110010011001",
			6882 => "0000001110000000000100010100000100",
			6883 => "11111111010001000110110010011001",
			6884 => "00000011000000110110110010011001",
			6885 => "0000001110000000001100110000000100",
			6886 => "11111101101000110110110010011001",
			6887 => "0000000110000000000101011100000100",
			6888 => "11111111000010100110110010011001",
			6889 => "00000010011000110110110010011001",
			6890 => "0000000110000000000100110101000000",
			6891 => "0000000011000000001010111100100000",
			6892 => "0000001110000000001101100000010000",
			6893 => "0000001000000000001001101000001000",
			6894 => "0000000011000000000101101100000100",
			6895 => "11111101111101000110110010011001",
			6896 => "11111111011101110110110010011001",
			6897 => "0000001110000000001001110000000100",
			6898 => "00000000000011010110110010011001",
			6899 => "11111110000100100110110010011001",
			6900 => "0000001101000000000001111100001000",
			6901 => "0000001000000000001001101000000100",
			6902 => "00000001110011010110110010011001",
			6903 => "11111111111000100110110010011001",
			6904 => "0000001111000000000111110000000100",
			6905 => "11111101010011000110110010011001",
			6906 => "11111111001111110110110010011001",
			6907 => "0000001110000000001100101000010000",
			6908 => "0000000010000000000010011100001000",
			6909 => "0000000010000000000101001000000100",
			6910 => "11111101101101100110110010011001",
			6911 => "00000000110011010110110010011001",
			6912 => "0000001001000000001101101000000100",
			6913 => "11111111100101100110110010011001",
			6914 => "11111101011000000110110010011001",
			6915 => "0000001010000000000111110100001000",
			6916 => "0000000100000000001011101100000100",
			6917 => "11111111111011110110110010011001",
			6918 => "11111101001011010110110010011001",
			6919 => "0000000010000000001110010000000100",
			6920 => "00000001101110110110110010011001",
			6921 => "11111111000111100110110010011001",
			6922 => "0000001100000000001010000000010100",
			6923 => "0000000110000000000100110100001000",
			6924 => "0000000010000000000111111100000100",
			6925 => "11111110001101000110110010011001",
			6926 => "00000000100001010110110010011001",
			6927 => "0000000010000000001010001000000100",
			6928 => "11111111101000000110110010011001",
			6929 => "0000001101000000000110000100000100",
			6930 => "11111110011010010110110010011001",
			6931 => "11111100100110010110110010011001",
			6932 => "0000001100000000001110111100001100",
			6933 => "0000000010000000001100010100001000",
			6934 => "0000001010000000001010110000000100",
			6935 => "00000001011011100110110010011001",
			6936 => "11111111001100100110110010011001",
			6937 => "00000010111110100110110010011001",
			6938 => "0000001000000000000001110000001000",
			6939 => "0000000010000000001100010100000100",
			6940 => "00000001111010000110110010011001",
			6941 => "11111111110000000110110010011001",
			6942 => "0000000000000000001000110000000100",
			6943 => "11111110011001010110110010011001",
			6944 => "00000000000111110110110010011001",
			6945 => "0000001010000000000111110100001000",
			6946 => "0000000010000000000001011100000100",
			6947 => "11111110100010010110110010011001",
			6948 => "00000001100101110110110010011001",
			6949 => "11111110011100000110110010011001",
			6950 => "0000001000000000000111000010011100",
			6951 => "0000001010000000000110011101111000",
			6952 => "0000001001000000001001111000111100",
			6953 => "0000000101000000001101100000100000",
			6954 => "0000000000000000000000110000010000",
			6955 => "0000000111000000000111111000001000",
			6956 => "0000000101000000001000111100000100",
			6957 => "00000001011100010110111001010101",
			6958 => "11111110000101000110111001010101",
			6959 => "0000001010000000000110011000000100",
			6960 => "00000000010011010110111001010101",
			6961 => "00000001011110010110111001010101",
			6962 => "0000000000000000000000110000001000",
			6963 => "0000001100000000000111111000000100",
			6964 => "11111110010100100110111001010101",
			6965 => "11111111100011000110111001010101",
			6966 => "0000001110000000000010011000000100",
			6967 => "11111111100111100110111001010101",
			6968 => "00000000001110100110111001010101",
			6969 => "0000001010000000000110011000010000",
			6970 => "0000001001000000000010001100001000",
			6971 => "0000001001000000000010001100000100",
			6972 => "11111110101110110110111001010101",
			6973 => "00000001011010110110111001010101",
			6974 => "0000001110000000000000110000000100",
			6975 => "11111110001010010110111001010101",
			6976 => "00000000000110110110111001010101",
			6977 => "0000000001000000000110000000000100",
			6978 => "11111111011100010110111001010101",
			6979 => "0000000000000000001110111100000100",
			6980 => "00000010100101000110111001010101",
			6981 => "00000001000010110110111001010101",
			6982 => "0000000001000000001110100000011100",
			6983 => "0000000101000000001100110000010000",
			6984 => "0000000101000000000011011100001000",
			6985 => "0000000110000000000100110100000100",
			6986 => "11111111100010010110111001010101",
			6987 => "00000001100000100110111001010101",
			6988 => "0000001111000000000100010000000100",
			6989 => "11111111010111110110111001010101",
			6990 => "11111110010000000110111001010101",
			6991 => "0000000111000000000100010100000100",
			6992 => "00000010000001100110111001010101",
			6993 => "0000001110000000000000110000000100",
			6994 => "11111110110011010110111001010101",
			6995 => "00000000010010000110111001010101",
			6996 => "0000001001000000000110101000010000",
			6997 => "0000000111000000000100010100001000",
			6998 => "0000001001000000000110101000000100",
			6999 => "00000000000011110110111001010101",
			7000 => "11111101101110110110111001010101",
			7001 => "0000001001000000000110101000000100",
			7002 => "00000000011001010110111001010101",
			7003 => "00000001110101110110111001010101",
			7004 => "0000001110000000000000101000001000",
			7005 => "0000000110000000000001111000000100",
			7006 => "11111111000111110110111001010101",
			7007 => "11111111110111100110111001010101",
			7008 => "0000001010000000000110011100000100",
			7009 => "11111111111111100110111001010101",
			7010 => "00000000100110100110111001010101",
			7011 => "0000001001000000000110101000000100",
			7012 => "00000011001010100110111001010101",
			7013 => "0000001011000000001000111100001000",
			7014 => "0000000000000000000000101000000100",
			7015 => "00000000011100100110111001010101",
			7016 => "11111110011000100110111001010101",
			7017 => "0000000101000000000100001000001000",
			7018 => "0000001110000000001101100000000100",
			7019 => "00000000000000000110111001010101",
			7020 => "00000010100011000110111001010101",
			7021 => "0000001111000000001001010000001000",
			7022 => "0000000110000000001001100100000100",
			7023 => "11111110011010000110111001010101",
			7024 => "00000000000000000110111001010101",
			7025 => "0000000001000000001001111000000100",
			7026 => "00000010000111110110111001010101",
			7027 => "11111110100000110110111001010101",
			7028 => "0000000010000000001100000001000000",
			7029 => "0000000010000000001001100000101100",
			7030 => "0000001111000000001111011100011000",
			7031 => "0000001110000000001000110000010000",
			7032 => "0000001100000000001010000000001000",
			7033 => "0000000010000000001110101000000100",
			7034 => "00000000000000000110111001010101",
			7035 => "00000001011010100110111001010101",
			7036 => "0000000110000000000100110100000100",
			7037 => "11111111100111100110111001010101",
			7038 => "11111110001111100110111001010101",
			7039 => "0000000001000000001110100000000100",
			7040 => "00000001010000110110111001010101",
			7041 => "11111110100011110110111001010101",
			7042 => "0000000111000000001011000100001000",
			7043 => "0000000010000000001010001000000100",
			7044 => "11111101111101010110111001010101",
			7045 => "11111111100000010110111001010101",
			7046 => "0000001011000000001100001000001000",
			7047 => "0000001101000000000110000100000100",
			7048 => "11111110111101010110111001010101",
			7049 => "00000000111101100110111001010101",
			7050 => "11111110011011110110111001010101",
			7051 => "0000000101000000001110001100000100",
			7052 => "11111110101001110110111001010101",
			7053 => "0000000110000000001010011000001000",
			7054 => "0000000111000000001010111100000100",
			7055 => "00000011100100010110111001010101",
			7056 => "00000000000000000110111001010101",
			7057 => "0000000110000000001011001100000100",
			7058 => "11111111010001110110111001010101",
			7059 => "00000001100110000110111001010101",
			7060 => "11111110010011010110111001010101",
			7061 => "0000001100000000000011011111001000",
			7062 => "0000000010000000001110101001011000",
			7063 => "0000000001000000000110000000101100",
			7064 => "0000001100000000000111111000011100",
			7065 => "0000000111000000001110111100001100",
			7066 => "0000001011000000001010000000001000",
			7067 => "0000000001000000001110011100000100",
			7068 => "11111110101111000111000000100001",
			7069 => "00000000001111000111000000100001",
			7070 => "11111110000010110111000000100001",
			7071 => "0000000111000000000111111000001000",
			7072 => "0000001011000000000111111000000100",
			7073 => "00000010110001100111000000100001",
			7074 => "11111111011011100111000000100001",
			7075 => "0000001100000000000111111000000100",
			7076 => "11111111100000000111000000100001",
			7077 => "00000100000001110111000000100001",
			7078 => "0000000111000000001011000100001000",
			7079 => "0000000111000000001110111100000100",
			7080 => "11111111011110010111000000100001",
			7081 => "11111110010001010111000000100001",
			7082 => "0000001011000000000100010100000100",
			7083 => "00000001111100100111000000100001",
			7084 => "11111110101001100111000000100001",
			7085 => "0000001001000000000010001100010000",
			7086 => "0000000111000000000100010100001000",
			7087 => "0000000000000000001110111100000100",
			7088 => "00000010001010100111000000100001",
			7089 => "11111111010001100111000000100001",
			7090 => "0000000101000000000011011100000100",
			7091 => "00000010101011000111000000100001",
			7092 => "00000100010101100111000000100001",
			7093 => "0000000110000000000111101000010000",
			7094 => "0000001101000000001100101100001000",
			7095 => "0000001111000000000000011100000100",
			7096 => "11111111110001100111000000100001",
			7097 => "00000010000000010111000000100001",
			7098 => "0000000100000000001111100100000100",
			7099 => "11111111101111000111000000100001",
			7100 => "11111110010000110111000000100001",
			7101 => "0000000001000000000010001100001000",
			7102 => "0000001101000000001100101000000100",
			7103 => "00000000101110110111000000100001",
			7104 => "11111110101111100111000000100001",
			7105 => "00000010010110010111000000100001",
			7106 => "0000001111000000001001010001000000",
			7107 => "0000001101000000000111001000100000",
			7108 => "0000001100000000000100010100010000",
			7109 => "0000001100000000000100010100001000",
			7110 => "0000000111000000001100001000000100",
			7111 => "00000000000110010111000000100001",
			7112 => "00000000110010000111000000100001",
			7113 => "0000001101000000000001111100000100",
			7114 => "11111111100011010111000000100001",
			7115 => "11111101001001110111000000100001",
			7116 => "0000001011000000001100001000001000",
			7117 => "0000000110000000000001111000000100",
			7118 => "11111111001100000111000000100001",
			7119 => "00000001000100100111000000100001",
			7120 => "0000001011000000001100001000000100",
			7121 => "11111111001110010111000000100001",
			7122 => "00000000010010000111000000100001",
			7123 => "0000000100000000001000011100010000",
			7124 => "0000000000000000001101010000001000",
			7125 => "0000000100000000000000010000000100",
			7126 => "00000001111110100111000000100001",
			7127 => "11111111011001010111000000100001",
			7128 => "0000001010000000000110011000000100",
			7129 => "00000001011101010111000000100001",
			7130 => "11111111110010010111000000100001",
			7131 => "0000000000000000000010011000001000",
			7132 => "0000000010000000000011001000000100",
			7133 => "11111100110011100111000000100001",
			7134 => "11111110101100010111000000100001",
			7135 => "0000001001000000001101011100000100",
			7136 => "11111111110011010111000000100001",
			7137 => "11111110110010110111000000100001",
			7138 => "0000001000000000001111001000011100",
			7139 => "0000000000000000000010011000010000",
			7140 => "0000001100000000000100000000001000",
			7141 => "0000001100000000000100000000000100",
			7142 => "00000001000111010111000000100001",
			7143 => "00000111011010100111000000100001",
			7144 => "0000001011000000000100001000000100",
			7145 => "11111110001100010111000000100001",
			7146 => "00000001101101000111000000100001",
			7147 => "0000001100000000001001110000001000",
			7148 => "0000000100000000001100001100000100",
			7149 => "11111101111011110111000000100001",
			7150 => "11111111011100110111000000100001",
			7151 => "00000001110001100111000000100001",
			7152 => "0000000100000000001001000000010000",
			7153 => "0000000110000000001101011000001000",
			7154 => "0000000110000000001101011000000100",
			7155 => "00000000110000010111000000100001",
			7156 => "00000010110011010111000000100001",
			7157 => "0000001111000000000111111100000100",
			7158 => "11111111111111100111000000100001",
			7159 => "00000001100011110111000000100001",
			7160 => "11111110010100100111000000100001",
			7161 => "0000001100000000001010111100011100",
			7162 => "0000000101000000001110101000011000",
			7163 => "0000001100000000000110000100010100",
			7164 => "0000000010000000000111011000001100",
			7165 => "0000000010000000001001100000001000",
			7166 => "0000001100000000001100110000000100",
			7167 => "11111110010110010111000000100001",
			7168 => "00000000000000000111000000100001",
			7169 => "00000000111100010111000000100001",
			7170 => "0000001011000000000011100000000100",
			7171 => "11111110010110100111000000100001",
			7172 => "00000000000000000111000000100001",
			7173 => "11111110011101000111000000100001",
			7174 => "00000010000101000111000000100001",
			7175 => "11111110011010110111000000100001",
			7176 => "0000001100000000001000111011010100",
			7177 => "0000001100000000000111111001101000",
			7178 => "0000001001000000000110101000111100",
			7179 => "0000000011000000001001110000100000",
			7180 => "0000000111000000001011000100010000",
			7181 => "0000000000000000000010111100001000",
			7182 => "0000000101000000000011011100000100",
			7183 => "00000010111101100111001001000101",
			7184 => "11111111010010000111001001000101",
			7185 => "0000000011000000001011000100000100",
			7186 => "11111111100111000111001001000101",
			7187 => "00000000001010010111001001000101",
			7188 => "0000001111000000001010011100001000",
			7189 => "0000000011000000000100010100000100",
			7190 => "11111110101111000111001001000101",
			7191 => "00000001011111010111001001000101",
			7192 => "0000000011000000000100000000000100",
			7193 => "11111110001010010111001001000101",
			7194 => "11111111010110100111001001000101",
			7195 => "0000001111000000000010001000001100",
			7196 => "0000001001000000001001111000000100",
			7197 => "00000000000000000111001001000101",
			7198 => "0000001111000000001011011100000100",
			7199 => "00000010100110100111001001000101",
			7200 => "00000001100110110111001001000101",
			7201 => "0000000101000000001101100000001000",
			7202 => "0000000010000000000011001000000100",
			7203 => "00000000000110000111001001000101",
			7204 => "00000010010011010111001001000101",
			7205 => "0000001010000000001010110000000100",
			7206 => "11111111000011100111001001000101",
			7207 => "00000000101010100111001001000101",
			7208 => "0000000101000000001100110000010000",
			7209 => "0000001011000000000000101000001100",
			7210 => "0000001110000000001000111100001000",
			7211 => "0000001111000000000101110100000100",
			7212 => "11111111000110010111001001000101",
			7213 => "11111101010100010111001001000101",
			7214 => "00000000010101110111001001000101",
			7215 => "11111100111010000111001001000101",
			7216 => "0000001100000000001110111100001100",
			7217 => "0000001010000000001001000100000100",
			7218 => "11111110110101010111001001000101",
			7219 => "0000001100000000001010000000000100",
			7220 => "11111111110111010111001001000101",
			7221 => "00000010001100010111001001000101",
			7222 => "0000000111000000001100001000001000",
			7223 => "0000001110000000001001110000000100",
			7224 => "11111111001110010111001001000101",
			7225 => "00000000000111010111001001000101",
			7226 => "0000000101000000001110001100000100",
			7227 => "00000010011010110111001001000101",
			7228 => "00000000000000000111001001000101",
			7229 => "0000001100000000000100010100101100",
			7230 => "0000001010000000001001000100010100",
			7231 => "0000000111000000000100010100000100",
			7232 => "00000010001001010111001001000101",
			7233 => "0000001100000000000111111000001000",
			7234 => "0000001111000000001011011100000100",
			7235 => "11111101110001100111001001000101",
			7236 => "11111110101011110111001001000101",
			7237 => "0000001001000000000110101000000100",
			7238 => "11111111010101110111001001000101",
			7239 => "00000010001101010111001001000101",
			7240 => "0000000010000000000011001000010000",
			7241 => "0000000111000000000100010100001000",
			7242 => "0000001011000000001110111100000100",
			7243 => "11111110001000110111001001000101",
			7244 => "00000000010100010111001001000101",
			7245 => "0000001001000000001100110100000100",
			7246 => "11111110101111000111001001000101",
			7247 => "00000010010011000111001001000101",
			7248 => "0000000110000000001100011000000100",
			7249 => "11111111000000010111001001000101",
			7250 => "00000001011101110111001001000101",
			7251 => "0000000011000000001100110000100000",
			7252 => "0000001001000000000110101000010000",
			7253 => "0000001100000000000100010100001000",
			7254 => "0000001100000000000100010100000100",
			7255 => "11111111011011000111001001000101",
			7256 => "00000000110111010111001001000101",
			7257 => "0000001111000000000101100100000100",
			7258 => "00000000000111000111001001000101",
			7259 => "11111111011111010111001001000101",
			7260 => "0000001000000000001011010100001000",
			7261 => "0000001101000000001101111000000100",
			7262 => "00000000101100000111001001000101",
			7263 => "11111101110111110111001001000101",
			7264 => "0000001111000000000110110100000100",
			7265 => "11111101111001000111001001000101",
			7266 => "00000000000000000111001001000101",
			7267 => "0000001001000000000111100100010000",
			7268 => "0000000011000000001101111000001000",
			7269 => "0000001111000000001010010100000100",
			7270 => "00000000101001100111001001000101",
			7271 => "11111111100101110111001001000101",
			7272 => "0000001100000000000100010100000100",
			7273 => "11111111111001000111001001000101",
			7274 => "00000001111111100111001001000101",
			7275 => "0000001011000000001100001000001000",
			7276 => "0000001100000000000000101000000100",
			7277 => "11111111001101110111001001000101",
			7278 => "00000000111111110111001001000101",
			7279 => "0000000011000000000101101100000100",
			7280 => "11111110110001100111001001000101",
			7281 => "00000000000101000111001001000101",
			7282 => "0000001111000000001101000100011000",
			7283 => "0000000101000000001000000000001100",
			7284 => "0000001110000000000110000100001000",
			7285 => "0000000000000000000000111000000100",
			7286 => "00000001001101100111001001000101",
			7287 => "11111110011101010111001001000101",
			7288 => "11111101110011100111001001000101",
			7289 => "0000000101000000001000000000001000",
			7290 => "0000000010000000000010011100000100",
			7291 => "00000000000000000111001001000101",
			7292 => "00000011011101110111001001000101",
			7293 => "11111110110011000111001001000101",
			7294 => "0000001001000000001111001100001000",
			7295 => "0000000110000000001101011000000100",
			7296 => "00000010110001110111001001000101",
			7297 => "11111110100000100111001001000101",
			7298 => "0000001011000000001101111000000100",
			7299 => "11111110010111100111001001000101",
			7300 => "0000001111000000001110010000010000",
			7301 => "0000000010000000001001100000001000",
			7302 => "0000001101000000000111010000000100",
			7303 => "11111110101010100111001001000101",
			7304 => "00000001001110110111001001000101",
			7305 => "0000001001000000000101011100000100",
			7306 => "00000010110101100111001001000101",
			7307 => "11111111001000000111001001000101",
			7308 => "0000001010000000000111110100001000",
			7309 => "0000000111000000001101010100000100",
			7310 => "00000001001011110111001001000101",
			7311 => "11111111001011100111001001000101",
			7312 => "11111110011110110111001001000101",
			7313 => "0000000010000000000000010011000100",
			7314 => "0000001010000000001010110001101000",
			7315 => "0000000000000000000111111001000000",
			7316 => "0000000010000000001110101000100000",
			7317 => "0000000110000000000111101000010000",
			7318 => "0000001100000000000111111000001000",
			7319 => "0000000000000000001111000100000100",
			7320 => "00000001101100110111001111100001",
			7321 => "00000000000000000111001111100001",
			7322 => "0000000011000000001001110000000100",
			7323 => "11111110101100010111001111100001",
			7324 => "11111111110100100111001111100001",
			7325 => "0000001100000000000111111000001000",
			7326 => "0000000011000000000111111000000100",
			7327 => "11111110100100010111001111100001",
			7328 => "00000000000101100111001111100001",
			7329 => "0000001111000000000001101000000100",
			7330 => "00000001101011000111001111100001",
			7331 => "00000000100000000111001111100001",
			7332 => "0000000001000000000110000000010000",
			7333 => "0000001101000000001101100000001000",
			7334 => "0000001011000000000100010100000100",
			7335 => "00000000110100010111001111100001",
			7336 => "11111111010010010111001111100001",
			7337 => "0000000111000000000100010100000100",
			7338 => "00000001111111010111001111100001",
			7339 => "11111110111101100111001111100001",
			7340 => "0000000011000000001000111000001000",
			7341 => "0000001011000000000100010100000100",
			7342 => "00000000010011010111001111100001",
			7343 => "11111111000111010111001111100001",
			7344 => "0000001111000000000101110100000100",
			7345 => "00000000001101010111001111100001",
			7346 => "11111111111010100111001111100001",
			7347 => "0000001011000000001011000100100000",
			7348 => "0000000110000000001101111100010000",
			7349 => "0000000100000000000011110100001000",
			7350 => "0000001101000000001100110000000100",
			7351 => "11111110001110110111001111100001",
			7352 => "11111111110010110111001111100001",
			7353 => "0000001000000000000001110100000100",
			7354 => "11111110001110000111001111100001",
			7355 => "00000001000001110111001111100001",
			7356 => "0000000110000000000100110100001000",
			7357 => "0000000100000000000011010100000100",
			7358 => "11111111001111000111001111100001",
			7359 => "00000001111110100111001111100001",
			7360 => "0000000010000000000100101000000100",
			7361 => "11111111101000100111001111100001",
			7362 => "11111110000010110111001111100001",
			7363 => "0000000100000000000010100100000100",
			7364 => "11111110000110000111001111100001",
			7365 => "11111111100101110111001111100001",
			7366 => "0000000100000000001001001100100100",
			7367 => "0000000010000000001100000000011100",
			7368 => "0000001011000000001001110000010000",
			7369 => "0000001111000000000111110000001000",
			7370 => "0000000100000000000101010100000100",
			7371 => "11111101110100110111001111100001",
			7372 => "11111111001000010111001111100001",
			7373 => "0000001100000000000000101000000100",
			7374 => "00000001010100100111001111100001",
			7375 => "11111111001100010111001111100001",
			7376 => "0000000000000000000000111000000100",
			7377 => "00000000111010100111001111100001",
			7378 => "0000001111000000001110000100000100",
			7379 => "11111101111011000111001111100001",
			7380 => "11111111011110010111001111100001",
			7381 => "0000001101000000001001001000000100",
			7382 => "00000010100001100111001111100001",
			7383 => "11111110101110000111001111100001",
			7384 => "0000000000000000000100010100011100",
			7385 => "0000001111000000000110110100001100",
			7386 => "0000000100000000000000010100000100",
			7387 => "11111111111000100111001111100001",
			7388 => "0000001011000000000000101000000100",
			7389 => "00000001011010100111001111100001",
			7390 => "00000011000001100111001111100001",
			7391 => "0000000100000000000000010100001000",
			7392 => "0000000100000000000000010100000100",
			7393 => "00000000101010010111001111100001",
			7394 => "00000010000110110111001111100001",
			7395 => "0000000111000000001101100000000100",
			7396 => "00000000000100000111001111100001",
			7397 => "00000001100111110111001111100001",
			7398 => "0000000100000000000011010100001100",
			7399 => "0000001000000000000010101000000100",
			7400 => "11111101111111110111001111100001",
			7401 => "0000000000000000001011000100000100",
			7402 => "00000001000000010111001111100001",
			7403 => "11111110000110110111001111100001",
			7404 => "0000000111000000000000101000001000",
			7405 => "0000000100000000000010100100000100",
			7406 => "11111111010000110111001111100001",
			7407 => "00000000000111110111001111100001",
			7408 => "0000001101000000001100110000000100",
			7409 => "00000011010110110111001111100001",
			7410 => "00000000011001110111001111100001",
			7411 => "0000001010000000000111110100001000",
			7412 => "0000001100000000001101010100000100",
			7413 => "00000001011101010111001111100001",
			7414 => "11111111100101100111001111100001",
			7415 => "11111110010110010111001111100001",
			7416 => "0000000010000000000010110101010100",
			7417 => "0000000110000000000100110101001100",
			7418 => "0000000110000000000001111000100100",
			7419 => "0000001000000000001100000100010100",
			7420 => "0000000010000000001110101100010000",
			7421 => "0000000101000000001100110000001000",
			7422 => "0000000000000000001111000100000100",
			7423 => "00000001010100110111010111111101",
			7424 => "11111111001111000111010111111101",
			7425 => "0000001111000000000000011100000100",
			7426 => "11111111000010010111010111111101",
			7427 => "00000001000011100111010111111101",
			7428 => "00000001100111010111010111111101",
			7429 => "0000001011000000000100010100001100",
			7430 => "0000000111000000000100010100001000",
			7431 => "0000001011000000001110111100000100",
			7432 => "00000001111101000111010111111101",
			7433 => "11111110110110100111010111111101",
			7434 => "00000010110000110111010111111101",
			7435 => "11111110011000110111010111111101",
			7436 => "0000001011000000000111111000010000",
			7437 => "0000000110000000001101111100001100",
			7438 => "0000001111000000000011100000001000",
			7439 => "0000001100000000001010000000000100",
			7440 => "00000000000000000111010111111101",
			7441 => "00000010010101110111010111111101",
			7442 => "11111110101110100111010111111101",
			7443 => "11111110011011100111010111111101",
			7444 => "0000001100000000000111111000001000",
			7445 => "0000001000000000000111000100000100",
			7446 => "11111111110101100111010111111101",
			7447 => "00000001011101100111010111111101",
			7448 => "0000000101000000000110000100001000",
			7449 => "0000000001000000000110000000000100",
			7450 => "00000000110100000111010111111101",
			7451 => "00000010010110100111010111111101",
			7452 => "0000001100000000000000101000000100",
			7453 => "11111111011101010111010111111101",
			7454 => "00000001011101110111010111111101",
			7455 => "0000001111000000001010111000000100",
			7456 => "00000000000000000111010111111101",
			7457 => "11111110011010110111010111111101",
			7458 => "0000001001000000001001111001101100",
			7459 => "0000000011000000001100001000111100",
			7460 => "0000001111000000000000011100011100",
			7461 => "0000000100000000000010111000001100",
			7462 => "0000001001000000001001111000001000",
			7463 => "0000001000000000001011010100000100",
			7464 => "00000000100110110111010111111101",
			7465 => "11111110011010110111010111111101",
			7466 => "11111110001111100111010111111101",
			7467 => "0000001110000000000011111100001000",
			7468 => "0000001000000000000110001000000100",
			7469 => "00000001010100000111010111111101",
			7470 => "11111111110111110111010111111101",
			7471 => "0000001000000000000001110100000100",
			7472 => "00000000100111100111010111111101",
			7473 => "00000010001111110111010111111101",
			7474 => "0000001011000000000100010100010000",
			7475 => "0000001011000000000111111000001000",
			7476 => "0000000001000000000110000000000100",
			7477 => "00000000000000000111010111111101",
			7478 => "11111110010111000111010111111101",
			7479 => "0000000111000000000111111000000100",
			7480 => "00000010101111010111010111111101",
			7481 => "11111111101010110111010111111101",
			7482 => "0000001001000000000010001100001000",
			7483 => "0000000110000000001101111100000100",
			7484 => "11111111000110100111010111111101",
			7485 => "00000001010001110111010111111101",
			7486 => "0000000000000000000100010100000100",
			7487 => "11111110000100010111010111111101",
			7488 => "11111110111011110111010111111101",
			7489 => "0000001111000000000010001000011000",
			7490 => "0000001000000000001100000100001000",
			7491 => "0000000011000000001000111000000100",
			7492 => "11111110010010000111010111111101",
			7493 => "00000000010011100111010111111101",
			7494 => "0000000100000000001001000000001000",
			7495 => "0000000100000000000011101100000100",
			7496 => "00000000110001100111010111111101",
			7497 => "00000010011100000111010111111101",
			7498 => "0000000011000000000100000000000100",
			7499 => "00000000000000000111010111111101",
			7500 => "11111110110011000111010111111101",
			7501 => "0000001000000000000010101000010000",
			7502 => "0000001000000000000001110100001000",
			7503 => "0000000100000000001010110100000100",
			7504 => "00000001001100000111010111111101",
			7505 => "11111111010111000111010111111101",
			7506 => "0000000111000000000100010100000100",
			7507 => "00000001111001100111010111111101",
			7508 => "00000000000001110111010111111101",
			7509 => "0000000111000000000000101000000100",
			7510 => "11111110001010100111010111111101",
			7511 => "00000000000000000111010111111101",
			7512 => "0000000001000000001110100000101100",
			7513 => "0000000101000000000011011100001100",
			7514 => "0000001100000000000111111000000100",
			7515 => "11111111010111110111010111111101",
			7516 => "0000001001000000001001111000000100",
			7517 => "00000010100111110111010111111101",
			7518 => "00000000010100100111010111111101",
			7519 => "0000001100000000000111111000010000",
			7520 => "0000000010000000000001000000001000",
			7521 => "0000000100000000000110001100000100",
			7522 => "11111111101100010111010111111101",
			7523 => "00000001111011000111010111111101",
			7524 => "0000000011000000001001110000000100",
			7525 => "11111110010100100111010111111101",
			7526 => "00000000001101000111010111111101",
			7527 => "0000001100000000000100010100001000",
			7528 => "0000000000000000000100000000000100",
			7529 => "11111111001100110111010111111101",
			7530 => "00000000110100000111010111111101",
			7531 => "0000001100000000000000101000000100",
			7532 => "00000000100001100111010111111101",
			7533 => "11111111000100010111010111111101",
			7534 => "0000000011000000001100001000000100",
			7535 => "00000001111111000111010111111101",
			7536 => "0000001100000000000111111000010000",
			7537 => "0000000101000000000101101100001000",
			7538 => "0000000101000000001101100000000100",
			7539 => "00000000011101000111010111111101",
			7540 => "11111110001010110111010111111101",
			7541 => "0000001000000000001100000100000100",
			7542 => "11111110110100010111010111111101",
			7543 => "00000000000010110111010111111101",
			7544 => "0000001011000000001100001000001000",
			7545 => "0000000111000000001100001000000100",
			7546 => "00000000001011110111010111111101",
			7547 => "00000001000001100111010111111101",
			7548 => "0000000011000000001001110000000100",
			7549 => "11111110100110100111010111111101",
			7550 => "11111111111100110111010111111101",
			7551 => "0000001000000000000111000011001000",
			7552 => "0000000110000000001101011001110100",
			7553 => "0000001100000000000000101000111000",
			7554 => "0000001100000000000100010100100000",
			7555 => "0000001100000000000100010100010000",
			7556 => "0000000111000000001100001000001000",
			7557 => "0000000111000000001100001000000100",
			7558 => "00000000000101010111100000011001",
			7559 => "11111110111111010111100000011001",
			7560 => "0000000010000000001100010100000100",
			7561 => "00000001000100110111100000011001",
			7562 => "11111111011100000111100000011001",
			7563 => "0000001100000000000100010100001000",
			7564 => "0000000100000000001011110000000100",
			7565 => "11111110001011100111100000011001",
			7566 => "11111111100101100111100000011001",
			7567 => "0000001101000000001100101100000100",
			7568 => "00000000110011110111100000011001",
			7569 => "11111111110001010111100000011001",
			7570 => "0000000111000000000000101000001100",
			7571 => "0000000100000000001001001100001000",
			7572 => "0000000111000000000000101000000100",
			7573 => "00000000011110110111100000011001",
			7574 => "00000010011111100111100000011001",
			7575 => "00000010110010000111100000011001",
			7576 => "0000001110000000001100101100001000",
			7577 => "0000000010000000000101110000000100",
			7578 => "00000000111011000111100000011001",
			7579 => "11111111001100100111100000011001",
			7580 => "00000001111110110111100000011001",
			7581 => "0000001100000000000000101000011100",
			7582 => "0000000010000000001110000100001100",
			7583 => "0000000001000000001100110100001000",
			7584 => "0000000111000000001100001000000100",
			7585 => "00000000111011000111100000011001",
			7586 => "11111110011000110111100000011001",
			7587 => "00000001101110000111100000011001",
			7588 => "0000001010000000001000010100001000",
			7589 => "0000000001000000000010001100000100",
			7590 => "11111100111011010111100000011001",
			7591 => "11111110111011110111100000011001",
			7592 => "0000000100000000000011001100000100",
			7593 => "00000000011001000111100000011001",
			7594 => "11111110111110100111100000011001",
			7595 => "0000001100000000000000101000010000",
			7596 => "0000001110000000001101111000001000",
			7597 => "0000001101000000001100101000000100",
			7598 => "00000000101101000111100000011001",
			7599 => "11111111010001110111100000011001",
			7600 => "0000001101000000000001111100000100",
			7601 => "00000000000000000111100000011001",
			7602 => "00000001111110100111100000011001",
			7603 => "0000001100000000000000101000001000",
			7604 => "0000000110000000000001111000000100",
			7605 => "11111110100001110111100000011001",
			7606 => "11111111100111110111100000011001",
			7607 => "0000001100000000000000101000000100",
			7608 => "00000000111101000111100000011001",
			7609 => "11111111111010100111100000011001",
			7610 => "0000000111000000001000111000100000",
			7611 => "0000001101000000001100101000001100",
			7612 => "0000000100000000000100001100001000",
			7613 => "0000000011000000000100001000000100",
			7614 => "00000000000000000111100000011001",
			7615 => "00000001110111000111100000011001",
			7616 => "11111110001100010111100000011001",
			7617 => "0000001001000000001101101000001000",
			7618 => "0000001011000000001000111100000100",
			7619 => "00000000000000000111100000011001",
			7620 => "00000010110001110111100000011001",
			7621 => "0000000001000000000010001100000100",
			7622 => "11111110101011110111100000011001",
			7623 => "0000001110000000001010111100000100",
			7624 => "00000000010000100111100000011001",
			7625 => "00000001010100000111100000011001",
			7626 => "0000000010000000000010000000010100",
			7627 => "0000000000000000000000111000001100",
			7628 => "0000000011000000001010011100000100",
			7629 => "00000001010001110111100000011001",
			7630 => "0000000011000000000000011100000100",
			7631 => "11111110000011100111100000011001",
			7632 => "00000000011100110111100000011001",
			7633 => "0000000010000000001100010100000100",
			7634 => "11111101110011110111100000011001",
			7635 => "11111110111001010111100000011001",
			7636 => "0000000110000000001011001100010000",
			7637 => "0000001100000000001000111000001000",
			7638 => "0000001011000000001101100000000100",
			7639 => "00000000001000000111100000011001",
			7640 => "00000001101100100111100000011001",
			7641 => "0000001110000000000110100100000100",
			7642 => "11111110011000100111100000011001",
			7643 => "00000000111101110111100000011001",
			7644 => "0000000011000000001111011100001000",
			7645 => "0000000000000000001011000100000100",
			7646 => "11111110011110100111100000011001",
			7647 => "00000000100100000111100000011001",
			7648 => "0000000011000000000100000100000100",
			7649 => "00000001101010100111100000011001",
			7650 => "11111111111001100111100000011001",
			7651 => "0000000010000000001100000001000100",
			7652 => "0000000010000000001001100000110100",
			7653 => "0000001100000000000111111000011000",
			7654 => "0000001011000000000100010100010000",
			7655 => "0000001001000000001100110100001000",
			7656 => "0000000011000000001000110000000100",
			7657 => "11111110111101000111100000011001",
			7658 => "00000001010100010111100000011001",
			7659 => "0000001110000000001000110000000100",
			7660 => "11111111010100010111100000011001",
			7661 => "11111110010001110111100000011001",
			7662 => "0000001101000000000011011100000100",
			7663 => "11111110111111010111100000011001",
			7664 => "00000011000100000111100000011001",
			7665 => "0000000111000000001011000100010000",
			7666 => "0000000100000000000010010000001000",
			7667 => "0000001101000000001001110000000100",
			7668 => "11111111001110010111100000011001",
			7669 => "11111110001000100111100000011001",
			7670 => "0000000110000000000100110100000100",
			7671 => "00000000111011100111100000011001",
			7672 => "11111111010001110111100000011001",
			7673 => "0000000111000000001100001000001000",
			7674 => "0000001000000000001000110000000100",
			7675 => "00000000111010110111100000011001",
			7676 => "11111111010110010111100000011001",
			7677 => "11111110011011000111100000011001",
			7678 => "0000001010000000000101000100000100",
			7679 => "11111110110000100111100000011001",
			7680 => "0000001110000000001100001000001000",
			7681 => "0000000010000000001100000000000100",
			7682 => "11111111000011100111100000011001",
			7683 => "00000000111110010111100000011001",
			7684 => "00000010010010100111100000011001",
			7685 => "11111110010110010111100000011001",
			7686 => "0000001110000000000101101111001000",
			7687 => "0000001100000000000100010101011100",
			7688 => "0000001100000000000100010101000000",
			7689 => "0000000100000000001101001000100000",
			7690 => "0000000000000000000011010000010000",
			7691 => "0000000100000000001000001000001000",
			7692 => "0000000010000000000101110000000100",
			7693 => "00000000000000000111101010100101",
			7694 => "11111101111111000111101010100101",
			7695 => "0000001110000000000100010100000100",
			7696 => "00000010010101110111101010100101",
			7697 => "00000000001111110111101010100101",
			7698 => "0000001110000000001011000100001000",
			7699 => "0000001000000000001011010100000100",
			7700 => "11111110100001110111101010100101",
			7701 => "11111111110001000111101010100101",
			7702 => "0000001010000000000001010000000100",
			7703 => "11111101110110000111101010100101",
			7704 => "00000000010111000111101010100101",
			7705 => "0000000010000000000010000000010000",
			7706 => "0000000000000000000100010100001000",
			7707 => "0000001000000000000001110100000100",
			7708 => "00000000010001000111101010100101",
			7709 => "00000010101001110111101010100101",
			7710 => "0000001010000000001010110000000100",
			7711 => "11111110010011110111101010100101",
			7712 => "00000000000010100111101010100101",
			7713 => "0000001100000000001110111100001000",
			7714 => "0000000100000000001011100000000100",
			7715 => "00000001000110000111101010100101",
			7716 => "11111110100101110111101010100101",
			7717 => "0000000101000000001100101100000100",
			7718 => "11111110010100010111101010100101",
			7719 => "11111111111101100111101010100101",
			7720 => "0000001011000000001011000100001000",
			7721 => "0000000000000000000111111000000100",
			7722 => "11111110010111010111101010100101",
			7723 => "00000000110011100111101010100101",
			7724 => "0000001000000000001100000100000100",
			7725 => "00000011110010010111101010100101",
			7726 => "0000000110000000000100110100001000",
			7727 => "0000000101000000000101101100000100",
			7728 => "00000010001110110111101010100101",
			7729 => "11111111100010000111101010100101",
			7730 => "0000000110000000001100011000000100",
			7731 => "00000011011010100111101010100101",
			7732 => "00000000011000110111101010100101",
			7733 => "0000001100000000000100010100101100",
			7734 => "0000001010000000000110011100011100",
			7735 => "0000000010000000001110000100010000",
			7736 => "0000001110000000000000101000001000",
			7737 => "0000001010000000001001000100000100",
			7738 => "11111110110110000111101010100101",
			7739 => "00000000011000100111101010100101",
			7740 => "0000001000000000000001110000000100",
			7741 => "11111111110001010111101010100101",
			7742 => "00000001101010100111101010100101",
			7743 => "0000001101000000001101100000000100",
			7744 => "00000000111100010111101010100101",
			7745 => "0000000011000000001101111000000100",
			7746 => "11111110111100110111101010100101",
			7747 => "11111111111011010111101010100101",
			7748 => "0000000111000000001100001000001100",
			7749 => "0000001011000000001100001000001000",
			7750 => "0000001010000000000101000100000100",
			7751 => "00000001000001110111101010100101",
			7752 => "11111111000101000111101010100101",
			7753 => "11111110010110000111101010100101",
			7754 => "00000010011110110111101010100101",
			7755 => "0000001011000000001100001000100000",
			7756 => "0000001011000000000000101000010000",
			7757 => "0000000101000000000101101100001000",
			7758 => "0000000001000000001110100000000100",
			7759 => "11111111111100010111101010100101",
			7760 => "00000000111110110111101010100101",
			7761 => "0000001110000000000000101000000100",
			7762 => "11111110000011100111101010100101",
			7763 => "00000000001100100111101010100101",
			7764 => "0000001100000000000100010100001000",
			7765 => "0000000111000000000000101000000100",
			7766 => "00000001111101100111101010100101",
			7767 => "00000011100011000111101010100101",
			7768 => "0000000011000000001101100000000100",
			7769 => "11111111001010010111101010100101",
			7770 => "00000001010000110111101010100101",
			7771 => "0000001011000000001100001000010000",
			7772 => "0000000101000000000110000100001000",
			7773 => "0000000110000000001101111100000100",
			7774 => "00000001011110010111101010100101",
			7775 => "11111110111001000111101010100101",
			7776 => "0000001100000000000000101000000100",
			7777 => "11111110000011110111101010100101",
			7778 => "00000000110010110111101010100101",
			7779 => "0000000010000000000101110000001000",
			7780 => "0000001101000000000001111100000100",
			7781 => "00000000100010100111101010100101",
			7782 => "11111110111000000111101010100101",
			7783 => "0000001000000000001011010100000100",
			7784 => "11111101111011110111101010100101",
			7785 => "11111111110110000111101010100101",
			7786 => "0000000000000000001111000101001000",
			7787 => "0000000100000000001000000100101100",
			7788 => "0000000000000000001101010000011000",
			7789 => "0000000100000000001011110000010000",
			7790 => "0000000110000000001010011000001000",
			7791 => "0000001010000000000111110100000100",
			7792 => "11111111010011110111101010100101",
			7793 => "00000000100000100111101010100101",
			7794 => "0000000100000000001000101000000100",
			7795 => "11111101100010000111101010100101",
			7796 => "00000000000000000111101010100101",
			7797 => "0000000000000000000111000100000100",
			7798 => "00000000011111110111101010100101",
			7799 => "11111101011011100111101010100101",
			7800 => "0000001100000000000000101000001000",
			7801 => "0000001010000000001000010100000100",
			7802 => "00000001101011100111101010100101",
			7803 => "11111101111000000111101010100101",
			7804 => "0000001011000000001110001100001000",
			7805 => "0000000001000000000111100100000100",
			7806 => "00000010010011100111101010100101",
			7807 => "00000000000000000111101010100101",
			7808 => "11111111001000110111101010100101",
			7809 => "0000000010000000001100010100001100",
			7810 => "0000000010000000000100101000000100",
			7811 => "11111111001001100111101010100101",
			7812 => "0000001000000000001100000100000100",
			7813 => "11111110010001010111101010100101",
			7814 => "11111100011001010111101010100101",
			7815 => "0000000100000000000110001100001100",
			7816 => "0000001000000000001001101000001000",
			7817 => "0000000000000000001101010000000100",
			7818 => "11111111111001110111101010100101",
			7819 => "00000001011000000111101010100101",
			7820 => "11111110111001110111101010100101",
			7821 => "11111110011100010111101010100101",
			7822 => "0000001000000000001001101000010100",
			7823 => "0000000100000000000110001100001100",
			7824 => "0000000001000000000010001100001000",
			7825 => "0000001010000000001000010100000100",
			7826 => "00000000100100000111101010100101",
			7827 => "00000001111011110111101010100101",
			7828 => "00000010001100110111101010100101",
			7829 => "0000000000000000000010111100000100",
			7830 => "11111110000110100111101010100101",
			7831 => "00000010101001010111101010100101",
			7832 => "0000000011000000000000001100000100",
			7833 => "11111110001001110111101010100101",
			7834 => "0000000010000000001110010000010000",
			7835 => "0000000110000000001010011000001000",
			7836 => "0000001101000000000001111100000100",
			7837 => "00000000101001110111101010100101",
			7838 => "00000001101001010111101010100101",
			7839 => "0000001100000000000100000000000100",
			7840 => "00000000111110110111101010100101",
			7841 => "11111110110101000111101010100101",
			7842 => "0000000110000000001100011000001000",
			7843 => "0000000101000000001100101100000100",
			7844 => "00000000101101010111101010100101",
			7845 => "11111111000000010111101010100101",
			7846 => "0000000101000000000100001000000100",
			7847 => "00000000101010000111101010100101",
			7848 => "00000000001001100111101010100101",
			7849 => "0000001100000000000100001010111000",
			7850 => "0000001111000000000010001001011000",
			7851 => "0000000011000000000100000000100000",
			7852 => "0000000111000000001100001000011100",
			7853 => "0000000001000000001110100000010000",
			7854 => "0000001001000000000010001100001000",
			7855 => "0000000011000000000100010100000100",
			7856 => "11111111110101100111110000011001",
			7857 => "00000000110000100111110000011001",
			7858 => "0000000010000000001110101000000100",
			7859 => "00000000001101000111110000011001",
			7860 => "11111111010010010111110000011001",
			7861 => "0000000011000000000000101000000100",
			7862 => "00000101011110000111110000011001",
			7863 => "0000001001000000000110101000000100",
			7864 => "11111110001111100111110000011001",
			7865 => "00000000111100100111110000011001",
			7866 => "11111110010000110111110000011001",
			7867 => "0000001001000000000110101000011100",
			7868 => "0000000011000000001101100000010000",
			7869 => "0000001111000000000001011000001000",
			7870 => "0000000011000000001000111000000100",
			7871 => "00000000111011010111110000011001",
			7872 => "00000010101000110111110000011001",
			7873 => "0000000010000000001001010000000100",
			7874 => "11111111011001110111110000011001",
			7875 => "00000000110011100111110000011001",
			7876 => "0000000001000000001110100000000100",
			7877 => "11111100111101010111110000011001",
			7878 => "0000001001000000000110101000000100",
			7879 => "00000010100110100111110000011001",
			7880 => "00000001010110000111110000011001",
			7881 => "0000000001000000001110100000001100",
			7882 => "0000001111000000001011011100001000",
			7883 => "0000001111000000000000011100000100",
			7884 => "11111110100011000111110000011001",
			7885 => "11111101000011100111110000011001",
			7886 => "11111111001111000111110000011001",
			7887 => "0000000110000000000001111000001000",
			7888 => "0000000101000000001110001100000100",
			7889 => "11111111110111110111110000011001",
			7890 => "11111110100100000111110000011001",
			7891 => "0000000000000000001011000100000100",
			7892 => "00000000100010100111110000011001",
			7893 => "11111110100101010111110000011001",
			7894 => "0000000011000000000101101100100000",
			7895 => "0000000011000000000101101100011000",
			7896 => "0000000011000000001100110000010000",
			7897 => "0000000111000000001011000100001000",
			7898 => "0000001010000000000110011000000100",
			7899 => "11111110000111110111110000011001",
			7900 => "00000000001000010111110000011001",
			7901 => "0000001100000000000111111000000100",
			7902 => "11111110001110000111110000011001",
			7903 => "11111111100111000111110000011001",
			7904 => "0000001100000000000100010100000100",
			7905 => "00000010000100000111110000011001",
			7906 => "11111111110100000111110000011001",
			7907 => "0000001111000000000101110100000100",
			7908 => "11111110110111100111110000011001",
			7909 => "11111101101101000111110000011001",
			7910 => "0000001000000000000010101000100000",
			7911 => "0000001001000000000110101000010000",
			7912 => "0000001111000000000111110000001000",
			7913 => "0000000111000000000100010100000100",
			7914 => "00000000101010010111110000011001",
			7915 => "00000011001100100111110000011001",
			7916 => "0000000110000000000100110100000100",
			7917 => "11111110100000010111110000011001",
			7918 => "00000001010000010111110000011001",
			7919 => "0000000011000000001100101100001000",
			7920 => "0000001001000000000111100100000100",
			7921 => "00000000000000000111110000011001",
			7922 => "11111110110000100111110000011001",
			7923 => "0000001001000000000111100100000100",
			7924 => "00000000010110100111110000011001",
			7925 => "00000000000000100111110000011001",
			7926 => "0000001010000000000110011100010000",
			7927 => "0000001100000000000000101000001000",
			7928 => "0000001111000000000001001000000100",
			7929 => "00000110000100110111110000011001",
			7930 => "00000001011010100111110000011001",
			7931 => "0000000100000000000011101100000100",
			7932 => "00000001011011100111110000011001",
			7933 => "11111110011111010111110000011001",
			7934 => "0000000000000000001011000100001000",
			7935 => "0000000100000000000010100100000100",
			7936 => "00000010011100010111110000011001",
			7937 => "11111110011000100111110000011001",
			7938 => "0000000111000000000000101000000100",
			7939 => "00000001111100110111110000011001",
			7940 => "11111111100000010111110000011001",
			7941 => "11111110011101000111110000011001",
			7942 => "0000000010000000001100010110110100",
			7943 => "0000000110000000001101011010000000",
			7944 => "0000000110000000001100011001000000",
			7945 => "0000000010000000000111111100100000",
			7946 => "0000000010000000000111111100010000",
			7947 => "0000000010000000000100101000001000",
			7948 => "0000000110000000001101111100000100",
			7949 => "11111111111010100111111100000111",
			7950 => "00000000001110100111111100000111",
			7951 => "0000001111000000000010001000000100",
			7952 => "00000001110010010111111100000111",
			7953 => "11111110010010100111111100000111",
			7954 => "0000000001000000001100110100001000",
			7955 => "0000001101000000001100110000000100",
			7956 => "00000011000000010111111100000111",
			7957 => "11111110100000000111111100000111",
			7958 => "0000000001000000001100110100000100",
			7959 => "00000010110010110111111100000111",
			7960 => "00000000100011000111111100000111",
			7961 => "0000000101000000000000001100010000",
			7962 => "0000000010000000001100010100001000",
			7963 => "0000001110000000001011000100000100",
			7964 => "11111111001101110111111100000111",
			7965 => "00000000000001100111111100000111",
			7966 => "0000001010000000001010110000000100",
			7967 => "00000000010101010111111100000111",
			7968 => "00000010100010000111111100000111",
			7969 => "0000001110000000000101101100001000",
			7970 => "0000001001000000000111100100000100",
			7971 => "00000001011110110111111100000111",
			7972 => "11111110000101110111111100000111",
			7973 => "0000000010000000000011001000000100",
			7974 => "00000000000101000111111100000111",
			7975 => "11111110010101100111111100000111",
			7976 => "0000000110000000001100011000100000",
			7977 => "0000001110000000001001110000010000",
			7978 => "0000001000000000000001110100001000",
			7979 => "0000000000000000000111111000000100",
			7980 => "00000000011001010111111100000111",
			7981 => "11111101111111110111111100000111",
			7982 => "0000000000000000000100010100000100",
			7983 => "00000011101001000111111100000111",
			7984 => "00000000011011110111111100000111",
			7985 => "0000001001000000001011101000001000",
			7986 => "0000001010000000000001010000000100",
			7987 => "00000001001001010111111100000111",
			7988 => "00000010100100010111111100000111",
			7989 => "0000001111000000000010110100000100",
			7990 => "11111111100011100111111100000111",
			7991 => "00000001111100110111111100000111",
			7992 => "0000001100000000000100000000010000",
			7993 => "0000001110000000001110001100001000",
			7994 => "0000001001000000000111100100000100",
			7995 => "00000000100010110111111100000111",
			7996 => "11111111001110110111111100000111",
			7997 => "0000000110000000001010011000000100",
			7998 => "00000001100011000111111100000111",
			7999 => "11111111110101100111111100000111",
			8000 => "0000001100000000001001110000001000",
			8001 => "0000001111000000000000110100000100",
			8002 => "11111110111010100111111100000111",
			8003 => "11111111111100000111111100000111",
			8004 => "0000001011000000001100101100000100",
			8005 => "00000011000110110111111100000111",
			8006 => "11111111111101000111111100000111",
			8007 => "0000000101000000000011100000100000",
			8008 => "0000000110000000001101011000010000",
			8009 => "0000000010000000001100010100001100",
			8010 => "0000000010000000000010011100000100",
			8011 => "11111111101101000111111100000111",
			8012 => "0000001110000000000110000100000100",
			8013 => "11111110010110010111111100000111",
			8014 => "11111101001110100111111100000111",
			8015 => "11111111011111010111111100000111",
			8016 => "0000000000000000000011111100000100",
			8017 => "11111101001111100111111100000111",
			8018 => "0000000000000000001110111100000100",
			8019 => "00000001101101000111111100000111",
			8020 => "0000001011000000001001110000000100",
			8021 => "00000000111000000111111100000111",
			8022 => "11111110000001010111111100000111",
			8023 => "0000001101000000000110100100001000",
			8024 => "0000001100000000000110000100000100",
			8025 => "00000100011010010111111100000111",
			8026 => "00000000000000000111111100000111",
			8027 => "0000001101000000001000011000000100",
			8028 => "11111111110101110111111100000111",
			8029 => "0000000101000000001000011000000100",
			8030 => "00000001100111010111111100000111",
			8031 => "00000000000000000111111100000111",
			8032 => "0000000110000000001100011001011000",
			8033 => "0000001100000000000111111000100100",
			8034 => "0000001010000000001010110000010000",
			8035 => "0000000010000000000110010000001000",
			8036 => "0000001000000000001111001000000100",
			8037 => "00000000000000000111111100000111",
			8038 => "00000010101011000111111100000111",
			8039 => "0000000100000000000011010100000100",
			8040 => "00000001100100010111111100000111",
			8041 => "11111110011010110111111100000111",
			8042 => "0000000010000000001110110100001100",
			8043 => "0000001011000000000100010100001000",
			8044 => "0000000010000000000010000000000100",
			8045 => "00000001110101110111111100000111",
			8046 => "11111110100111110111111100000111",
			8047 => "11111101101010000111111100000111",
			8048 => "0000001100000000001010000000000100",
			8049 => "11111111011001010111111100000111",
			8050 => "00000001111110110111111100000111",
			8051 => "0000000101000000000100001000011000",
			8052 => "0000001001000000001101101000010000",
			8053 => "0000001001000000000111100100001000",
			8054 => "0000000101000000001110001100000100",
			8055 => "11111111000101000111111100000111",
			8056 => "00000001110100110111111100000111",
			8057 => "0000001110000000001110001100000100",
			8058 => "11111101111010010111111100000111",
			8059 => "11111111110111010111111100000111",
			8060 => "0000000110000000001100011000000100",
			8061 => "11111110011011010111111100000111",
			8062 => "11111100000111110111111100000111",
			8063 => "0000000110000000001100011000001100",
			8064 => "0000000001000000000111100100000100",
			8065 => "11111101110100010111111100000111",
			8066 => "0000001110000000000011001000000100",
			8067 => "00000000101110010111111100000111",
			8068 => "11111111000001100111111100000111",
			8069 => "0000001111000000000001000000001000",
			8070 => "0000000100000000000000010100000100",
			8071 => "00000001100010000111111100000111",
			8072 => "11111110001110110111111100000111",
			8073 => "0000000010000000001001100000000100",
			8074 => "11111101010000110111111100000111",
			8075 => "11111111101010110111111100000111",
			8076 => "0000001001000000001011101001000000",
			8077 => "0000000100000000000100001100100000",
			8078 => "0000000101000000001010111100010000",
			8079 => "0000001001000000001101101000001000",
			8080 => "0000000101000000001101111000000100",
			8081 => "11111111111001010111111100000111",
			8082 => "00000010000010100111111100000111",
			8083 => "0000000001000000000010001100000100",
			8084 => "11111110001111100111111100000111",
			8085 => "11111111111000010111111100000111",
			8086 => "0000001111000000001101000100001000",
			8087 => "0000001100000000000100000000000100",
			8088 => "00000001111110110111111100000111",
			8089 => "11111111001011110111111100000111",
			8090 => "0000001110000000001101010100000100",
			8091 => "00000011000011110111111100000111",
			8092 => "00000001111111110111111100000111",
			8093 => "0000001011000000001100001000010000",
			8094 => "0000001010000000000110011100001000",
			8095 => "0000001110000000001000111000000100",
			8096 => "00000000010100100111111100000111",
			8097 => "00000011110001000111111100000111",
			8098 => "0000001111000000000010110100000100",
			8099 => "00000001001001000111111100000111",
			8100 => "11111110001001000111111100000111",
			8101 => "0000001011000000001000111100001000",
			8102 => "0000001001000000000110101000000100",
			8103 => "11111111110110100111111100000111",
			8104 => "11111110000111010111111100000111",
			8105 => "0000000110000000001101011000000100",
			8106 => "11111110111111100111111100000111",
			8107 => "00000000110001010111111100000111",
			8108 => "0000001100000000000100000000010100",
			8109 => "0000000110000000001101011000000100",
			8110 => "11111101101001010111111100000111",
			8111 => "0000000100000000001110111000001000",
			8112 => "0000001001000000001111001100000100",
			8113 => "00000001111101100111111100000111",
			8114 => "11111110111111110111111100000111",
			8115 => "0000001010000000000101000100000100",
			8116 => "11111101101111010111111100000111",
			8117 => "00000000000000000111111100000111",
			8118 => "0000001100000000000100000000001000",
			8119 => "0000000110000000001111000000000100",
			8120 => "00000010100000010111111100000111",
			8121 => "11111110110111010111111100000111",
			8122 => "0000001111000000001101000100001000",
			8123 => "0000000110000000001001100100000100",
			8124 => "11111101101111010111111100000111",
			8125 => "00000001011110000111111100000111",
			8126 => "0000000110000000001011001100000100",
			8127 => "00000000100110000111111100000111",
			8128 => "11111111011010110111111100000111",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(2792, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(5598, initial_addr_3'length));
	end generate gen_rom_14;

	gen_rom_15: if SELECT_ROM = 15 generate
		bank <= (
			0 => "00000000000000000000000000000101",
			1 => "00000000000000000000000000001001",
			2 => "00000000000000000000000000001101",
			3 => "00000000000000000000000000010001",
			4 => "00000000000000000000000000010101",
			5 => "00000000000000000000000000011001",
			6 => "00000000000000000000000000011101",
			7 => "00000000000000000000000000100001",
			8 => "00000000000000000000000000100101",
			9 => "00000000000000000000000000101001",
			10 => "00000000000000000000000000101101",
			11 => "00000000000000000000000000110001",
			12 => "00000000000000000000000000110101",
			13 => "00000000000000000000000000111001",
			14 => "00000000000000000000000000111101",
			15 => "00000000000000000000000001000001",
			16 => "00000000000000000000000001000101",
			17 => "00000000000000000000000001001001",
			18 => "00000000000000000000000001001101",
			19 => "0000001011000000001101010100000100",
			20 => "00000000000000000000000001011001",
			21 => "11111111110010000000000001011001",
			22 => "0000000111000000001110001100000100",
			23 => "00000000000000010000000001100101",
			24 => "00000000000000000000000001100101",
			25 => "0000001100000000001010000000000100",
			26 => "00000000000000000000000001110001",
			27 => "11111111111111100000000001110001",
			28 => "0000001100000000001010000000000100",
			29 => "00000000000000000000000010000101",
			30 => "0000001010000000000000001000000100",
			31 => "00000000000000000000000010000101",
			32 => "11111111110101000000000010000101",
			33 => "0000000111000000001110001100001000",
			34 => "0000001011000000000000111000000100",
			35 => "00000000000000000000000010011001",
			36 => "00000000000011100000000010011001",
			37 => "00000000000000000000000010011001",
			38 => "0000000110000000000001000100000100",
			39 => "00000000000000000000000010101101",
			40 => "0000000110000000001010011000000100",
			41 => "11111111111011110000000010101101",
			42 => "00000000000000000000000010101101",
			43 => "0000000110000000001101111100001000",
			44 => "0000000110000000001101011100000100",
			45 => "00000000000000000000000011000001",
			46 => "00000000000001000000000011000001",
			47 => "00000000000000000000000011000001",
			48 => "0000000001000000001110100000001000",
			49 => "0000001001000000001100100000000100",
			50 => "00000000000000000000000011010101",
			51 => "00000000000000000000000011010101",
			52 => "11111111111011110000000011010101",
			53 => "0000000110000000001110010100000100",
			54 => "00000000000000000000000011101001",
			55 => "0000000110000000001111000000000100",
			56 => "11111111111100110000000011101001",
			57 => "00000000000000000000000011101001",
			58 => "0000000110000000000001111000000100",
			59 => "00000000000000000000000100000101",
			60 => "0000000110000000001010011000001000",
			61 => "0000000100000000001101000000000100",
			62 => "11111111100010110000000100000101",
			63 => "00000000000000000000000100000101",
			64 => "00000000000000000000000100000101",
			65 => "0000000111000000001110001100001100",
			66 => "0000001111000000001001001000000100",
			67 => "00000000000000000000000100100001",
			68 => "0000001100000000001100110000000100",
			69 => "00000000001101000000000100100001",
			70 => "00000000000000000000000100100001",
			71 => "00000000000000000000000100100001",
			72 => "0000000110000000000001111000001100",
			73 => "0000000110000000001101011100000100",
			74 => "00000000000000000000000100111101",
			75 => "0000000110000000001011111100000100",
			76 => "00000000001000000000000100111101",
			77 => "00000000000000000000000100111101",
			78 => "11111111110100110000000100111101",
			79 => "0000000111000000001110001100001100",
			80 => "0000001111000000000100011000000100",
			81 => "00000000000000000000000101011001",
			82 => "0000000001000000001011101000000100",
			83 => "00000000010000100000000101011001",
			84 => "00000000000000000000000101011001",
			85 => "00000000000000000000000101011001",
			86 => "0000000110000000001101111100001100",
			87 => "0000001010000000001001100100000100",
			88 => "00000000000000000000000101111101",
			89 => "0000001010000000000011101000000100",
			90 => "00000000010000100000000101111101",
			91 => "00000000000000000000000101111101",
			92 => "0000000110000000001001100100000100",
			93 => "11111111100101010000000101111101",
			94 => "00000000000000000000000101111101",
			95 => "0000000001000000000110000000001100",
			96 => "0000000001000000001110011100000100",
			97 => "00000000000000000000000110100001",
			98 => "0000000010000000001010010100000100",
			99 => "00000000000000000000000110100001",
			100 => "00000000000101010000000110100001",
			101 => "0000000010000000001100010100000100",
			102 => "11111111111011000000000110100001",
			103 => "00000000000000000000000110100001",
			104 => "0000000001000000000000011000001100",
			105 => "0000001100000000000111111000001000",
			106 => "0000001111000000001010111100000100",
			107 => "00000000000000000000000111001101",
			108 => "00000000010101110000000111001101",
			109 => "00000000000000000000000111001101",
			110 => "0000000000000000001001101000000100",
			111 => "00000000000000000000000111001101",
			112 => "0000000110000000001011111100000100",
			113 => "00000000000000000000000111001101",
			114 => "11111111001111000000000111001101",
			115 => "0000000111000000001110001100010000",
			116 => "0000001010000000001000100100001100",
			117 => "0000001101000000000100000000000100",
			118 => "00000000000000000000000111110001",
			119 => "0000001000000000000000001000000100",
			120 => "00000000000000000000000111110001",
			121 => "00000000011110100000000111110001",
			122 => "00000000000000000000000111110001",
			123 => "11111111100110110000000111110001",
			124 => "0000000110000000000001000100000100",
			125 => "00000000000000000000001000010101",
			126 => "0000001100000000000000110000000100",
			127 => "00000000000000000000001000010101",
			128 => "0000001100000000001110001100001000",
			129 => "0000000110000000001101111100000100",
			130 => "00000000000000000000001000010101",
			131 => "11111111101111100000001000010101",
			132 => "00000000000000000000001000010101",
			133 => "0000001011000000001010111000010000",
			134 => "0000001111000000001110110000000100",
			135 => "00000000000000000000001000111001",
			136 => "0000001100000000001100110000001000",
			137 => "0000000111000000001110001100000100",
			138 => "00000000010001000000001000111001",
			139 => "00000000000000000000001000111001",
			140 => "00000000000000000000001000111001",
			141 => "00000000000000000000001000111001",
			142 => "0000000111000000001110001100010000",
			143 => "0000001111000000001010111100000100",
			144 => "00000000000000000000001001011101",
			145 => "0000001010000000001001100100000100",
			146 => "00000000000000000000001001011101",
			147 => "0000001100000000001100110000000100",
			148 => "00000000010000010000001001011101",
			149 => "00000000000000000000001001011101",
			150 => "00000000000000000000001001011101",
			151 => "0000001111000000001010111100000100",
			152 => "00000000000000000000001010000001",
			153 => "0000001100000000000100001000001100",
			154 => "0000001111000000001100111000001000",
			155 => "0000000111000000001110110000000100",
			156 => "00000000001000010000001010000001",
			157 => "00000000000000000000001010000001",
			158 => "00000000000000000000001010000001",
			159 => "00000000000000000000001010000001",
			160 => "0000000111000000000110000100010000",
			161 => "0000000110000000001101111100001100",
			162 => "0000000110000000001001011000000100",
			163 => "00000000000000000000001010101101",
			164 => "0000001011000000000000111000000100",
			165 => "00000000000000000000001010101101",
			166 => "00000000001110100000001010101101",
			167 => "00000000000000000000001010101101",
			168 => "0000001011000000001001110100000100",
			169 => "11111111110101110000001010101101",
			170 => "00000000000000000000001010101101",
			171 => "0000000010000000001110010000001100",
			172 => "0000000001000000000000011000000100",
			173 => "00000000000000000000001011100001",
			174 => "0000001100000000000000111000000100",
			175 => "00000000000000000000001011100001",
			176 => "11111111110100010000001011100001",
			177 => "0000000111000000001110001100001100",
			178 => "0000000001000000001011101000001000",
			179 => "0000001100000000000011011100000100",
			180 => "00000000100111010000001011100001",
			181 => "00000000000000000000001011100001",
			182 => "00000000000000000000001011100001",
			183 => "00000000000000000000001011100001",
			184 => "0000000001000000001110100000010000",
			185 => "0000001001000000001100100000000100",
			186 => "00000000000000000000001100010101",
			187 => "0000000101000000000100000000000100",
			188 => "00000000000000000000001100010101",
			189 => "0000000111000000000000101000000100",
			190 => "00000000001101110000001100010101",
			191 => "00000000000000000000001100010101",
			192 => "0000000110000000001010011000001000",
			193 => "0000000001000000001110100000000100",
			194 => "00000000000000000000001100010101",
			195 => "11111111101001010000001100010101",
			196 => "00000000000000000000001100010101",
			197 => "0000000111000000001110001100011000",
			198 => "0000001111000000000101100100001100",
			199 => "0000000110000000000001000100000100",
			200 => "00000000000000000000001101010001",
			201 => "0000000001000000001100100000000100",
			202 => "00000000000000000000001101010001",
			203 => "11111111110011000000001101010001",
			204 => "0000000001000000001011101000001000",
			205 => "0000001010000000001000100100000100",
			206 => "00000000100011110000001101010001",
			207 => "00000000000000000000001101010001",
			208 => "00000000000000000000001101010001",
			209 => "0000000110000000001001100100000100",
			210 => "11111111110110000000001101010001",
			211 => "00000000000000000000001101010001",
			212 => "0000000111000000001110001100010100",
			213 => "0000001111000000001010111100000100",
			214 => "00000000000000000000001101111101",
			215 => "0000001010000000001001100100000100",
			216 => "00000000000000000000001101111101",
			217 => "0000001100000000001100110000001000",
			218 => "0000001011000000000000111000000100",
			219 => "00000000000000000000001101111101",
			220 => "00000000001111000000001101111101",
			221 => "00000000000000000000001101111101",
			222 => "00000000000000000000001101111101",
			223 => "0000001100000000001010000000000100",
			224 => "00000000000000000000001110101001",
			225 => "0000000110000000000101011100000100",
			226 => "00000000000000000000001110101001",
			227 => "0000000110000000001001100100001100",
			228 => "0000000111000000001010000000000100",
			229 => "00000000000000000000001110101001",
			230 => "0000000110000000001011111100000100",
			231 => "00000000000000000000001110101001",
			232 => "11111111110110100000001110101001",
			233 => "00000000000000000000001110101001",
			234 => "0000001100000000001010000000010100",
			235 => "0000000010000000000001001000000100",
			236 => "00000000000000000000001111100101",
			237 => "0000000001000000001110100000001100",
			238 => "0000001001000000001100100000000100",
			239 => "00000000000000000000001111100101",
			240 => "0000001011000000000000111000000100",
			241 => "00000000000000000000001111100101",
			242 => "00000000010111010000001111100101",
			243 => "00000000000000000000001111100101",
			244 => "0000000110000000001010011000001000",
			245 => "0000000110000000000001111000000100",
			246 => "00000000000000000000001111100101",
			247 => "11111111011100010000001111100101",
			248 => "00000000000000000000001111100101",
			249 => "0000001100000000001010000000010100",
			250 => "0000000001000000001110100000010000",
			251 => "0000001101000000000000101000000100",
			252 => "00000000000000000000010000100001",
			253 => "0000001001000000001100100000000100",
			254 => "00000000000000000000010000100001",
			255 => "0000000111000000000100010100000100",
			256 => "00000000001011110000010000100001",
			257 => "00000000000000000000010000100001",
			258 => "00000000000000000000010000100001",
			259 => "0000000111000000000111001000001000",
			260 => "0000000001000000001110100000000100",
			261 => "00000000000000000000010000100001",
			262 => "11111111110000010000010000100001",
			263 => "00000000000000000000010000100001",
			264 => "0000000001000000000110000000010000",
			265 => "0000001100000000000100000000001100",
			266 => "0000001001000000001100100000000100",
			267 => "00000000000000000000010001100101",
			268 => "0000000001000000001110011100000100",
			269 => "00000000000000000000010001100101",
			270 => "00000000000101110000010001100101",
			271 => "00000000000000000000010001100101",
			272 => "0000001100000000001100110000010000",
			273 => "0000000110000000001010011000001100",
			274 => "0000001100000000001010000000000100",
			275 => "00000000000000000000010001100101",
			276 => "0000000110000000001001011000000100",
			277 => "00000000000000000000010001100101",
			278 => "11111111101111000000010001100101",
			279 => "00000000000000000000010001100101",
			280 => "00000000000000000000010001100101",
			281 => "0000001001000000000010001100001100",
			282 => "0000000011000000001010101100000100",
			283 => "00000000000000000000010010110001",
			284 => "0000000111000000001100001000000100",
			285 => "00000000100010110000010010110001",
			286 => "00000000000000000000010010110001",
			287 => "0000001110000000000101001000010000",
			288 => "0000001010000000000000001000000100",
			289 => "00000000000000000000010010110001",
			290 => "0000001100000000000000111000000100",
			291 => "00000000000000000000010010110001",
			292 => "0000000110000000001011111100000100",
			293 => "00000000000000000000010010110001",
			294 => "11111111000111000000010010110001",
			295 => "0000001110000000001001010000000100",
			296 => "00000000000110000000010010110001",
			297 => "0000000010000000001100111000000100",
			298 => "11111111111000010000010010110001",
			299 => "00000000000000000000010010110001",
			300 => "0000001100000000001010000000010100",
			301 => "0000000010000000001010010100000100",
			302 => "00000000000000000000010011111101",
			303 => "0000001011000000001011000100001100",
			304 => "0000001011000000000000111000000100",
			305 => "00000000000000000000010011111101",
			306 => "0000000111000000000100010100000100",
			307 => "00000000010101000000010011111101",
			308 => "00000000000000000000010011111101",
			309 => "00000000000000000000010011111101",
			310 => "0000000010000000001100010100001000",
			311 => "0000000111000000001010000000000100",
			312 => "00000000000000000000010011111101",
			313 => "11111111110010110000010011111101",
			314 => "0000000111000000001110001100001000",
			315 => "0000000111000000000101101100000100",
			316 => "00000000000000000000010011111101",
			317 => "00000000001010000000010011111101",
			318 => "00000000000000000000010011111101",
			319 => "0000001000000000000101000100011000",
			320 => "0000001110000000000010111100000100",
			321 => "00000000000000000000010101001001",
			322 => "0000001110000000001001010000001100",
			323 => "0000001010000000000011101000001000",
			324 => "0000000000000000001010110000000100",
			325 => "00000000000000000000010101001001",
			326 => "00000000011101100000010101001001",
			327 => "00000000000000000000010101001001",
			328 => "0000001000000000001010110000000100",
			329 => "11111111111101100000010101001001",
			330 => "00000000000000000000010101001001",
			331 => "0000001110000000000111010100001100",
			332 => "0000001110000000001000110000000100",
			333 => "00000000000000000000010101001001",
			334 => "0000001010000000000111110100000100",
			335 => "00000000000000000000010101001001",
			336 => "11111111100101110000010101001001",
			337 => "00000000000000000000010101001001",
			338 => "0000000001000000001110100000011000",
			339 => "0000000010000000000100101000010000",
			340 => "0000000110000000000001000100001000",
			341 => "0000000011000000000000111000000100",
			342 => "00000000000000000000010110100101",
			343 => "00000000011001010000010110100101",
			344 => "0000001110000000001110111100000100",
			345 => "11111111100101110000010110100101",
			346 => "00000000000000000000010110100101",
			347 => "0000001100000000000100010100000100",
			348 => "00000000110111100000010110100101",
			349 => "00000000000000000000010110100101",
			350 => "0000001101000000000010001000001000",
			351 => "0000001010000000000111101100000100",
			352 => "00000000000000000000010110100101",
			353 => "11111110110111100000010110100101",
			354 => "0000001001000000001011001100001100",
			355 => "0000001100000000000100001000001000",
			356 => "0000001101000000001110101100000100",
			357 => "00000000011000110000010110100101",
			358 => "00000000000000000000010110100101",
			359 => "00000000000000000000010110100101",
			360 => "11111111110010000000010110100101",
			361 => "0000000001000000000000011000010100",
			362 => "0000001100000000000111111000010000",
			363 => "0000001001000000001100100000000100",
			364 => "00000000000000000000010111110001",
			365 => "0000001011000000000000111000000100",
			366 => "00000000000000000000010111110001",
			367 => "0000000001000000001110011100000100",
			368 => "00000000000000000000010111110001",
			369 => "00000000010001010000010111110001",
			370 => "00000000000000000000010111110001",
			371 => "0000000010000000001011111000010000",
			372 => "0000001100000000001100110000001100",
			373 => "0000001000000000001001000100000100",
			374 => "00000000000000000000010111110001",
			375 => "0000001100000000000000111000000100",
			376 => "00000000000000000000010111110001",
			377 => "11111111100010010000010111110001",
			378 => "00000000000000000000010111110001",
			379 => "00000000000000000000010111110001",
			380 => "0000000110000000001101111100100000",
			381 => "0000001111000000000010001000010100",
			382 => "0000000110000000000001000100001100",
			383 => "0000000001000000000110000000001000",
			384 => "0000000001000000001110011100000100",
			385 => "00000000000000000000011001001101",
			386 => "00000000001101110000011001001101",
			387 => "00000000000000000000011001001101",
			388 => "0000000001000000001100100000000100",
			389 => "00000000000000000000011001001101",
			390 => "11111111100101100000011001001101",
			391 => "0000001011000000001101010100001000",
			392 => "0000001010000000000011101000000100",
			393 => "00000000100111110000011001001101",
			394 => "00000000000000000000011001001101",
			395 => "00000000000000000000011001001101",
			396 => "0000001010000000001000110000001100",
			397 => "0000001111000000001000001100001000",
			398 => "0000000100000000000110111100000100",
			399 => "00000000000000000000011001001101",
			400 => "11111111001010110000011001001101",
			401 => "00000000000000000000011001001101",
			402 => "00000000000000000000011001001101",
			403 => "0000001100000000000100001000011000",
			404 => "0000001111000000001110110000000100",
			405 => "00000000000000000000011010000001",
			406 => "0000001010000000001000100100010000",
			407 => "0000000011000000000010000000001100",
			408 => "0000001010000000001001100100000100",
			409 => "00000000000000000000011010000001",
			410 => "0000001101000000001110101100000100",
			411 => "00000000010010110000011010000001",
			412 => "00000000000000000000011010000001",
			413 => "00000000000000000000011010000001",
			414 => "00000000000000000000011010000001",
			415 => "00000000000000000000011010000001",
			416 => "0000000110000000001110010100010100",
			417 => "0000001001000000001001111000001000",
			418 => "0000000010000000000101110100000100",
			419 => "11010011100111100000011011100101",
			420 => "11111000111110000000011011100101",
			421 => "0000000001000000001110100000001000",
			422 => "0000001110000000000000110000000100",
			423 => "11001000010110000000011011100101",
			424 => "11011111011101100000011011100101",
			425 => "11000111111110010000011011100101",
			426 => "0000000110000000000111101000001000",
			427 => "0000000010000000001110010000000100",
			428 => "11001000000001110000011011100101",
			429 => "11110101011101110000011011100101",
			430 => "0000001100000000000000110000001000",
			431 => "0000000010000000001100010100000100",
			432 => "11000111111110010000011011100101",
			433 => "11110011010000010000011011100101",
			434 => "0000000111000000001110111100001100",
			435 => "0000001101000000001000111100000100",
			436 => "11000111111111010000011011100101",
			437 => "0000001011000000001110111100000100",
			438 => "11010011111001110000011011100101",
			439 => "11001000001110110000011011100101",
			440 => "11000111111110110000011011100101",
			441 => "0000000010000000001100010100010100",
			442 => "0000000110000000000001111000010000",
			443 => "0000000010000000000001101000000100",
			444 => "00000000000000000000011100111001",
			445 => "0000000110000000001011111100001000",
			446 => "0000000001000000001110100000000100",
			447 => "00000000010111000000011100111001",
			448 => "00000000000000000000011100111001",
			449 => "00000000000000000000011100111001",
			450 => "11111111011001000000011100111001",
			451 => "0000000001000000001101011100010100",
			452 => "0000001100000000000100001000010000",
			453 => "0000001001000000001100100000000100",
			454 => "00000000000000000000011100111001",
			455 => "0000000100000000001101001100001000",
			456 => "0000000010000000000011000000000100",
			457 => "00000000101111100000011100111001",
			458 => "00000000000000000000011100111001",
			459 => "00000000000000000000011100111001",
			460 => "00000000000000000000011100111001",
			461 => "00000000000000000000011100111001",
			462 => "0000000001000000000110000000010000",
			463 => "0000001111000000001110110000001000",
			464 => "0000000111000000000000110000000100",
			465 => "00000000000000000000011110010101",
			466 => "11111111110111010000011110010101",
			467 => "0000000111000000001100001000000100",
			468 => "00000000111111010000011110010101",
			469 => "00000000000000000000011110010101",
			470 => "0000000111000000001101100000001000",
			471 => "0000000001000000001110100000000100",
			472 => "00000000000000000000011110010101",
			473 => "11111110101011010000011110010101",
			474 => "0000000111000000000111001000010100",
			475 => "0000001000000000000001110000010000",
			476 => "0000000001000000001001011000001100",
			477 => "0000001111000000001010010100000100",
			478 => "00000000000000000000011110010101",
			479 => "0000001000000000000111110100000100",
			480 => "00000000000000000000011110010101",
			481 => "00000000101100110000011110010101",
			482 => "00000000000000000000011110010101",
			483 => "00000000000000000000011110010101",
			484 => "11111111011110100000011110010101",
			485 => "0000001000000000000101000100100000",
			486 => "0000000011000000000010000000011100",
			487 => "0000000010000000001100010100010100",
			488 => "0000000001000000001110100000001100",
			489 => "0000001110000000000010111100000100",
			490 => "00000000000000000000100000000001",
			491 => "0000001000000000001100011100000100",
			492 => "00000000100110100000100000000001",
			493 => "00000000000000000000100000000001",
			494 => "0000001000000000000111110100000100",
			495 => "00000000000000000000100000000001",
			496 => "11111111100111100000100000000001",
			497 => "0000000001000000001011111100000100",
			498 => "00000000111011000000100000000001",
			499 => "00000000000000000000100000000001",
			500 => "11111111111001000000100000000001",
			501 => "0000001001000000001100110100001100",
			502 => "0000001100000000001010000000001000",
			503 => "0000001101000000000000101000000100",
			504 => "00000000000000000000100000000001",
			505 => "00000000001001000000100000000001",
			506 => "00000000000000000000100000000001",
			507 => "0000000010000000001100010000001000",
			508 => "0000000101000000001000111100000100",
			509 => "00000000000000000000100000000001",
			510 => "11111110110111100000100000000001",
			511 => "00000000000000000000100000000001",
			512 => "0000000001000000000000011000010100",
			513 => "0000001111000000001011000000001000",
			514 => "0000001100000000000000110000000100",
			515 => "00000000000000000000100001101101",
			516 => "11111111111011010000100001101101",
			517 => "0000001101000000000001111100001000",
			518 => "0000001001000000001100110100000100",
			519 => "00000001010010100000100001101101",
			520 => "00000000000000000000100001101101",
			521 => "00000000000000000000100001101101",
			522 => "0000000000000000000111000000011100",
			523 => "0000000001000000001101011100011000",
			524 => "0000001111000000000011001000001100",
			525 => "0000000001000000001110100000001000",
			526 => "0000001110000000000000101000000100",
			527 => "00000000000000000000100001101101",
			528 => "00000000110011100000100001101101",
			529 => "11111111000100000000100001101101",
			530 => "0000001001000000001011001100001000",
			531 => "0000000101000000000001001000000100",
			532 => "00000001001011000000100001101101",
			533 => "00000000000000000000100001101101",
			534 => "00000000000000000000100001101101",
			535 => "11111111010010010000100001101101",
			536 => "0000000110000000001011111100000100",
			537 => "00000000000000000000100001101101",
			538 => "11111110100110010000100001101101",
			539 => "0000000001000000000110000000011000",
			540 => "0000001111000000001110110000000100",
			541 => "00000000000000000000100011011001",
			542 => "0000001101000000000001111100010000",
			543 => "0000001101000000000100000000000100",
			544 => "00000000000000000000100011011001",
			545 => "0000001100000000000100010100001000",
			546 => "0000001100000000000011111100000100",
			547 => "00000000000000000000100011011001",
			548 => "00000000101101110000100011011001",
			549 => "00000000000000000000100011011001",
			550 => "00000000000000000000100011011001",
			551 => "0000001001000000001100011000001100",
			552 => "0000000111000000000111111000000100",
			553 => "00000000000000000000100011011001",
			554 => "0000000110000000001001011000000100",
			555 => "00000000000000000000100011011001",
			556 => "11111110111110110000100011011001",
			557 => "0000000001000000001101011100010000",
			558 => "0000000111000000001110110000001100",
			559 => "0000001100000000001000111000000100",
			560 => "00000000000000000000100011011001",
			561 => "0000000101000000001001010100000100",
			562 => "00000000010100110000100011011001",
			563 => "00000000000000000000100011011001",
			564 => "00000000000000000000100011011001",
			565 => "00000000000000000000100011011001",
			566 => "0000000001000000000110000000011000",
			567 => "0000001111000000001011000000001100",
			568 => "0000001100000000000000110000000100",
			569 => "00000000000000000000100101010101",
			570 => "0000001110000000001100011100000100",
			571 => "00000000000000000000100101010101",
			572 => "11111111101011000000100101010101",
			573 => "0000001101000000000001111100001000",
			574 => "0000000001000000000000011000000100",
			575 => "00000001010100100000100101010101",
			576 => "00000000000010100000100101010101",
			577 => "00000000000000000000100101010101",
			578 => "0000000000000000000111000000011100",
			579 => "0000000001000000001101011100011000",
			580 => "0000001111000000000011001000001100",
			581 => "0000000001000000001110100000001000",
			582 => "0000000011000000000110000100000100",
			583 => "00000000000000000000100101010101",
			584 => "00000000011010110000100101010101",
			585 => "11111111000110110000100101010101",
			586 => "0000001001000000001011001100001000",
			587 => "0000000101000000000001001000000100",
			588 => "00000001000110010000100101010101",
			589 => "00000000000000000000100101010101",
			590 => "00000000000000000000100101010101",
			591 => "11111111010101000000100101010101",
			592 => "0000001001000000000010001100000100",
			593 => "00000000000000000000100101010101",
			594 => "0000001011000000001110111100000100",
			595 => "00000000000000000000100101010101",
			596 => "11111110100111010000100101010101",
			597 => "0000001010000000001000100100100000",
			598 => "0000001001000000001011001100011100",
			599 => "0000001111000000001011011100001000",
			600 => "0000000001000000000110000000000100",
			601 => "00000000100111110000100111000001",
			602 => "11111111010111010000100111000001",
			603 => "0000001100000000000100001000010000",
			604 => "0000001000000000000011101000000100",
			605 => "00000000000000000000100111000001",
			606 => "0000000101000000001010010100001000",
			607 => "0000001000000000000101000100000100",
			608 => "00000000111111010000100111000001",
			609 => "00000000000000000000100111000001",
			610 => "00000000000000000000100111000001",
			611 => "00000000000000000000100111000001",
			612 => "11111111011100100000100111000001",
			613 => "0000000110000000000001111000010000",
			614 => "0000000100000000001111100000000100",
			615 => "11111111111011010000100111000001",
			616 => "0000000111000000000100010100001000",
			617 => "0000000011000000000001110100000100",
			618 => "00000000000000000000100111000001",
			619 => "00000000110001000000100111000001",
			620 => "00000000000000000000100111000001",
			621 => "0000001100000000000000111000000100",
			622 => "00000000000000000000100111000001",
			623 => "11111110100101110000100111000001",
			624 => "0000000110000000000001111000100100",
			625 => "0000000010000000000101001000011100",
			626 => "0000001010000000000011101000010100",
			627 => "0000001111000000001110110000000100",
			628 => "11111111011111100000101001000101",
			629 => "0000000111000000000110000100001100",
			630 => "0000000000000000000011101000000100",
			631 => "00000000000000000000101001000101",
			632 => "0000001010000000000010101100000100",
			633 => "00000001010100110000101001000101",
			634 => "00000000000000000000101001000101",
			635 => "00000000000000000000101001000101",
			636 => "0000000110000000001011111100000100",
			637 => "00000000000000000000101001000101",
			638 => "11111110101110000000101001000101",
			639 => "0000000111000000000000101000000100",
			640 => "00000001011001010000101001000101",
			641 => "11111111111010110000101001000101",
			642 => "0000000000000000000111000000010100",
			643 => "0000000101000000000110110100001000",
			644 => "0000001111000000000011001000000100",
			645 => "11111111001101100000101001000101",
			646 => "00000000111101100000101001000101",
			647 => "0000001000000000000001110000000100",
			648 => "11111110101001100000101001000101",
			649 => "0000000011000000000010010100000100",
			650 => "00000000011001110000101001000101",
			651 => "00000000000000000000101001000101",
			652 => "0000001100000000000000111000000100",
			653 => "00000000000000000000101001000101",
			654 => "0000000111000000001110111100000100",
			655 => "00000000000000000000101001000101",
			656 => "11111110011101010000101001000101",
			657 => "0000001100000000001010000000010000",
			658 => "0000000010000000000100101000001000",
			659 => "0000000110000000001110010100000100",
			660 => "00000001000111100000101010111001",
			661 => "11111111000101000000101010111001",
			662 => "0000000001000000001110100000000100",
			663 => "00000001101100110000101010111001",
			664 => "00000000000000000000101010111001",
			665 => "0000001000000000000001110000100000",
			666 => "0000001100000000000000001100011100",
			667 => "0000001010000000001000100100010100",
			668 => "0000001001000000001001111000001000",
			669 => "0000001110000000000011111100000100",
			670 => "00000000000000000000101010111001",
			671 => "00000000111100110000101010111001",
			672 => "0000000000000000001001101000001000",
			673 => "0000000010000000000101110000000100",
			674 => "00000000000000000000101010111001",
			675 => "00000000110001110000101010111001",
			676 => "11111110101100100000101010111001",
			677 => "0000001110000000000100101000000100",
			678 => "00000000000000000000101010111001",
			679 => "00000001011001110000101010111001",
			680 => "11111110111001000000101010111001",
			681 => "0000000110000000001011111100000100",
			682 => "00000000000000000000101010111001",
			683 => "0000000111000000001010000000000100",
			684 => "00000000000000000000101010111001",
			685 => "11111110011110100000101010111001",
			686 => "0000000110000000000111101000101000",
			687 => "0000000001000000000110000000010100",
			688 => "0000001111000000001010111100000100",
			689 => "11111110111111010000101101001101",
			690 => "0000000110000000001110010100000100",
			691 => "00000001101110110000101101001101",
			692 => "0000001100000000000000110000000100",
			693 => "00000001100101010000101101001101",
			694 => "0000000110000000000111101000000100",
			695 => "11111111011011010000101101001101",
			696 => "00000001000101010000101101001101",
			697 => "0000001111000000001011011100001100",
			698 => "0000000110000000001001011000001000",
			699 => "0000001111000000001110110000000100",
			700 => "11111111010000100000101101001101",
			701 => "00000001110000110000101101001101",
			702 => "11111110011010000000101101001101",
			703 => "0000000001000000001100110100000100",
			704 => "00000010001010010000101101001101",
			705 => "11111110111100000000101101001101",
			706 => "0000001100000000001010000000010000",
			707 => "0000000010000000000110010000001100",
			708 => "0000000010000000000011001000000100",
			709 => "11111110011100000000101101001101",
			710 => "0000001111000000000010001000000100",
			711 => "00000001010100100000101101001101",
			712 => "11111110111001000000101101001101",
			713 => "00000010100011010000101101001101",
			714 => "0000000000000000000111000000010000",
			715 => "0000001100000000000000001100001100",
			716 => "0000000010000000000010000100000100",
			717 => "11111110100101100000101101001101",
			718 => "0000001000000000000110011100000100",
			719 => "00000000111101000000101101001101",
			720 => "00000100010000000000101101001101",
			721 => "11111110011010010000101101001101",
			722 => "11111110011001010000101101001101",
			723 => "0000000110000000001110010100010000",
			724 => "0000001111000000000111001000001000",
			725 => "0000000000000000000001110100000100",
			726 => "11111111000001000000101111010001",
			727 => "00000000000000000000101111010001",
			728 => "0000001001000000000110101000000100",
			729 => "00000001100100010000101111010001",
			730 => "11111111010001100000101111010001",
			731 => "0000000000000000000111000000011000",
			732 => "0000000111000000000111001000010100",
			733 => "0000000111000000000101101100000100",
			734 => "11111111000010000000101111010001",
			735 => "0000000111000000001110001100000100",
			736 => "00000010010110110000101111010001",
			737 => "0000000111000000000111001000000100",
			738 => "11111110100110100000101111010001",
			739 => "0000000001000000001001011000000100",
			740 => "00000001110110110000101111010001",
			741 => "00000000000000000000101111010001",
			742 => "11111110100001010000101111010001",
			743 => "0000001011000000001110111100001100",
			744 => "0000000010000000001110010000000100",
			745 => "11111110101101000000101111010001",
			746 => "0000000100000000000010010000000100",
			747 => "00000000000000000000101111010001",
			748 => "00000001010110000000101111010001",
			749 => "0000001000000000000101000100000100",
			750 => "00000000000000000000101111010001",
			751 => "0000000101000000000100000000000100",
			752 => "00000000000000000000101111010001",
			753 => "0000001110000000000001010100000100",
			754 => "00000000000000000000101111010001",
			755 => "11111110011010010000101111010001",
			756 => "0000000110000000001110010100010100",
			757 => "0000001111000000000111001000001000",
			758 => "0000001100000000001010000000000100",
			759 => "00000000000000000000110001011101",
			760 => "11111111000001110000110001011101",
			761 => "0000001001000000000110101000001000",
			762 => "0000000001000000001110100000000100",
			763 => "00000001100110010000110001011101",
			764 => "00000000011011110000110001011101",
			765 => "11111111010101110000110001011101",
			766 => "0000000000000000000111000000011000",
			767 => "0000001100000000000000001100010100",
			768 => "0000001100000000001000111000000100",
			769 => "11111110111010000000110001011101",
			770 => "0000000111000000001110001100000100",
			771 => "00000010000111110000110001011101",
			772 => "0000000111000000000111001000000100",
			773 => "11111110101101100000110001011101",
			774 => "0000000001000000000000111100000100",
			775 => "00000001110000000000110001011101",
			776 => "00000000000000000000110001011101",
			777 => "11111110100010010000110001011101",
			778 => "0000000111000000001110111100010000",
			779 => "0000000010000000000010000000001100",
			780 => "0000000110000000000111101000000100",
			781 => "00000000000000000000110001011101",
			782 => "0000001000000000001011000100000100",
			783 => "11111110110101100000110001011101",
			784 => "00000000000000000000110001011101",
			785 => "00000001000010100000110001011101",
			786 => "0000001000000000000101000100000100",
			787 => "00000000000000000000110001011101",
			788 => "0000001100000000000000111000000100",
			789 => "00000000000000000000110001011101",
			790 => "11111110011011010000110001011101",
			791 => "0000000110000000000111101000011100",
			792 => "0000001001000000001001111000011000",
			793 => "0000000000000000001001101000001000",
			794 => "0000001101000000001100110000000100",
			795 => "00000011010100000000110011011001",
			796 => "00000100111101000000110011011001",
			797 => "0000000010000000000001001000000100",
			798 => "11111110001110100000110011011001",
			799 => "0000001100000000000111111000001000",
			800 => "0000000011000000000001110100000100",
			801 => "11111111001101100000110011011001",
			802 => "00000010011111000000110011011001",
			803 => "11111111100101010000110011011001",
			804 => "11111110011001100000110011011001",
			805 => "0000001100000000000000110000001000",
			806 => "0000000010000000001100010100000100",
			807 => "11111110011001100000110011011001",
			808 => "00000010011101110000110011011001",
			809 => "0000000100000000000101110000000100",
			810 => "00000011000101010000110011011001",
			811 => "0000000111000000000000110000001000",
			812 => "0000001100000000001010000000000100",
			813 => "11111110100101010000110011011001",
			814 => "00000011101000110000110011011001",
			815 => "0000000100000000001000110100001100",
			816 => "0000001101000000001101000100001000",
			817 => "0000001101000000000101100100000100",
			818 => "11111110011000100000110011011001",
			819 => "00000000111100100000110011011001",
			820 => "11111110011000010000110011011001",
			821 => "11111110011000010000110011011001",
			822 => "0000000001000000000000011000010000",
			823 => "0000001111000000001110110000000100",
			824 => "00000000000000000000110101011101",
			825 => "0000000111000000001100001000001000",
			826 => "0000001101000000000100000000000100",
			827 => "00000000000000000000110101011101",
			828 => "00000001000000000000110101011101",
			829 => "00000000000000000000110101011101",
			830 => "0000000000000000001000110000101000",
			831 => "0000000100000000000110111000011100",
			832 => "0000000100000000001010000100010000",
			833 => "0000001111000000001011000000000100",
			834 => "00000000000000000000110101011101",
			835 => "0000000111000000000110000100001000",
			836 => "0000001000000000000000001000000100",
			837 => "00000000000000000000110101011101",
			838 => "00000000110001010000110101011101",
			839 => "00000000000000000000110101011101",
			840 => "0000001011000000001001110100001000",
			841 => "0000000001000000001110100000000100",
			842 => "00000000000000000000110101011101",
			843 => "11111110111100000000110101011101",
			844 => "00000000000000000000110101011101",
			845 => "0000001100000000001110001100001000",
			846 => "0000000000000000001000101100000100",
			847 => "00000000110100110000110101011101",
			848 => "00000000000000000000110101011101",
			849 => "00000000000000000000110101011101",
			850 => "0000001010000000001000100100000100",
			851 => "00000000000000000000110101011101",
			852 => "0000001100000000000000111000000100",
			853 => "00000000000000000000110101011101",
			854 => "11111110110000000000110101011101",
			855 => "0000000110000000000111101000101100",
			856 => "0000000001000000000110000000011100",
			857 => "0000000110000000001110010100001100",
			858 => "0000000100000000001111011000001000",
			859 => "0000001111000000001110110000000100",
			860 => "00000000101110110000111000010001",
			861 => "00000001101010100000111000010001",
			862 => "00000000001001110000111000010001",
			863 => "0000000111000000001110111100001000",
			864 => "0000000010000000001110010000000100",
			865 => "00000000000000000000111000010001",
			866 => "00000001101011010000111000010001",
			867 => "0000000011000000000000111000000100",
			868 => "00000000010101110000111000010001",
			869 => "11111110101100100000111000010001",
			870 => "0000001111000000000100010000001000",
			871 => "0000001111000000001011011100000100",
			872 => "11111110011011010000111000010001",
			873 => "00000000000000000000111000010001",
			874 => "0000000001000000001100110100000100",
			875 => "00000001111011100000111000010001",
			876 => "11111111110011000000111000010001",
			877 => "0000001100000000001010000000010000",
			878 => "0000001010000000000111000100001100",
			879 => "0000000010000000000011001000000100",
			880 => "11111110011110110000111000010001",
			881 => "0000000001000000000000011000000100",
			882 => "00000001100100100000111000010001",
			883 => "11111110110000100000111000010001",
			884 => "00001000001111000000111000010001",
			885 => "0000000100000000000110101100010000",
			886 => "0000001000000000000110011000000100",
			887 => "11111110011110010000111000010001",
			888 => "0000001110000000001110101000000100",
			889 => "11111111001100100000111000010001",
			890 => "0000000001000000001011111100000100",
			891 => "00000010110101100000111000010001",
			892 => "11111111101000110000111000010001",
			893 => "0000000000000000000111000000001100",
			894 => "0000001001000000000100111100001000",
			895 => "0000001111000000001010000100000100",
			896 => "11111110101101000000111000010001",
			897 => "00000010010110000000111000010001",
			898 => "11111110011101010000111000010001",
			899 => "11111110011001110000111000010001",
			900 => "0000000110000000001110010100010000",
			901 => "0000001111000000000111001000001000",
			902 => "0000001011000000001110111100000100",
			903 => "00000000000000000000111010011101",
			904 => "11111110111101110000111010011101",
			905 => "0000001001000000000110101000000100",
			906 => "00000001100110000000111010011101",
			907 => "11111111001101100000111010011101",
			908 => "0000000000000000000111000000011000",
			909 => "0000001100000000000000001100010100",
			910 => "0000001100000000001000111000000100",
			911 => "11111110110111000000111010011101",
			912 => "0000000111000000001110001100000100",
			913 => "00000010101010110000111010011101",
			914 => "0000000111000000000111001000000100",
			915 => "11111110101000000000111010011101",
			916 => "0000000001000000000000111100000100",
			917 => "00000001111111000000111010011101",
			918 => "00000000000000000000111010011101",
			919 => "11111110100000000000111010011101",
			920 => "0000000111000000001110111100010000",
			921 => "0000000011000000000001110100000100",
			922 => "11111111000100010000111010011101",
			923 => "0000000100000000000001100100001000",
			924 => "0000001000000000001011010100000100",
			925 => "00000000000000000000111010011101",
			926 => "11111111000000110000111010011101",
			927 => "00000001010011000000111010011101",
			928 => "0000001100000000000000111000000100",
			929 => "00000000000000000000111010011101",
			930 => "0000001000000000000101000100000100",
			931 => "00000000000000000000111010011101",
			932 => "0000001011000000000000110000000100",
			933 => "00000000000000000000111010011101",
			934 => "11111110011010100000111010011101",
			935 => "0000000110000000000111101000100100",
			936 => "0000000001000000001110100000011000",
			937 => "0000001111000000001101010100001000",
			938 => "0000000010000000001110101100000100",
			939 => "11111110010110010000111100111001",
			940 => "00000000101101000000111100111001",
			941 => "0000001000000000001000010100000100",
			942 => "00000101010001100000111100111001",
			943 => "0000000010000000000001001000000100",
			944 => "00000000101101000000111100111001",
			945 => "0000000010000000000010110100000100",
			946 => "00000010101000010000111100111001",
			947 => "00000011101111110000111100111001",
			948 => "0000000001000000001110100000001000",
			949 => "0000001100000000000100010100000100",
			950 => "11111110011110110000111100111001",
			951 => "00000101010011010000111100111001",
			952 => "11111110011001000000111100111001",
			953 => "0000001100000000000000110000001000",
			954 => "0000000010000000001100010100000100",
			955 => "11111110010111110000111100111001",
			956 => "00000100010000010000111100111001",
			957 => "0000000111000000001110111100001100",
			958 => "0000000011000000001000101100000100",
			959 => "11111110011001000000111100111001",
			960 => "0000000100000000001101110100000100",
			961 => "11111110100000110000111100111001",
			962 => "00001011011001110000111100111001",
			963 => "0000000100000000000110111000010100",
			964 => "0000001000000000000110011000000100",
			965 => "11111110010111100000111100111001",
			966 => "0000000100000000000110101100001000",
			967 => "0000000100000000000111010100000100",
			968 => "00000001001101000000111100111001",
			969 => "11111111100111100000111100111001",
			970 => "0000000100000000000110111000000100",
			971 => "11111110011100100000111100111001",
			972 => "11111111010100100000111100111001",
			973 => "11111110010111010000111100111001",
			974 => "0000000001000000000000011000011000",
			975 => "0000001001000000001100100000001000",
			976 => "0000000100000000001111101100000100",
			977 => "00000000000000000000111111000101",
			978 => "11111111111111010000111111000101",
			979 => "0000000111000000001100001000001100",
			980 => "0000001111000000001010111100000100",
			981 => "00000000000000000000111111000101",
			982 => "0000001101000000000100000000000100",
			983 => "00000000000000000000111111000101",
			984 => "00000001100011000000111111000101",
			985 => "00000000000000000000111111000101",
			986 => "0000001000000000000001110000101000",
			987 => "0000001100000000000100001000100100",
			988 => "0000001111000000001010010100010100",
			989 => "0000000110000000000001000100001100",
			990 => "0000001111000000001001001000000100",
			991 => "11111111110100110000111111000101",
			992 => "0000000001000000001001111000000100",
			993 => "00000000101110110000111111000101",
			994 => "00000000000000000000111111000101",
			995 => "0000001010000000001010100000000100",
			996 => "00000000000000000000111111000101",
			997 => "11111111000110000000111111000101",
			998 => "0000000001000000001101011100001100",
			999 => "0000000101000000001001010100001000",
			1000 => "0000000111000000001010111100000100",
			1001 => "00000000011001010000111111000101",
			1002 => "00000001010111000000111111000101",
			1003 => "00000000000000000000111111000101",
			1004 => "00000000000000000000111111000101",
			1005 => "11111111001001000000111111000101",
			1006 => "0000000110000000001110010100000100",
			1007 => "00000000000000000000111111000101",
			1008 => "11111110100000000000111111000101",
			1009 => "0000000110000000000001111000101000",
			1010 => "0000000010000000001111010000100000",
			1011 => "0000001010000000000011101000011000",
			1012 => "0000001111000000001110110000000100",
			1013 => "11111111010001000001000001010001",
			1014 => "0000000001000000000111100100010000",
			1015 => "0000001010000000001010100100001000",
			1016 => "0000001000000000000000001000000100",
			1017 => "00000000000000000001000001010001",
			1018 => "00000001101001110001000001010001",
			1019 => "0000000111000000000100010100000100",
			1020 => "00000000101000100001000001010001",
			1021 => "11111111101001100001000001010001",
			1022 => "11111111101010010001000001010001",
			1023 => "0000000110000000001011111100000100",
			1024 => "00000000100110100001000001010001",
			1025 => "11111110100011000001000001010001",
			1026 => "0000000111000000000000101000000100",
			1027 => "00000001100100110001000001010001",
			1028 => "11111111001110010001000001010001",
			1029 => "0000000010000000001110110100000100",
			1030 => "11111110011011100001000001010001",
			1031 => "0000001100000000000100001000011000",
			1032 => "0000000000000000000111000000010000",
			1033 => "0000001011000000001001110100001000",
			1034 => "0000001111000000000010000100000100",
			1035 => "00000000100101100001000001010001",
			1036 => "11111111011000100001000001010001",
			1037 => "0000001011000000000001101000000100",
			1038 => "00000001010111110001000001010001",
			1039 => "00000000000000000001000001010001",
			1040 => "0000001011000000001011000100000100",
			1041 => "00000000100111100001000001010001",
			1042 => "11111110101010000001000001010001",
			1043 => "11111110100001100001000001010001",
			1044 => "0000000110000000000111101000011100",
			1045 => "0000001001000000000110101000011000",
			1046 => "0000000110000000001011111100001100",
			1047 => "0000001111000000000111001000000100",
			1048 => "00000000001010110001000011101101",
			1049 => "0000001000000000000111110100000100",
			1050 => "00000010101000110001000011101101",
			1051 => "00000001101110000001000011101101",
			1052 => "0000000010000000001010001000000100",
			1053 => "11111110010111100001000011101101",
			1054 => "0000000101000000001000111000000100",
			1055 => "00000001101010110001000011101101",
			1056 => "00000000011100100001000011101101",
			1057 => "11111110100001000001000011101101",
			1058 => "0000001100000000001010000000010000",
			1059 => "0000000010000000000011001000000100",
			1060 => "11111110011011100001000011101101",
			1061 => "0000000001000000000000011000001000",
			1062 => "0000001100000000000000111000000100",
			1063 => "00000001100101010001000011101101",
			1064 => "00000010111100000001000011101101",
			1065 => "11111110110010000001000011101101",
			1066 => "0000000100000000001000110100100000",
			1067 => "0000000100000000001000000100010100",
			1068 => "0000000101000000001001010100010000",
			1069 => "0000001011000000001000011000001000",
			1070 => "0000001111000000000110010000000100",
			1071 => "11111110011011100001000011101101",
			1072 => "11111111110111000001000011101101",
			1073 => "0000000010000000001010000100000100",
			1074 => "00000000000000000001000011101101",
			1075 => "00000100001100010001000011101101",
			1076 => "11111110011010110001000011101101",
			1077 => "0000001010000000001001000100000100",
			1078 => "11111110111110110001000011101101",
			1079 => "0000000001000000000111100100000100",
			1080 => "11111111111101010001000011101101",
			1081 => "00000100001101010001000011101101",
			1082 => "11111110011001010001000011101101",
			1083 => "0000000110000000000111101000100000",
			1084 => "0000000001000000001110100000011100",
			1085 => "0000000010000000000010110100001100",
			1086 => "0000000110000000001011111100001000",
			1087 => "0000001101000000000011011100000100",
			1088 => "00000000000111000001000110001001",
			1089 => "00000001101101010001000110001001",
			1090 => "11111110011101100001000110001001",
			1091 => "0000000110000000001110010100001000",
			1092 => "0000000100000000000100100100000100",
			1093 => "00000001101011000001000110001001",
			1094 => "00000000011010110001000110001001",
			1095 => "0000000001000000000000011000000100",
			1096 => "00000001010010100001000110001001",
			1097 => "11111111000100100001000110001001",
			1098 => "11111110100111110001000110001001",
			1099 => "0000000100000000000101110000000100",
			1100 => "00000011001001000001000110001001",
			1101 => "0000000000000000000111000000010000",
			1102 => "0000000111000000001110110000001100",
			1103 => "0000001111000000000011001000000100",
			1104 => "11111110101101100001000110001001",
			1105 => "0000000001000000001001011000000100",
			1106 => "00000010100010110001000110001001",
			1107 => "11111110111101110001000110001001",
			1108 => "11111110011011100001000110001001",
			1109 => "0000000111000000001110111100001100",
			1110 => "0000000010000000000011001000000100",
			1111 => "11111110100011100001000110001001",
			1112 => "0000000110000000000001111000000100",
			1113 => "00000001100000100001000110001001",
			1114 => "00000000011011010001000110001001",
			1115 => "0000001100000000000000110000001100",
			1116 => "0000001110000000000001110100001000",
			1117 => "0000000101000000000100000000000100",
			1118 => "11111111100100010001000110001001",
			1119 => "00000000100011100001000110001001",
			1120 => "11111111000001000001000110001001",
			1121 => "11111110011001110001000110001001",
			1122 => "0000001001000000001100110100010000",
			1123 => "0000001111000000001010111100000100",
			1124 => "11111111110000100001001000001101",
			1125 => "0000000101000000001100101000001000",
			1126 => "0000001001000000001100110100000100",
			1127 => "00000001011001110001001000001101",
			1128 => "00000000000000000001001000001101",
			1129 => "00000000000000000001001000001101",
			1130 => "0000001000000000000001110000101100",
			1131 => "0000001100000000000100001000101000",
			1132 => "0000001111000000001010010100010100",
			1133 => "0000000110000000000001000100001100",
			1134 => "0000001111000000001001001000000100",
			1135 => "00000000000000000001001000001101",
			1136 => "0000000010000000000001101000000100",
			1137 => "00000000000000000001001000001101",
			1138 => "00000000001111100001001000001101",
			1139 => "0000001010000000001010100000000100",
			1140 => "00000000000000000001001000001101",
			1141 => "11111111001000110001001000001101",
			1142 => "0000001001000000000100111100010000",
			1143 => "0000000111000000000111001000001000",
			1144 => "0000000111000000000110000100000100",
			1145 => "00000000111011010001001000001101",
			1146 => "11111111001111000001001000001101",
			1147 => "0000000101000000000000110100000100",
			1148 => "00000001010011110001001000001101",
			1149 => "00000000000000000001001000001101",
			1150 => "00000000000000000001001000001101",
			1151 => "11111111001100100001001000001101",
			1152 => "0000000110000000001110010100000100",
			1153 => "00000000000000000001001000001101",
			1154 => "11111110100000110001001000001101",
			1155 => "0000000110000000001110010100010000",
			1156 => "0000000101000000001101010100001100",
			1157 => "0000000010000000001101000100001000",
			1158 => "0000000110000000000001000100000100",
			1159 => "00000001011011100001001010100011",
			1160 => "11111110100110100001001010100011",
			1161 => "00000001101000010001001010100011",
			1162 => "11111110110000110001001010100011",
			1163 => "0000000100000000000101110000000100",
			1164 => "00000001100111010001001010100011",
			1165 => "0000001001000000001110100000011100",
			1166 => "0000001111000000000100000100010000",
			1167 => "0000000110000000000111101000001000",
			1168 => "0000000010000000001110010000000100",
			1169 => "00000000000000000001001010100011",
			1170 => "00000000110110000001001010100011",
			1171 => "0000001111000000001111011100000100",
			1172 => "11111110100110010001001010100011",
			1173 => "00000000000000000001001010100011",
			1174 => "0000000110000000001010011000001000",
			1175 => "0000000101000000001010111000000100",
			1176 => "00000001001000110001001010100011",
			1177 => "00000000000000000001001010100011",
			1178 => "00000100010111000001001010100011",
			1179 => "0000000100000000000001011100010000",
			1180 => "0000000000000000001011010100000100",
			1181 => "11111110011101110001001010100011",
			1182 => "0000001110000000001110101000000100",
			1183 => "11111110111001010001001010100011",
			1184 => "0000000011000000000010000000000100",
			1185 => "00000010000000000001001010100011",
			1186 => "11111110111101010001001010100011",
			1187 => "0000000110000000000111101000001000",
			1188 => "0000001000000000000001010100000100",
			1189 => "00000000000011000001001010100011",
			1190 => "11111111000101000001001010100011",
			1191 => "11111110011100110001001010100011",
			1192 => "00000000000000000001001010100101",
			1193 => "00000000000000000001001010101001",
			1194 => "00000000000000000001001010101101",
			1195 => "00000000000000000001001010110001",
			1196 => "00000000000000000001001010110101",
			1197 => "00000000000000000001001010111001",
			1198 => "00000000000000000001001010111101",
			1199 => "00000000000000000001001011000001",
			1200 => "00000000000000000001001011000101",
			1201 => "00000000000000000001001011001001",
			1202 => "00000000000000000001001011001101",
			1203 => "00000000000000000001001011010001",
			1204 => "00000000000000000001001011010101",
			1205 => "00000000000000000001001011011001",
			1206 => "00000000000000000001001011011101",
			1207 => "00000000000000000001001011100001",
			1208 => "00000000000000000001001011100101",
			1209 => "00000000000000000001001011101001",
			1210 => "00000000000000000001001011101101",
			1211 => "0000000111000000001110001100000100",
			1212 => "00000000000101000001001011111001",
			1213 => "00000000000000000001001011111001",
			1214 => "0000000111000000000100010100000100",
			1215 => "00000000000000000001001100000101",
			1216 => "11111111111011110001001100000101",
			1217 => "0000000001000000000110000000001000",
			1218 => "0000000001000000001110011100000100",
			1219 => "00000000000000000001001100011001",
			1220 => "00000000000011010001001100011001",
			1221 => "00000000000000000001001100011001",
			1222 => "0000000110000000000001111000001000",
			1223 => "0000000110000000001101011100000100",
			1224 => "00000000000000000001001100101101",
			1225 => "00000000000000010001001100101101",
			1226 => "11111111111000110001001100101101",
			1227 => "0000000001000000000110000000001000",
			1228 => "0000000001000000001110011100000100",
			1229 => "00000000000000000001001101000001",
			1230 => "00000000000011100001001101000001",
			1231 => "00000000000000000001001101000001",
			1232 => "0000000111000000000111111000000100",
			1233 => "00000000000000000001001101010101",
			1234 => "0000000111000000000111001000000100",
			1235 => "11111111111110000001001101010101",
			1236 => "00000000000000000001001101010101",
			1237 => "0000000111000000001110001100001000",
			1238 => "0000001001000000001100100000000100",
			1239 => "00000000000000000001001101101001",
			1240 => "00000000000110010001001101101001",
			1241 => "00000000000000000001001101101001",
			1242 => "0000000110000000001110010100000100",
			1243 => "00000000000000000001001101111101",
			1244 => "0000000110000000001111000000000100",
			1245 => "11111111111011110001001101111101",
			1246 => "00000000000000000001001101111101",
			1247 => "0000000001000000001110100000001100",
			1248 => "0000000001000000001110011100000100",
			1249 => "00000000000000000001001110011001",
			1250 => "0000000001000000000110000000000100",
			1251 => "00000000000011100001001110011001",
			1252 => "00000000000000000001001110011001",
			1253 => "11111111111111110001001110011001",
			1254 => "0000001111000000001001001000000100",
			1255 => "00000000000000000001001110110101",
			1256 => "0000001011000000001010111000001000",
			1257 => "0000001100000000001100110000000100",
			1258 => "00000000010000000001001110110101",
			1259 => "00000000000000000001001110110101",
			1260 => "00000000000000000001001110110101",
			1261 => "0000001011000000001010111000001100",
			1262 => "0000001111000000001110110000000100",
			1263 => "00000000000000000001001111010001",
			1264 => "0000000111000000001110001100000100",
			1265 => "00000000001110000001001111010001",
			1266 => "00000000000000000001001111010001",
			1267 => "00000000000000000001001111010001",
			1268 => "0000000110000000000001111000001100",
			1269 => "0000000110000000001101011100000100",
			1270 => "00000000000000000001001111101101",
			1271 => "0000000110000000001011111100000100",
			1272 => "00000000001000000001001111101101",
			1273 => "00000000000000000001001111101101",
			1274 => "11111111110111010001001111101101",
			1275 => "0000000110000000001110010100000100",
			1276 => "00000000000000000001010000001001",
			1277 => "0000000110000000001010011000001000",
			1278 => "0000000110000000001110010100000100",
			1279 => "00000000000000000001010000001001",
			1280 => "11111111110010110001010000001001",
			1281 => "00000000000000000001010000001001",
			1282 => "0000000110000000001101111100001100",
			1283 => "0000001010000000001001100100000100",
			1284 => "00000000000000000001010000101101",
			1285 => "0000001010000000001111001000000100",
			1286 => "00000000001100110001010000101101",
			1287 => "00000000000000000001010000101101",
			1288 => "0000000110000000001001100100000100",
			1289 => "11111111100111110001010000101101",
			1290 => "00000000000000000001010000101101",
			1291 => "0000000110000000001011111100001000",
			1292 => "0000000110000000001101011100000100",
			1293 => "00000000000000000001010001010001",
			1294 => "00000000000000110001010001010001",
			1295 => "0000001100000000000000110000000100",
			1296 => "00000000000000000001010001010001",
			1297 => "0000001011000000000000110000000100",
			1298 => "00000000000000000001010001010001",
			1299 => "11111111101101100001010001010001",
			1300 => "0000000110000000001101111100001100",
			1301 => "0000001000000000000000001000000100",
			1302 => "00000000000000000001010001111101",
			1303 => "0000001010000000000011101000000100",
			1304 => "00000000010011110001010001111101",
			1305 => "00000000000000000001010001111101",
			1306 => "0000000110000000001001100100001000",
			1307 => "0000000100000000000110101100000100",
			1308 => "00000000000000000001010001111101",
			1309 => "11111111011011000001010001111101",
			1310 => "00000000000000000001010001111101",
			1311 => "0000000111000000000111001000010000",
			1312 => "0000001111000000000101100100000100",
			1313 => "00000000000000000001010010100001",
			1314 => "0000001000000000000011101000000100",
			1315 => "00000000000000000001010010100001",
			1316 => "0000000001000000001101011100000100",
			1317 => "00000000010010100001010010100001",
			1318 => "00000000000000000001010010100001",
			1319 => "00000000000000000001010010100001",
			1320 => "0000000111000000000110000100010000",
			1321 => "0000001101000000000100000000000100",
			1322 => "00000000000000000001010011000101",
			1323 => "0000000110000000001101111100001000",
			1324 => "0000000110000000001001011000000100",
			1325 => "00000000000000000001010011000101",
			1326 => "00000000000100000001010011000101",
			1327 => "00000000000000000001010011000101",
			1328 => "11111111101000010001010011000101",
			1329 => "0000000111000000001110001100010000",
			1330 => "0000001111000000000100011000000100",
			1331 => "00000000000000000001010011101001",
			1332 => "0000000001000000001011101000001000",
			1333 => "0000001100000000001100110000000100",
			1334 => "00000000010011010001010011101001",
			1335 => "00000000000000000001010011101001",
			1336 => "00000000000000000001010011101001",
			1337 => "00000000000000000001010011101001",
			1338 => "0000000111000000001110001100010000",
			1339 => "0000001111000000001010111100000100",
			1340 => "00000000000000000001010100001101",
			1341 => "0000001100000000001100110000001000",
			1342 => "0000001011000000000000111000000100",
			1343 => "00000000000000000001010100001101",
			1344 => "00000000001101000001010100001101",
			1345 => "00000000000000000001010100001101",
			1346 => "00000000000000000001010100001101",
			1347 => "0000000001000000000110000000010000",
			1348 => "0000001111000000001110110000000100",
			1349 => "00000000000000000001010100111001",
			1350 => "0000000101000000001100101000001000",
			1351 => "0000001100000000000100010100000100",
			1352 => "00000000011001010001010100111001",
			1353 => "00000000000000000001010100111001",
			1354 => "00000000000000000001010100111001",
			1355 => "0000000000000000001001101000000100",
			1356 => "00000000000000000001010100111001",
			1357 => "11111111001101000001010100111001",
			1358 => "0000000111000000001110001100010100",
			1359 => "0000001011000000000100001000001100",
			1360 => "0000000110000000001110010100001000",
			1361 => "0000000110000000001101011100000100",
			1362 => "00000000000000000001010101100101",
			1363 => "00000000000111110001010101100101",
			1364 => "11111111110001110001010101100101",
			1365 => "0000000110000000000111101000000100",
			1366 => "00000000000000000001010101100101",
			1367 => "00000000011101110001010101100101",
			1368 => "11111111100101000001010101100101",
			1369 => "0000000110000000001101111100010000",
			1370 => "0000001111000000001001001000000100",
			1371 => "00000000000000000001010110011001",
			1372 => "0000000111000000000110000100001000",
			1373 => "0000001010000000000111110100000100",
			1374 => "00000000010010110001010110011001",
			1375 => "00000000000000000001010110011001",
			1376 => "00000000000000000001010110011001",
			1377 => "0000000100000000000110111100000100",
			1378 => "00000000000000000001010110011001",
			1379 => "0000000110000000001001100100000100",
			1380 => "11111111010111000001010110011001",
			1381 => "00000000000000000001010110011001",
			1382 => "0000000001000000001110100000010000",
			1383 => "0000000101000000001010111000001100",
			1384 => "0000001101000000000011011100000100",
			1385 => "00000000000000000001010111010101",
			1386 => "0000000101000000001000111000000100",
			1387 => "00000000000000000001010111010101",
			1388 => "00000000011011000001010111010101",
			1389 => "00000000000000000001010111010101",
			1390 => "0000001101000000000010001000001000",
			1391 => "0000000110000000001001011000000100",
			1392 => "00000000000000000001010111010101",
			1393 => "11111111100111110001010111010101",
			1394 => "0000001001000000001011001100000100",
			1395 => "00000000000001110001010111010101",
			1396 => "00000000000000000001010111010101",
			1397 => "0000001100000000001010000000010000",
			1398 => "0000001011000000001011000100001100",
			1399 => "0000001001000000001100100000000100",
			1400 => "00000000000000000001011000010001",
			1401 => "0000000001000000001110100000000100",
			1402 => "00000000001101110001011000010001",
			1403 => "00000000000000000001011000010001",
			1404 => "00000000000000000001011000010001",
			1405 => "0000000110000000001010011000001100",
			1406 => "0000000110000000001011111100000100",
			1407 => "00000000000000000001011000010001",
			1408 => "0000000111000000001010000000000100",
			1409 => "00000000000000000001011000010001",
			1410 => "11111111100000100001011000010001",
			1411 => "00000000000000000001011000010001",
			1412 => "0000000111000000001110110000010100",
			1413 => "0000001111000000001110110000000100",
			1414 => "00000000000000000001011000111101",
			1415 => "0000000001000000001110011100000100",
			1416 => "00000000000000000001011000111101",
			1417 => "0000000001000000001101011100001000",
			1418 => "0000000101000000001001010100000100",
			1419 => "00000000001001010001011000111101",
			1420 => "00000000000000000001011000111101",
			1421 => "00000000000000000001011000111101",
			1422 => "00000000000000000001011000111101",
			1423 => "0000000010000000001100010100011000",
			1424 => "0000000110000000001011111100001100",
			1425 => "0000001001000000000110101000001000",
			1426 => "0000000110000000001001011000000100",
			1427 => "00000000000000000001011010000001",
			1428 => "00000000000101100001011010000001",
			1429 => "00000000000000000001011010000001",
			1430 => "0000001010000000000111101100000100",
			1431 => "00000000000000000001011010000001",
			1432 => "0000001001000000000000011000000100",
			1433 => "00000000000000000001011010000001",
			1434 => "11111111010111100001011010000001",
			1435 => "0000000111000000001110001100001000",
			1436 => "0000000001000000001011101000000100",
			1437 => "00000000100111010001011010000001",
			1438 => "00000000000000000001011010000001",
			1439 => "00000000000000000001011010000001",
			1440 => "0000000010000000001100010100001100",
			1441 => "0000000110000000000001000100000100",
			1442 => "00000000000000000001011010111101",
			1443 => "0000001010000000000111101100000100",
			1444 => "00000000000000000001011010111101",
			1445 => "11111111100010000001011010111101",
			1446 => "0000000111000000001110110000010000",
			1447 => "0000000001000000001101011100001100",
			1448 => "0000000100000000001101001100001000",
			1449 => "0000000010000000000011000000000100",
			1450 => "00000000100110100001011010111101",
			1451 => "00000000000000000001011010111101",
			1452 => "00000000000000000001011010111101",
			1453 => "00000000000000000001011010111101",
			1454 => "00000000000000000001011010111101",
			1455 => "0000001100000000001010000000010100",
			1456 => "0000000010000000001010010100000100",
			1457 => "00000000000000000001011100000001",
			1458 => "0000000001000000001110100000001100",
			1459 => "0000000001000000001110011100000100",
			1460 => "00000000000000000001011100000001",
			1461 => "0000000111000000000100010100000100",
			1462 => "00000000010110110001011100000001",
			1463 => "00000000000000000001011100000001",
			1464 => "00000000000000000001011100000001",
			1465 => "0000000010000000000111010100001100",
			1466 => "0000001011000000001001110100001000",
			1467 => "0000000111000000001010000000000100",
			1468 => "00000000000000000001011100000001",
			1469 => "11111111110011110001011100000001",
			1470 => "00000000000000000001011100000001",
			1471 => "00000000000000000001011100000001",
			1472 => "0000000001000000001110100000010000",
			1473 => "0000001111000000001011000000000100",
			1474 => "00000000000000000001011101001101",
			1475 => "0000001100000000000100010100001000",
			1476 => "0000000110000000001110010100000100",
			1477 => "00000000111001010001011101001101",
			1478 => "00000000000000000001011101001101",
			1479 => "00000000000000000001011101001101",
			1480 => "0000001111000000001100010000001000",
			1481 => "0000001010000000000100101100000100",
			1482 => "00000000000000000001011101001101",
			1483 => "11111111000100000001011101001101",
			1484 => "0000001001000000001111000000001100",
			1485 => "0000001011000000000001101000001000",
			1486 => "0000001001000000001100011000000100",
			1487 => "00000000000000000001011101001101",
			1488 => "00000000001100000001011101001101",
			1489 => "00000000000000000001011101001101",
			1490 => "00000000000000000001011101001101",
			1491 => "0000001001000000000010001100001100",
			1492 => "0000000011000000001010101100000100",
			1493 => "00000000000000000001011110011001",
			1494 => "0000000111000000001100001000000100",
			1495 => "00000000100000100001011110011001",
			1496 => "00000000000000000001011110011001",
			1497 => "0000000110000000001101011000010000",
			1498 => "0000000000000000001001101000000100",
			1499 => "00000000000000000001011110011001",
			1500 => "0000000110000000001011111100000100",
			1501 => "00000000000000000001011110011001",
			1502 => "0000001100000000000000111000000100",
			1503 => "00000000000000000001011110011001",
			1504 => "11111111000011110001011110011001",
			1505 => "0000000001000000001101011100001000",
			1506 => "0000000001000000001101011100000100",
			1507 => "00000000000000000001011110011001",
			1508 => "00000000010101110001011110011001",
			1509 => "00000000000000000001011110011001",
			1510 => "0000000110000000001101111100011100",
			1511 => "0000001111000000000010001000010100",
			1512 => "0000000110000000000001000100001100",
			1513 => "0000000001000000000110000000001000",
			1514 => "0000000001000000001110011100000100",
			1515 => "00000000000000000001011111101101",
			1516 => "00000000001110110001011111101101",
			1517 => "00000000000000000001011111101101",
			1518 => "0000000001000000001100100000000100",
			1519 => "00000000000000000001011111101101",
			1520 => "11111111100010000001011111101101",
			1521 => "0000001011000000001101010100000100",
			1522 => "00000000101010000001011111101101",
			1523 => "00000000000000000001011111101101",
			1524 => "0000000010000000001011111000001000",
			1525 => "0000001011000000001001110100000100",
			1526 => "11111111000100010001011111101101",
			1527 => "00000000000000000001011111101101",
			1528 => "0000001100000000000011011100000100",
			1529 => "00000000011100010001011111101101",
			1530 => "00000000000000000001011111101101",
			1531 => "0000000111000000001110001100100000",
			1532 => "0000000010000000001110010000010100",
			1533 => "0000001010000000001010100000001100",
			1534 => "0000001110000000000100000000000100",
			1535 => "00000000000000000001100000111001",
			1536 => "0000000110000000001001011000000100",
			1537 => "00000000000000000001100000111001",
			1538 => "00000000000110110001100000111001",
			1539 => "0000000110000000000001000100000100",
			1540 => "00000000000000000001100000111001",
			1541 => "11111111011100010001100000111001",
			1542 => "0000000001000000001011101000001000",
			1543 => "0000001100000000000011011100000100",
			1544 => "00000000100100010001100000111001",
			1545 => "00000000000000000001100000111001",
			1546 => "00000000000000000001100000111001",
			1547 => "0000000110000000001001100100000100",
			1548 => "11111111110111000001100000111001",
			1549 => "00000000000000000001100000111001",
			1550 => "0000001000000000000001110000011000",
			1551 => "0000000111000000001110110000010100",
			1552 => "0000001111000000001110110000000100",
			1553 => "00000000000000000001100001111101",
			1554 => "0000000001000000001001011000001100",
			1555 => "0000001000000000000000001000000100",
			1556 => "00000000000000000001100001111101",
			1557 => "0000000101000000001001010100000100",
			1558 => "00000000100011010001100001111101",
			1559 => "00000000000000000001100001111101",
			1560 => "00000000000000000001100001111101",
			1561 => "00000000000000000001100001111101",
			1562 => "0000000110000000001110010100000100",
			1563 => "00000000000000000001100001111101",
			1564 => "0000001001000000000110000000000100",
			1565 => "00000000000000000001100001111101",
			1566 => "11111111000110110001100001111101",
			1567 => "0000001011000000001011000100011000",
			1568 => "0000001101000000000000101000000100",
			1569 => "00000000000000000001100011001001",
			1570 => "0000001100000000001010000000010000",
			1571 => "0000001001000000001001111000001100",
			1572 => "0000000111000000000100010100001000",
			1573 => "0000001001000000001100100000000100",
			1574 => "00000000000000000001100011001001",
			1575 => "00000000010001010001100011001001",
			1576 => "00000000000000000001100011001001",
			1577 => "00000000000000000001100011001001",
			1578 => "00000000000000000001100011001001",
			1579 => "0000001101000000000010001000001000",
			1580 => "0000001001000000000010001100000100",
			1581 => "00000000000000000001100011001001",
			1582 => "11111111101000110001100011001001",
			1583 => "0000001001000000001011001100000100",
			1584 => "00000000000010100001100011001001",
			1585 => "00000000000000000001100011001001",
			1586 => "0000000110000000001101111100100000",
			1587 => "0000001111000000001010010100010100",
			1588 => "0000000110000000001011111100001100",
			1589 => "0000001111000000000111001000000100",
			1590 => "00000000000000000001100100101101",
			1591 => "0000000101000000000100011000000100",
			1592 => "00000000110111000001100100101101",
			1593 => "00000000000000000001100100101101",
			1594 => "0000001001000000000110000000000100",
			1595 => "00000000000000000001100100101101",
			1596 => "11111111000100000001100100101101",
			1597 => "0000000111000000000110000100001000",
			1598 => "0000001010000000000001010000000100",
			1599 => "00000000111101010001100100101101",
			1600 => "00000000000000000001100100101101",
			1601 => "00000000000000000001100100101101",
			1602 => "0000000010000000001100111000001000",
			1603 => "0000000111000000000111001000000100",
			1604 => "11111110101101000001100100101101",
			1605 => "00000000000000000001100100101101",
			1606 => "0000000111000000000111001000001000",
			1607 => "0000000010000000000011000000000100",
			1608 => "00000000101110000001100100101101",
			1609 => "00000000000000000001100100101101",
			1610 => "00000000000000000001100100101101",
			1611 => "0000001000000000000101000100011000",
			1612 => "0000001100000000000100001000010100",
			1613 => "0000001110000000000010111100000100",
			1614 => "00000000000000000001100101111001",
			1615 => "0000001110000000000011001000001100",
			1616 => "0000001010000000000011101000001000",
			1617 => "0000001000000000000000001000000100",
			1618 => "00000000000000000001100101111001",
			1619 => "00000000011111000001100101111001",
			1620 => "00000000000000000001100101111001",
			1621 => "00000000000000000001100101111001",
			1622 => "00000000000000000001100101111001",
			1623 => "0000001100000000000000110000000100",
			1624 => "00000000000000000001100101111001",
			1625 => "0000001110000000000111010100001000",
			1626 => "0000001110000000000001010100000100",
			1627 => "00000000000000000001100101111001",
			1628 => "11111111011111110001100101111001",
			1629 => "00000000000000000001100101111001",
			1630 => "0000000110000000001101111100100100",
			1631 => "0000001111000000001010010100011000",
			1632 => "0000000110000000000001000100001100",
			1633 => "0000001111000000001010111100000100",
			1634 => "00000000000000000001100111101101",
			1635 => "0000000101000000000100011000000100",
			1636 => "00000000110011010001100111101101",
			1637 => "00000000000000000001100111101101",
			1638 => "0000000001000000000000011000000100",
			1639 => "00000000000000000001100111101101",
			1640 => "0000001010000000001010100000000100",
			1641 => "00000000000000000001100111101101",
			1642 => "11111111000001100001100111101101",
			1643 => "0000000111000000000110000100001000",
			1644 => "0000001010000000000001010000000100",
			1645 => "00000000111010000001100111101101",
			1646 => "00000000000000000001100111101101",
			1647 => "00000000000000000001100111101101",
			1648 => "0000000010000000001100111000001100",
			1649 => "0000000111000000000111001000001000",
			1650 => "0000000001000000001100100000000100",
			1651 => "00000000000000000001100111101101",
			1652 => "11111110101110000001100111101101",
			1653 => "00000000000000000001100111101101",
			1654 => "0000000111000000000111001000001000",
			1655 => "0000000010000000000011000000000100",
			1656 => "00000000101010000001100111101101",
			1657 => "00000000000000000001100111101101",
			1658 => "00000000000000000001100111101101",
			1659 => "0000000010000000001100010100010100",
			1660 => "0000000110000000000001111000010000",
			1661 => "0000000010000000000001101000000100",
			1662 => "00000000000000000001101001000001",
			1663 => "0000000110000000001011111100001000",
			1664 => "0000000001000000001110100000000100",
			1665 => "00000000010101100001101001000001",
			1666 => "00000000000000000001101001000001",
			1667 => "00000000000000000001101001000001",
			1668 => "11111111011011000001101001000001",
			1669 => "0000000001000000001101011100010100",
			1670 => "0000001100000000000100001000010000",
			1671 => "0000001001000000001100100000000100",
			1672 => "00000000000000000001101001000001",
			1673 => "0000000000000000000110110100001000",
			1674 => "0000000010000000000011000000000100",
			1675 => "00000000101011010001101001000001",
			1676 => "00000000000000000001101001000001",
			1677 => "00000000000000000001101001000001",
			1678 => "00000000000000000001101001000001",
			1679 => "00000000000000000001101001000001",
			1680 => "0000000001000000000110000000011000",
			1681 => "0000000010000000000100101000010000",
			1682 => "0000000110000000001011111100001000",
			1683 => "0000000011000000000000111000000100",
			1684 => "00000000000000000001101010111101",
			1685 => "00000000001000010001101010111101",
			1686 => "0000001110000000000000110000000100",
			1687 => "11111111110001100001101010111101",
			1688 => "00000000000000000001101010111101",
			1689 => "0000000111000000000000101000000100",
			1690 => "00000000110100110001101010111101",
			1691 => "00000000000000000001101010111101",
			1692 => "0000000111000000000101101100010000",
			1693 => "0000000000000000000101000100000100",
			1694 => "00000000000000000001101010111101",
			1695 => "0000000010000000001100010000001000",
			1696 => "0000001100000000000000111000000100",
			1697 => "00000000000000000001101010111101",
			1698 => "11111110111110110001101010111101",
			1699 => "00000000000000000001101010111101",
			1700 => "0000000111000000001110001100001100",
			1701 => "0000000110000000001010011000001000",
			1702 => "0000000010000000000000110100000100",
			1703 => "00000000000000000001101010111101",
			1704 => "00000000101111110001101010111101",
			1705 => "00000000000000000001101010111101",
			1706 => "0000000110000000001001100100001000",
			1707 => "0000000100000000000110111100000100",
			1708 => "00000000000000000001101010111101",
			1709 => "11111111011100000001101010111101",
			1710 => "00000000000000000001101010111101",
			1711 => "0000001010000000001001000100100100",
			1712 => "0000000111000000001110110000100000",
			1713 => "0000001110000000001110101000010100",
			1714 => "0000000001000000001110100000001100",
			1715 => "0000001101000000000100000000000100",
			1716 => "00000000000000000001101100011001",
			1717 => "0000000110000000001110010100000100",
			1718 => "00000000101110110001101100011001",
			1719 => "00000000000000000001101100011001",
			1720 => "0000000100000000001110010000000100",
			1721 => "00000000000000000001101100011001",
			1722 => "11111111011110000001101100011001",
			1723 => "0000001001000000001011001100001000",
			1724 => "0000000000000000001001101000000100",
			1725 => "00000000000000000001101100011001",
			1726 => "00000000111000110001101100011001",
			1727 => "00000000000000000001101100011001",
			1728 => "00000000000000000001101100011001",
			1729 => "0000000110000000000001111000000100",
			1730 => "00000000000000000001101100011001",
			1731 => "0000000001000000001100100000000100",
			1732 => "00000000000000000001101100011001",
			1733 => "11111111001010100001101100011001",
			1734 => "0000000001000000000110000000011000",
			1735 => "0000000010000000000100101000010000",
			1736 => "0000000110000000001011111100001000",
			1737 => "0000000011000000001000101100000100",
			1738 => "00000000000000000001101110000101",
			1739 => "00000000101100000001101110000101",
			1740 => "0000001110000000000000110000000100",
			1741 => "11111111011011100001101110000101",
			1742 => "00000000000000000001101110000101",
			1743 => "0000000111000000000000101000000100",
			1744 => "00000001001111110001101110000101",
			1745 => "00000000000000000001101110000101",
			1746 => "0000001100000000000011011100001000",
			1747 => "0000000110000000001110010100000100",
			1748 => "00000000000000000001101110000101",
			1749 => "11111110101011010001101110000101",
			1750 => "0000001100000000000000001100010100",
			1751 => "0000001110000000001011011100000100",
			1752 => "00000000000000000001101110000101",
			1753 => "0000000000000000000111000000001100",
			1754 => "0000000000000000000110011100000100",
			1755 => "00000000000000000001101110000101",
			1756 => "0000000111000000000111001000000100",
			1757 => "00000001001010010001101110000101",
			1758 => "00000000000000000001101110000101",
			1759 => "00000000000000000001101110000101",
			1760 => "11111111010100010001101110000101",
			1761 => "0000000001000000000110000000011000",
			1762 => "0000001111000000001110110000000100",
			1763 => "00000000000000000001101111110001",
			1764 => "0000001101000000000001111100010000",
			1765 => "0000001101000000000100000000000100",
			1766 => "00000000000000000001101111110001",
			1767 => "0000001100000000000100010100001000",
			1768 => "0000001100000000000011111100000100",
			1769 => "00000000000000000001101111110001",
			1770 => "00000000101010010001101111110001",
			1771 => "00000000000000000001101111110001",
			1772 => "00000000000000000001101111110001",
			1773 => "0000000001000000001101101000001100",
			1774 => "0000000111000000001110111100000100",
			1775 => "00000000000000000001101111110001",
			1776 => "0000000110000000001001011000000100",
			1777 => "00000000000000000001101111110001",
			1778 => "11111111000011010001101111110001",
			1779 => "0000000001000000001101011100010000",
			1780 => "0000001100000000000100001000001100",
			1781 => "0000001100000000001000111000000100",
			1782 => "00000000000000000001101111110001",
			1783 => "0000000111000000001110110000000100",
			1784 => "00000000001101010001101111110001",
			1785 => "00000000000000000001101111110001",
			1786 => "00000000000000000001101111110001",
			1787 => "00000000000000000001101111110001",
			1788 => "0000000001000000000110000000011000",
			1789 => "0000001111000000001011000000001100",
			1790 => "0000001100000000000000110000000100",
			1791 => "00000000000000000001110001101101",
			1792 => "0000000111000000000000110000000100",
			1793 => "00000000000000000001110001101101",
			1794 => "11111111101010100001110001101101",
			1795 => "0000001101000000000001111100001000",
			1796 => "0000000001000000000000011000000100",
			1797 => "00000001001001110001110001101101",
			1798 => "00000000000000000001110001101101",
			1799 => "00000000000000000001110001101101",
			1800 => "0000000000000000000111000000011100",
			1801 => "0000000001000000001101011100011000",
			1802 => "0000001111000000000011001000001100",
			1803 => "0000000001000000001110100000001000",
			1804 => "0000000011000000000110000100000100",
			1805 => "00000000000000000001110001101101",
			1806 => "00000000011000100001110001101101",
			1807 => "11111111001001110001110001101101",
			1808 => "0000001001000000001011001100001000",
			1809 => "0000001101000000000010110100000100",
			1810 => "00000001000001110001110001101101",
			1811 => "00000000000000000001110001101101",
			1812 => "00000000000000000001110001101101",
			1813 => "11111111010111110001110001101101",
			1814 => "0000001001000000000010001100000100",
			1815 => "00000000000000000001110001101101",
			1816 => "0000001000000000000101000100000100",
			1817 => "00000000000000000001110001101101",
			1818 => "11111110100101100001110001101101",
			1819 => "0000001000000000000101000100100100",
			1820 => "0000000011000000000010000000100000",
			1821 => "0000000010000000001100010100011000",
			1822 => "0000001010000000001010100000001100",
			1823 => "0000001101000000001010011100001000",
			1824 => "0000000010000000000001101000000100",
			1825 => "00000000000000000001110011100001",
			1826 => "00000000101100000001110011100001",
			1827 => "00000000000000000001110011100001",
			1828 => "0000000001000000000110000000000100",
			1829 => "00000000000000000001110011100001",
			1830 => "0000001011000000001011000100000100",
			1831 => "00000000000000000001110011100001",
			1832 => "11111111011101110001110011100001",
			1833 => "0000000001000000001011111100000100",
			1834 => "00000001000001000001110011100001",
			1835 => "00000000000000000001110011100001",
			1836 => "11111111110011100001110011100001",
			1837 => "0000000110000000001110010100001000",
			1838 => "0000001101000000001100110000000100",
			1839 => "00000000011000010001110011100001",
			1840 => "00000000000000000001110011100001",
			1841 => "0000001001000000000110000000000100",
			1842 => "00000000000000000001110011100001",
			1843 => "0000000000000000000111000000000100",
			1844 => "00000000000000000001110011100001",
			1845 => "0000001100000000000000111000000100",
			1846 => "00000000000000000001110011100001",
			1847 => "11111110110000100001110011100001",
			1848 => "0000001100000000001010000000011000",
			1849 => "0000000001000000000000011000001000",
			1850 => "0000001111000000001010111100000100",
			1851 => "00000000000000000001110101100101",
			1852 => "00000001010001010001110101100101",
			1853 => "0000001110000000001011000100001000",
			1854 => "0000001111000000000111110000000100",
			1855 => "11111111100101010001110101100101",
			1856 => "00000000000000000001110101100101",
			1857 => "0000001010000000001001000100000100",
			1858 => "00000000101011010001110101100101",
			1859 => "00000000000000000001110101100101",
			1860 => "0000000000000000000111000000011100",
			1861 => "0000001100000000000000001100011000",
			1862 => "0000001100000000000011011100001100",
			1863 => "0000000001000000001110100000001000",
			1864 => "0000001110000000001110111100000100",
			1865 => "00000000000000000001110101100101",
			1866 => "00000000001001100001110101100101",
			1867 => "11111111001111010001110101100101",
			1868 => "0000001000000000000111110100000100",
			1869 => "00000000000000000001110101100101",
			1870 => "0000000001000000000101011100000100",
			1871 => "00000001001100100001110101100101",
			1872 => "00000000000000000001110101100101",
			1873 => "11111111011101110001110101100101",
			1874 => "0000001000000000000101000100000100",
			1875 => "00000000000000000001110101100101",
			1876 => "0000000111000000001010000000000100",
			1877 => "00000000000000000001110101100101",
			1878 => "0000001011000000000000110000000100",
			1879 => "00000000000000000001110101100101",
			1880 => "11111110101011100001110101100101",
			1881 => "0000000110000000000001111000100100",
			1882 => "0000000010000000000101001000011100",
			1883 => "0000001010000000000011101000010100",
			1884 => "0000001111000000001110110000000100",
			1885 => "11111111100001010001110111110001",
			1886 => "0000000111000000000110000100001100",
			1887 => "0000000000000000000011101000000100",
			1888 => "00000000000000000001110111110001",
			1889 => "0000001010000000000010101100000100",
			1890 => "00000001010000100001110111110001",
			1891 => "00000000000000000001110111110001",
			1892 => "00000000000000000001110111110001",
			1893 => "0000000110000000001011111100000100",
			1894 => "00000000000000000001110111110001",
			1895 => "11111110101111100001110111110001",
			1896 => "0000000111000000000000101000000100",
			1897 => "00000001010111110001110111110001",
			1898 => "00000000000000000001110111110001",
			1899 => "0000000000000000000111000000011000",
			1900 => "0000000000000000000010101000001100",
			1901 => "0000001110000000001001010000001000",
			1902 => "0000001111000000001100010100000100",
			1903 => "11111111010100110001110111110001",
			1904 => "00000000110110010001110111110001",
			1905 => "11111110101110010001110111110001",
			1906 => "0000001100000000001110001100001000",
			1907 => "0000001010000000000111110100000100",
			1908 => "00000000000000000001110111110001",
			1909 => "00000001000010010001110111110001",
			1910 => "11111111110011100001110111110001",
			1911 => "0000001100000000000000111000000100",
			1912 => "00000000000000000001110111110001",
			1913 => "0000000111000000001110111100000100",
			1914 => "00000000000000000001110111110001",
			1915 => "11111110011101110001110111110001",
			1916 => "0000001100000000001010000000011100",
			1917 => "0000001001000000001100110100001100",
			1918 => "0000001111000000001010111100000100",
			1919 => "00000000000000000001111001110101",
			1920 => "0000001101000000000100000000000100",
			1921 => "00000000000000000001111001110101",
			1922 => "00000001101010110001111001110101",
			1923 => "0000001110000000001000111100001000",
			1924 => "0000001110000000001011000100000100",
			1925 => "11111111011001000001111001110101",
			1926 => "00000000000000000001111001110101",
			1927 => "0000001010000000001001000100000100",
			1928 => "00000000111100100001111001110101",
			1929 => "00000000000000000001111001110101",
			1930 => "0000001000000000000001110000100000",
			1931 => "0000001100000000000000001100011100",
			1932 => "0000001010000000001000100100010100",
			1933 => "0000001001000000001001111000001000",
			1934 => "0000001110000000000011111100000100",
			1935 => "00000000000000000001111001110101",
			1936 => "00000000111000110001111001110101",
			1937 => "0000000000000000001001101000001000",
			1938 => "0000001111000000001001011100000100",
			1939 => "00000000000000000001111001110101",
			1940 => "00000000101111010001111001110101",
			1941 => "11111110101111000001111001110101",
			1942 => "0000001110000000000100101000000100",
			1943 => "00000000000000000001111001110101",
			1944 => "00000001010101100001111001110101",
			1945 => "11111110111100000001111001110101",
			1946 => "0000000111000000001010000000000100",
			1947 => "00000000000000000001111001110101",
			1948 => "11111110100001110001111001110101",
			1949 => "0000000110000000000111101000100000",
			1950 => "0000000001000000001110100000010100",
			1951 => "0000001111000000001010111100000100",
			1952 => "11111110110000100001111100000001",
			1953 => "0000001000000000001000010100000100",
			1954 => "00000011101000110001111100000001",
			1955 => "0000001100000000000100010100001000",
			1956 => "0000000011000000000000001100000100",
			1957 => "00000010010000010001111100000001",
			1958 => "00000010110111010001111100000001",
			1959 => "11111111101101110001111100000001",
			1960 => "0000000001000000001110100000001000",
			1961 => "0000001101000000000110000100000100",
			1962 => "11111110101010100001111100000001",
			1963 => "00000001101010000001111100000001",
			1964 => "11111110011010110001111100000001",
			1965 => "0000001100000000000000110000001100",
			1966 => "0000001111000000001110110000000100",
			1967 => "11111110011010010001111100000001",
			1968 => "0000000001000000000000011000000100",
			1969 => "00000010011110000001111100000001",
			1970 => "11111110011000100001111100000001",
			1971 => "0000000100000000000101110000000100",
			1972 => "00000010100110000001111100000001",
			1973 => "0000000111000000000000110000001000",
			1974 => "0000001100000000001010000000000100",
			1975 => "11111110100111110001111100000001",
			1976 => "00000010110001110001111100000001",
			1977 => "0000000100000000001000110100001100",
			1978 => "0000000101000000001001010100001000",
			1979 => "0000001110000000000011001000000100",
			1980 => "11111110101110110001111100000001",
			1981 => "00000101110100000001111100000001",
			1982 => "11111110011000100001111100000001",
			1983 => "11111110011000100001111100000001",
			1984 => "0000000110000000001110010100010000",
			1985 => "0000001001000000000110101000001100",
			1986 => "0000001111000000000111001000000100",
			1987 => "00000000000000000001111110010101",
			1988 => "0000000100000000001111011000000100",
			1989 => "00000001101000010001111110010101",
			1990 => "00000000000001000001111110010101",
			1991 => "11111110111000010001111110010101",
			1992 => "0000001100000000001010000000011000",
			1993 => "0000000010000000001110010000001000",
			1994 => "0000000010000000001010001000000100",
			1995 => "11111110011110110001111110010101",
			1996 => "00000000000000000001111110010101",
			1997 => "0000000001000000000110000000001000",
			1998 => "0000000110000000001101111100000100",
			1999 => "00000001100100100001111110010101",
			2000 => "00000011111101100001111110010101",
			2001 => "0000000100000000000000010100000100",
			2002 => "00000000000000010001111110010101",
			2003 => "11111110111101110001111110010101",
			2004 => "0000000100000000000110101100010000",
			2005 => "0000001000000000000110011000000100",
			2006 => "11111110100001010001111110010101",
			2007 => "0000001111000000000011001000000100",
			2008 => "11111111001110010001111110010101",
			2009 => "0000001100000000000100001000000100",
			2010 => "00000010010111000001111110010101",
			2011 => "11111111101010110001111110010101",
			2012 => "0000000000000000000111000000001100",
			2013 => "0000000111000000000111001000001000",
			2014 => "0000000010000000001000001100000100",
			2015 => "11111110101111010001111110010101",
			2016 => "00000010011110110001111110010101",
			2017 => "11111110011110110001111110010101",
			2018 => "0000000111000000001010000000000100",
			2019 => "00000000000000000001111110010101",
			2020 => "11111110011001100001111110010101",
			2021 => "0000000110000000001110010100010100",
			2022 => "0000000001000000000110000000001000",
			2023 => "0000000010000000000001001000000100",
			2024 => "00000000010111010010000000010001",
			2025 => "00000001100101100010000000010001",
			2026 => "0000001111000000001010011100000100",
			2027 => "11111110101111110010000000010001",
			2028 => "0000001001000000000110101000000100",
			2029 => "00000000101111110010000000010001",
			2030 => "11111111001111110010000000010001",
			2031 => "0000000100000000000101110000000100",
			2032 => "00000010001011000010000000010001",
			2033 => "0000001100000000001010000000010100",
			2034 => "0000000010000000001100010100001000",
			2035 => "0000001000000000000100010100000100",
			2036 => "11111110100001110010000000010001",
			2037 => "00000000000000000010000000010001",
			2038 => "0000001011000000001011000100001000",
			2039 => "0000000000000000001010011100000100",
			2040 => "00000001010101100010000000010001",
			2041 => "00000011100101100010000000010001",
			2042 => "11111111100100110010000000010001",
			2043 => "0000000100000000000001011100010000",
			2044 => "0000000000000000001011010100000100",
			2045 => "11111110011100110010000000010001",
			2046 => "0000001100000000000011011100000100",
			2047 => "11111110110001100010000000010001",
			2048 => "0000000111000000001110110000000100",
			2049 => "00000010001110010010000000010001",
			2050 => "11111111000011110010000000010001",
			2051 => "11111110011100010010000000010001",
			2052 => "0000000110000000001110010100011100",
			2053 => "0000000010000000000010110100010100",
			2054 => "0000000001000000000110000000001000",
			2055 => "0000000101000000000011011100000100",
			2056 => "00000000000000000010000010110101",
			2057 => "00000001000001010010000010110101",
			2058 => "0000001110000000001000111000000100",
			2059 => "11111110111101010010000010110101",
			2060 => "0000001011000000000101101100000100",
			2061 => "00000000010110100010000010110101",
			2062 => "00000000000000000010000010110101",
			2063 => "0000000001000000001110100000000100",
			2064 => "00000001100000010010000010110101",
			2065 => "00000000000000000010000010110101",
			2066 => "0000000010000000000111010100100100",
			2067 => "0000001111000000000011001000010100",
			2068 => "0000000001000000000000011000001100",
			2069 => "0000000010000000001010001000000100",
			2070 => "11111111001100110010000010110101",
			2071 => "0000000101000000000100011000000100",
			2072 => "00000000111101010010000010110101",
			2073 => "00000000000000000010000010110101",
			2074 => "0000000101000000000100000000000100",
			2075 => "00000000000000000010000010110101",
			2076 => "11111110011101110010000010110101",
			2077 => "0000000111000000000110000100001000",
			2078 => "0000000000000000001000110000000100",
			2079 => "00000001011100110010000010110101",
			2080 => "00000000000000000010000010110101",
			2081 => "0000001000000000001010110000000100",
			2082 => "11111110110010100010000010110101",
			2083 => "00000000000000000010000010110101",
			2084 => "0000001100000000000000001100010000",
			2085 => "0000000110000000001000010000001100",
			2086 => "0000000001000000001101011100001000",
			2087 => "0000000010000000000011000000000100",
			2088 => "00000010000011010010000010110101",
			2089 => "00000000000000000010000010110101",
			2090 => "00000000000000000010000010110101",
			2091 => "00000000000000000010000010110101",
			2092 => "11111110101010110010000010110101",
			2093 => "0000000110000000000001111000110100",
			2094 => "0000000001000000000110000000011000",
			2095 => "0000000110000000001110010100001100",
			2096 => "0000000001000000001110011100000100",
			2097 => "00000000000000000010000101101001",
			2098 => "0000001101000000001100001000000100",
			2099 => "00000000000000000010000101101001",
			2100 => "00000001100101110010000101101001",
			2101 => "0000000010000000001010001000000100",
			2102 => "11111110101101000010000101101001",
			2103 => "0000000111000000001110111100000100",
			2104 => "00000001011100110010000101101001",
			2105 => "00000000000000000010000101101001",
			2106 => "0000000110000000000111101000010100",
			2107 => "0000000111000000000111111000001000",
			2108 => "0000000010000000001110101000000100",
			2109 => "00000000000000000010000101101001",
			2110 => "00000000110000110010000101101001",
			2111 => "0000000110000000000101011100001000",
			2112 => "0000001101000000001110110000000100",
			2113 => "00000000101100100010000101101001",
			2114 => "11111111100011010010000101101001",
			2115 => "11111110100011100010000101101001",
			2116 => "0000000100000000001110010000000100",
			2117 => "00000011100101100010000101101001",
			2118 => "00000000000000000010000101101001",
			2119 => "0000000100000000000001011100010000",
			2120 => "0000000000000000001011010100000100",
			2121 => "11111110011101100010000101101001",
			2122 => "0000001001000000001011001100001000",
			2123 => "0000000011000000000111100000000100",
			2124 => "11111111000010110010000101101001",
			2125 => "00000001110101100010000101101001",
			2126 => "11111110111111110010000101101001",
			2127 => "0000001110000000001001101000001000",
			2128 => "0000000010000000001111010100000100",
			2129 => "11111110101110000010000101101001",
			2130 => "00000011001010000010000101101001",
			2131 => "0000000111000000001110111100001100",
			2132 => "0000000111000000001110111100001000",
			2133 => "0000000101000000001000111100000100",
			2134 => "00000000000000000010000101101001",
			2135 => "11111111011001010010000101101001",
			2136 => "00000000000000000010000101101001",
			2137 => "11111110011101100010000101101001",
			2138 => "0000000110000000000111101000011100",
			2139 => "0000000001000000001110100000011000",
			2140 => "0000001010000000000100101100000100",
			2141 => "00000100010101010010000111101101",
			2142 => "0000001100000000000100010100010000",
			2143 => "0000000011000000000001110100000100",
			2144 => "11111111001011010010000111101101",
			2145 => "0000000010000000000001001000000100",
			2146 => "00000000110100110010000111101101",
			2147 => "0000000011000000000000001100000100",
			2148 => "00000010001000000010000111101101",
			2149 => "00000010110110000010000111101101",
			2150 => "11111110011111000010000111101101",
			2151 => "11111110011010010010000111101101",
			2152 => "0000000111000000001110111100001100",
			2153 => "0000000010000000000011001000000100",
			2154 => "11111110011001110010000111101101",
			2155 => "0000000010000000001001100000000100",
			2156 => "00000001110000100010000111101101",
			2157 => "00000011000010000010000111101101",
			2158 => "0000001100000000000000111000001000",
			2159 => "0000001000000000001110111100000100",
			2160 => "11111111011101110010000111101101",
			2161 => "00000000101000010010000111101101",
			2162 => "0000000100000000001000110100010000",
			2163 => "0000000100000000001000000100000100",
			2164 => "11111110100000000010000111101101",
			2165 => "0000001000000000000001110000000100",
			2166 => "11111110101001110010000111101101",
			2167 => "0000000000000000001000110000000100",
			2168 => "00000111111001100010000111101101",
			2169 => "11111110111100010010000111101101",
			2170 => "11111110011001000010000111101101",
			2171 => "0000000001000000000000011000010100",
			2172 => "0000001100000000000100010100010000",
			2173 => "0000001111000000001010111100000100",
			2174 => "11111111011001110010001001100001",
			2175 => "0000000001000000000000011000000100",
			2176 => "00000001101110100010001001100001",
			2177 => "0000001010000000001001000100000100",
			2178 => "00000000110100010010001001100001",
			2179 => "00000000000000000010001001100001",
			2180 => "11111111000101010010001001100001",
			2181 => "0000001000000000000001110000100100",
			2182 => "0000001100000000000100001000100000",
			2183 => "0000001111000000001010010100010000",
			2184 => "0000001001000000000010001100001000",
			2185 => "0000001101000000000011011100000100",
			2186 => "11111111101110110010001001100001",
			2187 => "00000000101001110010001001100001",
			2188 => "0000001010000000000100111100000100",
			2189 => "00000000000000000010001001100001",
			2190 => "11111110110011000010001001100001",
			2191 => "0000000001000000001101011100001100",
			2192 => "0000000010000000001100010000001000",
			2193 => "0000000100000000001010000100000100",
			2194 => "00000001100011110010001001100001",
			2195 => "00000000000000000010001001100001",
			2196 => "00000001101110100010001001100001",
			2197 => "00000000000000000010001001100001",
			2198 => "11111110101100010010001001100001",
			2199 => "11111110011110110010001001100001",
			2200 => "0000000110000000000111101000011100",
			2201 => "0000000001000000001110100000011000",
			2202 => "0000000110000000001110010100010000",
			2203 => "0000001000000000000111110100000100",
			2204 => "00000011010000010010001011111101",
			2205 => "0000001001000000000010001100000100",
			2206 => "00000001110100110010001011111101",
			2207 => "0000001011000000000100010100000100",
			2208 => "00000001111101110010001011111101",
			2209 => "11111111111100010010001011111101",
			2210 => "0000000010000000001110010000000100",
			2211 => "11111110001110010010001011111101",
			2212 => "00000001101010000010001011111101",
			2213 => "11111110011110010010001011111101",
			2214 => "0000000111000000001110111100001100",
			2215 => "0000000010000000000011001000000100",
			2216 => "11111110011100000010001011111101",
			2217 => "0000001101000000001000111000000100",
			2218 => "00000010010000100010001011111101",
			2219 => "00000001000011000010001011111101",
			2220 => "0000001010000000000011101000010000",
			2221 => "0000000101000000000111110000001100",
			2222 => "0000001100000000001000111000000100",
			2223 => "11111110110001010010001011111101",
			2224 => "0000001001000000001011001100000100",
			2225 => "00000110100011100010001011111101",
			2226 => "11111111011010110010001011111101",
			2227 => "11111110011010100010001011111101",
			2228 => "0000001100000000001010000000010100",
			2229 => "0000001100000000001010000000001100",
			2230 => "0000001100000000000000110000001000",
			2231 => "0000001001000000000110000000000100",
			2232 => "00000000000000000010001011111101",
			2233 => "11111110100000010010001011111101",
			2234 => "11111110011100100010001011111101",
			2235 => "0000000011000000001010000000000100",
			2236 => "00000111100100010010001011111101",
			2237 => "11111111101011010010001011111101",
			2238 => "11111110011001110010001011111101",
			2239 => "0000000110000000000111101000011100",
			2240 => "0000001001000000000110101000011000",
			2241 => "0000000110000000001110010100010000",
			2242 => "0000001111000000001101010100000100",
			2243 => "11111111110101110010001110010001",
			2244 => "0000001000000000000111110100000100",
			2245 => "00000011000110000010001110010001",
			2246 => "0000001001000000000010001100000100",
			2247 => "00000001110010110010001110010001",
			2248 => "00000000111110100010001110010001",
			2249 => "0000000010000000001110010000000100",
			2250 => "11111110010001100010001110010001",
			2251 => "00000001100100110010001110010001",
			2252 => "11111110011111000010001110010001",
			2253 => "0000000111000000001110111100001100",
			2254 => "0000000010000000000011001000000100",
			2255 => "11111110011100110010001110010001",
			2256 => "0000001111000000000110110100000100",
			2257 => "00000010001000110010001110010001",
			2258 => "00000000101111010010001110010001",
			2259 => "0000000100000000000101110000000100",
			2260 => "00000010000011110010001110010001",
			2261 => "0000000100000000000110101100001100",
			2262 => "0000001100000000000100001000001000",
			2263 => "0000000010000000001100010100000100",
			2264 => "11111110101110000010001110010001",
			2265 => "00000101010001010010001110010001",
			2266 => "11111110011011010010001110010001",
			2267 => "0000001100000000001010000000010000",
			2268 => "0000001100000000001010000000001000",
			2269 => "0000001100000000000000110000000100",
			2270 => "11111111011010010010001110010001",
			2271 => "11111110011101010010001110010001",
			2272 => "0000000011000000001010000000000100",
			2273 => "00000101001010010010001110010001",
			2274 => "11111111101111000010001110010001",
			2275 => "11111110011010000010001110010001",
			2276 => "0000000110000000001110010100011100",
			2277 => "0000000010000000000010110100010100",
			2278 => "0000000001000000000110000000001000",
			2279 => "0000000101000000000011011100000100",
			2280 => "00000000000000000010010001001101",
			2281 => "00000000111011010010010001001101",
			2282 => "0000001110000000001000111000000100",
			2283 => "11111111000011100010010001001101",
			2284 => "0000001101000000001110110000000100",
			2285 => "00000000001110100010010001001101",
			2286 => "00000000000000000010010001001101",
			2287 => "0000000001000000001110100000000100",
			2288 => "00000001011100010010010001001101",
			2289 => "00000000000000000010010001001101",
			2290 => "0000000010000000000111010100110000",
			2291 => "0000001111000000000011001000011100",
			2292 => "0000000001000000000000011000001100",
			2293 => "0000000010000000001010001000000100",
			2294 => "11111111010111110010010001001101",
			2295 => "0000000101000000000100011000000100",
			2296 => "00000000110100110010010001001101",
			2297 => "00000000000000000010010001001101",
			2298 => "0000000101000000000100000000000100",
			2299 => "00000000000000000010010001001101",
			2300 => "0000000010000000001100010000000100",
			2301 => "11111110011100100010010001001101",
			2302 => "0000000010000000001100010000000100",
			2303 => "00000000000000000010010001001101",
			2304 => "11111111100101110010010001001101",
			2305 => "0000000110000000001101111100001000",
			2306 => "0000001110000000000111111100000100",
			2307 => "00000001001110110010010001001101",
			2308 => "00000000000000000010010001001101",
			2309 => "0000001111000000001100010000000100",
			2310 => "11111110111000000010010001001101",
			2311 => "0000001111000000001100000000000100",
			2312 => "00000000000000000010010001001101",
			2313 => "11111111110111110010010001001101",
			2314 => "0000001100000000000000001100010000",
			2315 => "0000000110000000001000010000001100",
			2316 => "0000000001000000001101011100001000",
			2317 => "0000000010000000000011000000000100",
			2318 => "00000001101110110010010001001101",
			2319 => "00000000000000000010010001001101",
			2320 => "00000000000000000010010001001101",
			2321 => "00000000000000000010010001001101",
			2322 => "11111110101111100010010001001101",
			2323 => "0000000110000000000111101000100000",
			2324 => "0000001001000000000110101000011100",
			2325 => "0000000010000000000010110100001100",
			2326 => "0000000110000000001011111100001000",
			2327 => "0000000011000000000100000000000100",
			2328 => "00000000010001010010010011100001",
			2329 => "00000001110111100010010011100001",
			2330 => "11111110011001010010010011100001",
			2331 => "0000000110000000001110010100001000",
			2332 => "0000000011000000000000001100000100",
			2333 => "00000001101001010010010011100001",
			2334 => "00000010011011110010010011100001",
			2335 => "0000000001000000000000011000000100",
			2336 => "00000001011010000010010011100001",
			2337 => "11111111000010010010010011100001",
			2338 => "11111110100100000010010011100001",
			2339 => "0000000100000000000101110000000100",
			2340 => "00000110001101110010010011100001",
			2341 => "0000000111000000001110111100001000",
			2342 => "0000000010000000000011001000000100",
			2343 => "11111110100000100010010011100001",
			2344 => "00000001011001100010010011100001",
			2345 => "0000000000000000000111000000010000",
			2346 => "0000001100000000000100001000001100",
			2347 => "0000001111000000000011001000000100",
			2348 => "11111110101011100010010011100001",
			2349 => "0000000001000000001001011000000100",
			2350 => "00000011100000000010010011100001",
			2351 => "11111110110101100010010011100001",
			2352 => "11111110011010110010010011100001",
			2353 => "0000001100000000000000110000001100",
			2354 => "0000001011000000000111111000001000",
			2355 => "0000001011000000001110111100000100",
			2356 => "00000000000000000010010011100001",
			2357 => "11111110111110000010010011100001",
			2358 => "00000000000000000010010011100001",
			2359 => "11111110011001100010010011100001",
			2360 => "0000000110000000001110010100011100",
			2361 => "0000000010000000000010110100010100",
			2362 => "0000000001000000000110000000001000",
			2363 => "0000000101000000000011011100000100",
			2364 => "00000000000000000010010110100101",
			2365 => "00000000111110010010010110100101",
			2366 => "0000000011000000000101101100000100",
			2367 => "11111111000001110010010110100101",
			2368 => "0000001011000000000101101100000100",
			2369 => "00000000001100110010010110100101",
			2370 => "00000000000000000010010110100101",
			2371 => "0000000001000000001110100000000100",
			2372 => "00000001011110010010010110100101",
			2373 => "00000000000000000010010110100101",
			2374 => "0000000010000000000111010100110000",
			2375 => "0000001111000000000011001000011100",
			2376 => "0000000001000000000000011000001100",
			2377 => "0000000010000000001010001000000100",
			2378 => "11111111010010000010010110100101",
			2379 => "0000000101000000000100011000000100",
			2380 => "00000000111001010010010110100101",
			2381 => "00000000000000000010010110100101",
			2382 => "0000000010000000001100010000001000",
			2383 => "0000000101000000000100000000000100",
			2384 => "00000000000000000010010110100101",
			2385 => "11111110011100000010010110100101",
			2386 => "0000000101000000000101101100000100",
			2387 => "00000000000000000010010110100101",
			2388 => "11111111100000010010010110100101",
			2389 => "0000000110000000001101111100001000",
			2390 => "0000001001000000001010011000000100",
			2391 => "00000001010111100010010110100101",
			2392 => "00000000000000000010010110100101",
			2393 => "0000001111000000001100010000000100",
			2394 => "11111110110101100010010110100101",
			2395 => "0000001111000000001100000000000100",
			2396 => "00000000000000000010010110100101",
			2397 => "11111111110101000010010110100101",
			2398 => "0000000111000000000111001000010100",
			2399 => "0000000110000000001000010000010000",
			2400 => "0000000001000000001101011100001100",
			2401 => "0000000010000000000011000000001000",
			2402 => "0000000100000000000011000100000100",
			2403 => "00000001111000010010010110100101",
			2404 => "00000000000000000010010110100101",
			2405 => "00000000000000000010010110100101",
			2406 => "00000000000000000010010110100101",
			2407 => "00000000000000000010010110100101",
			2408 => "11111110101101000010010110100101",
			2409 => "0000000110000000000111101000100000",
			2410 => "0000001001000000000110101000011100",
			2411 => "0000000110000000001011111100001000",
			2412 => "0000000000000000000101000100000100",
			2413 => "00000010101100100010011001011011",
			2414 => "00000001101110110010011001011011",
			2415 => "0000001011000000000111111000001100",
			2416 => "0000000011000000000001110100000100",
			2417 => "00000000000000000010011001011011",
			2418 => "0000000100000000000000100000000100",
			2419 => "00000000000000000010011001011011",
			2420 => "00000001101101100010011001011011",
			2421 => "0000000101000000001101100000000100",
			2422 => "11111111110000010010011001011011",
			2423 => "11111110000111000010011001011011",
			2424 => "11111110011111110010011001011011",
			2425 => "0000001100000000001010000000011000",
			2426 => "0000001000000000000000101000010100",
			2427 => "0000000011000000001010101100000100",
			2428 => "11111110011100110010011001011011",
			2429 => "0000001001000000001110100000001100",
			2430 => "0000000111000000000111111000001000",
			2431 => "0000001101000000000100000000000100",
			2432 => "00000000011101010010011001011011",
			2433 => "00000010000001000010011001011011",
			2434 => "00000000000000000010011001011011",
			2435 => "11111110011100100010011001011011",
			2436 => "00000011100010000010011001011011",
			2437 => "0000000100000000001000110100100000",
			2438 => "0000000100000000001000000100010100",
			2439 => "0000001101000000001110101100010000",
			2440 => "0000000101000000001010010100001000",
			2441 => "0000000011000000000111100000000100",
			2442 => "11111110011011000010011001011011",
			2443 => "11111111111110100010011001011011",
			2444 => "0000000101000000001001010100000100",
			2445 => "00000100101000110010011001011011",
			2446 => "00000000000000000010011001011011",
			2447 => "11111110011010010010011001011011",
			2448 => "0000001010000000001001000100000100",
			2449 => "11111110111010100010011001011011",
			2450 => "0000001000000000001001101000000100",
			2451 => "00000101101000000010011001011011",
			2452 => "11111111111101000010011001011011",
			2453 => "11111110011001010010011001011011",
			2454 => "00000000000000000010011001011101",
			2455 => "00000000000000000010011001100001",
			2456 => "00000000000000000010011001100101",
			2457 => "00000000000000000010011001101001",
			2458 => "00000000000000000010011001101101",
			2459 => "00000000000000000010011001110001",
			2460 => "00000000000000000010011001110101",
			2461 => "00000000000000000010011001111001",
			2462 => "00000000000000000010011001111101",
			2463 => "00000000000000000010011010000001",
			2464 => "00000000000000000010011010000101",
			2465 => "00000000000000000010011010001001",
			2466 => "00000000000000000010011010001101",
			2467 => "00000000000000000010011010010001",
			2468 => "00000000000000000010011010010101",
			2469 => "00000000000000000010011010011001",
			2470 => "00000000000000000010011010011101",
			2471 => "00000000000000000010011010100001",
			2472 => "0000001100000000001010000000000100",
			2473 => "00000000000000000010011010101101",
			2474 => "11111111111110100010011010101101",
			2475 => "0000000111000000001110001100000100",
			2476 => "00000000000100110010011010111001",
			2477 => "00000000000000000010011010111001",
			2478 => "0000000111000000000100010100000100",
			2479 => "00000000000000000010011011000101",
			2480 => "11111111111100010010011011000101",
			2481 => "0000000110000000000001111000000100",
			2482 => "00000000000000000010011011011001",
			2483 => "0000001100000000000011011100000100",
			2484 => "11111111110000110010011011011001",
			2485 => "00000000000000000010011011011001",
			2486 => "0000000111000000001110001100001000",
			2487 => "0000001011000000000000111000000100",
			2488 => "00000000000000000010011011101101",
			2489 => "00000000000011110010011011101101",
			2490 => "00000000000000000010011011101101",
			2491 => "0000000110000000000001111000000100",
			2492 => "00000000000000000010011100000001",
			2493 => "0000000110000000001010011000000100",
			2494 => "11111111100111110010011100000001",
			2495 => "00000000000000000010011100000001",
			2496 => "0000000110000000001101111100001000",
			2497 => "0000000110000000001101011100000100",
			2498 => "00000000000000000010011100010101",
			2499 => "00000000000000110010011100010101",
			2500 => "00000000000000000010011100010101",
			2501 => "0000000110000000001110010100000100",
			2502 => "00000000000000000010011100101001",
			2503 => "0000000110000000001010011000000100",
			2504 => "11111111110010000010011100101001",
			2505 => "00000000000000000010011100101001",
			2506 => "0000000110000000001110010100000100",
			2507 => "00000000000000000010011100111101",
			2508 => "0000000110000000001111000000000100",
			2509 => "11111111111100010010011100111101",
			2510 => "00000000000000000010011100111101",
			2511 => "0000000111000000001110001100001100",
			2512 => "0000001100000000001100110000001000",
			2513 => "0000001011000000000000111000000100",
			2514 => "00000000000000000010011101011001",
			2515 => "00000000000100110010011101011001",
			2516 => "00000000000000000010011101011001",
			2517 => "00000000000000000010011101011001",
			2518 => "0000000111000000001110001100001100",
			2519 => "0000001111000000001001001000000100",
			2520 => "00000000000000000010011101110101",
			2521 => "0000001100000000001100110000000100",
			2522 => "00000000001110010010011101110101",
			2523 => "00000000000000000010011101110101",
			2524 => "00000000000000000010011101110101",
			2525 => "0000000110000000000001111000001100",
			2526 => "0000000110000000001101011100000100",
			2527 => "00000000000000000010011110010001",
			2528 => "0000000110000000001011111100000100",
			2529 => "00000000000111110010011110010001",
			2530 => "00000000000000000010011110010001",
			2531 => "11111111110100000010011110010001",
			2532 => "0000000111000000000110000100001100",
			2533 => "0000001111000000000100011000000100",
			2534 => "00000000000000000010011110101101",
			2535 => "0000000110000000001101111100000100",
			2536 => "00000000010110000010011110101101",
			2537 => "00000000000000000010011110101101",
			2538 => "00000000000000000010011110101101",
			2539 => "0000000110000000001110010100000100",
			2540 => "00000000000000000010011111001001",
			2541 => "0000000110000000001010011000001000",
			2542 => "0000000110000000001110010100000100",
			2543 => "00000000000000000010011111001001",
			2544 => "11111111110100000010011111001001",
			2545 => "00000000000000000010011111001001",
			2546 => "0000000111000000000110000100001100",
			2547 => "0000000110000000001101111100001000",
			2548 => "0000000110000000001001011000000100",
			2549 => "00000000000000000010011111101101",
			2550 => "00000000001101000010011111101101",
			2551 => "00000000000000000010011111101101",
			2552 => "0000000111000000000111001000000100",
			2553 => "11111111111110010010011111101101",
			2554 => "00000000000000000010011111101101",
			2555 => "0000000110000000001011111100001000",
			2556 => "0000000110000000001101011100000100",
			2557 => "00000000000000000010100000010001",
			2558 => "00000000000000110010100000010001",
			2559 => "0000001100000000000000110000000100",
			2560 => "00000000000000000010100000010001",
			2561 => "0000001011000000000000110000000100",
			2562 => "00000000000000000010100000010001",
			2563 => "11111111101111110010100000010001",
			2564 => "0000000110000000001101111100001100",
			2565 => "0000001111000000001001001000000100",
			2566 => "00000000000000000010100000111101",
			2567 => "0000000111000000000110000100000100",
			2568 => "00000000001010110010100000111101",
			2569 => "00000000000000000010100000111101",
			2570 => "0000000100000000000110111100000100",
			2571 => "00000000000000000010100000111101",
			2572 => "0000000110000000001001100100000100",
			2573 => "11111111011011010010100000111101",
			2574 => "00000000000000000010100000111101",
			2575 => "0000001100000000001010000000000100",
			2576 => "00000000000000000010100001100001",
			2577 => "0000001010000000000111101100000100",
			2578 => "00000000000000000010100001100001",
			2579 => "0000001111000000001100010000001000",
			2580 => "0000001011000000001001110100000100",
			2581 => "11111111100010100010100001100001",
			2582 => "00000000000000000010100001100001",
			2583 => "00000000000000000010100001100001",
			2584 => "0000000111000000000110000100010000",
			2585 => "0000001101000000000100000000000100",
			2586 => "00000000000000000010100010000101",
			2587 => "0000000110000000001101111100001000",
			2588 => "0000000110000000001001011000000100",
			2589 => "00000000000000000010100010000101",
			2590 => "00000000000100000010100010000101",
			2591 => "00000000000000000010100010000101",
			2592 => "11111111101001110010100010000101",
			2593 => "0000000110000000001011111100000100",
			2594 => "00000000000000000010100010101001",
			2595 => "0000000100000000001010000100000100",
			2596 => "00000000000000000010100010101001",
			2597 => "0000001100000000000000110000000100",
			2598 => "00000000000000000010100010101001",
			2599 => "0000001011000000000000110000000100",
			2600 => "00000000000000000010100010101001",
			2601 => "11111111100001110010100010101001",
			2602 => "0000001111000000001010111100000100",
			2603 => "00000000000000000010100011001101",
			2604 => "0000001100000000000100001000001100",
			2605 => "0000001111000000001100111000001000",
			2606 => "0000000111000000001110110000000100",
			2607 => "00000000001000010010100011001101",
			2608 => "00000000000000000010100011001101",
			2609 => "00000000000000000010100011001101",
			2610 => "00000000000000000010100011001101",
			2611 => "0000000111000000000110000100010000",
			2612 => "0000000110000000001101111100001100",
			2613 => "0000000110000000001001011000000100",
			2614 => "00000000000000000010100011111001",
			2615 => "0000001011000000000000111000000100",
			2616 => "00000000000000000010100011111001",
			2617 => "00000000010000010010100011111001",
			2618 => "00000000000000000010100011111001",
			2619 => "0000001011000000001001110100000100",
			2620 => "11111111110101010010100011111001",
			2621 => "00000000000000000010100011111001",
			2622 => "0000000111000000000111001000010100",
			2623 => "0000000010000000001100010100001000",
			2624 => "0000000110000000001011111100000100",
			2625 => "00000000000000000010100100100101",
			2626 => "00000000000000000010100100100101",
			2627 => "0000000001000000001101011100001000",
			2628 => "0000000000000000000110110100000100",
			2629 => "00000000011000010010100100100101",
			2630 => "00000000000000000010100100100101",
			2631 => "00000000000000000010100100100101",
			2632 => "00000000000000000010100100100101",
			2633 => "0000000110000000001101111100010000",
			2634 => "0000001111000000001001001000000100",
			2635 => "00000000000000000010100101011001",
			2636 => "0000000111000000000110000100001000",
			2637 => "0000001010000000000111110100000100",
			2638 => "00000000010001110010100101011001",
			2639 => "00000000000000000010100101011001",
			2640 => "00000000000000000010100101011001",
			2641 => "0000001011000000001001110100001000",
			2642 => "0000001100000000000000111000000100",
			2643 => "00000000000000000010100101011001",
			2644 => "11111111011100100010100101011001",
			2645 => "00000000000000000010100101011001",
			2646 => "0000000001000000001110100000010000",
			2647 => "0000001100000000000100000000001100",
			2648 => "0000001101000000000011011100000100",
			2649 => "00000000000000000010100110010101",
			2650 => "0000000101000000001000111000000100",
			2651 => "00000000000000000010100110010101",
			2652 => "00000000011001000010100110010101",
			2653 => "00000000000000000010100110010101",
			2654 => "0000001101000000000010001000001000",
			2655 => "0000000110000000001001011000000100",
			2656 => "00000000000000000010100110010101",
			2657 => "11111111101001100010100110010101",
			2658 => "0000001001000000001011001100000100",
			2659 => "00000000000001110010100110010101",
			2660 => "00000000000000000010100110010101",
			2661 => "0000000110000000001101111100010100",
			2662 => "0000001111000000001110110000000100",
			2663 => "00000000000000000010100111001001",
			2664 => "0000001010000000000111110100001100",
			2665 => "0000000111000000000110000100001000",
			2666 => "0000001010000000000100111100000100",
			2667 => "00000000000000000010100111001001",
			2668 => "00000000011110100010100111001001",
			2669 => "00000000000000000010100111001001",
			2670 => "00000000000000000010100111001001",
			2671 => "0000000110000000001101011000000100",
			2672 => "11111111111110000010100111001001",
			2673 => "00000000000000000010100111001001",
			2674 => "0000001100000000001010000000000100",
			2675 => "00000000000000000010100111110101",
			2676 => "0000000110000000000101011100000100",
			2677 => "00000000000000000010100111110101",
			2678 => "0000000110000000001001100100001100",
			2679 => "0000000110000000001011111100000100",
			2680 => "00000000000000000010100111110101",
			2681 => "0000000111000000001010000000000100",
			2682 => "00000000000000000010100111110101",
			2683 => "11111111110101000010100111110101",
			2684 => "00000000000000000010100111110101",
			2685 => "0000000001000000000000011000010100",
			2686 => "0000001100000000000111111000010000",
			2687 => "0000001001000000001100100000000100",
			2688 => "00000000000000000010101000110001",
			2689 => "0000001011000000000000111000000100",
			2690 => "00000000000000000010101000110001",
			2691 => "0000000001000000001110011100000100",
			2692 => "00000000000000000010101000110001",
			2693 => "00000000010010000010101000110001",
			2694 => "00000000000000000010101000110001",
			2695 => "0000000110000000001010011000001000",
			2696 => "0000000110000000000001111000000100",
			2697 => "00000000000000000010101000110001",
			2698 => "11111111010110110010101000110001",
			2699 => "00000000000000000010101000110001",
			2700 => "0000000010000000001100010100001100",
			2701 => "0000000110000000000001000100000100",
			2702 => "00000000000000000010101001101101",
			2703 => "0000001010000000000111101100000100",
			2704 => "00000000000000000010101001101101",
			2705 => "11111111100100000010101001101101",
			2706 => "0000001100000000000100001000010000",
			2707 => "0000000001000000001101011100001100",
			2708 => "0000000100000000001101001100001000",
			2709 => "0000000010000000000011000000000100",
			2710 => "00000000100010000010101001101101",
			2711 => "00000000000000000010101001101101",
			2712 => "00000000000000000010101001101101",
			2713 => "00000000000000000010101001101101",
			2714 => "00000000000000000010101001101101",
			2715 => "0000000010000000001100010100010000",
			2716 => "0000000110000000000001000100000100",
			2717 => "00000000000000000010101010110001",
			2718 => "0000001010000000000111101100000100",
			2719 => "00000000000000000010101010110001",
			2720 => "0000000001000000001100100000000100",
			2721 => "00000000000000000010101010110001",
			2722 => "11111111011111000010101010110001",
			2723 => "0000000111000000001110110000010000",
			2724 => "0000000001000000001101011100001100",
			2725 => "0000000100000000001101001100001000",
			2726 => "0000000010000000000011000000000100",
			2727 => "00000000101010000010101010110001",
			2728 => "00000000000000000010101010110001",
			2729 => "00000000000000000010101010110001",
			2730 => "00000000000000000010101010110001",
			2731 => "00000000000000000010101010110001",
			2732 => "0000001100000000001010000000010100",
			2733 => "0000001111000000001110110000000100",
			2734 => "00000000000000000010101011111101",
			2735 => "0000001001000000001001111000001100",
			2736 => "0000000111000000000100010100001000",
			2737 => "0000001101000000000100000000000100",
			2738 => "00000000000000000010101011111101",
			2739 => "00000000100011100010101011111101",
			2740 => "00000000000000000010101011111101",
			2741 => "00000000000000000010101011111101",
			2742 => "0000001001000000001100011000001100",
			2743 => "0000000110000000001011111100000100",
			2744 => "00000000000000000010101011111101",
			2745 => "0000000111000000001010000000000100",
			2746 => "00000000000000000010101011111101",
			2747 => "11111111000001010010101011111101",
			2748 => "0000001001000000001011001100000100",
			2749 => "00000000001100110010101011111101",
			2750 => "00000000000000000010101011111101",
			2751 => "0000001001000000000010001100001100",
			2752 => "0000000011000000001010101100000100",
			2753 => "00000000000000000010101101001001",
			2754 => "0000000111000000001100001000000100",
			2755 => "00000000011110000010101101001001",
			2756 => "00000000000000000010101101001001",
			2757 => "0000000110000000001101011000010000",
			2758 => "0000000000000000001001101000000100",
			2759 => "00000000000000000010101101001001",
			2760 => "0000001100000000000000111000000100",
			2761 => "00000000000000000010101101001001",
			2762 => "0000000110000000001011111100000100",
			2763 => "00000000000000000010101101001001",
			2764 => "11111111000101110010101101001001",
			2765 => "0000000001000000001101011100001000",
			2766 => "0000000001000000001101011100000100",
			2767 => "00000000000000000010101101001001",
			2768 => "00000000010101000010101101001001",
			2769 => "00000000000000000010101101001001",
			2770 => "0000000110000000001101111100011100",
			2771 => "0000001111000000000010001000010100",
			2772 => "0000000110000000000001000100001100",
			2773 => "0000000001000000000110000000001000",
			2774 => "0000000001000000001110011100000100",
			2775 => "00000000000000000010101110011101",
			2776 => "00000000001110010010101110011101",
			2777 => "00000000000000000010101110011101",
			2778 => "0000000001000000001100100000000100",
			2779 => "00000000000000000010101110011101",
			2780 => "11111111100100000010101110011101",
			2781 => "0000001011000000001101010100000100",
			2782 => "00000000100111110010101110011101",
			2783 => "00000000000000000010101110011101",
			2784 => "0000000010000000001011111000001000",
			2785 => "0000001011000000001001110100000100",
			2786 => "11111111000110110010101110011101",
			2787 => "00000000000000000010101110011101",
			2788 => "0000001100000000000011011100000100",
			2789 => "00000000011010100010101110011101",
			2790 => "00000000000000000010101110011101",
			2791 => "0000000001000000000110000000011000",
			2792 => "0000001011000000001110111100000100",
			2793 => "00000000000000000010101111011001",
			2794 => "0000000111000000000000101000010000",
			2795 => "0000000011000000000010111100000100",
			2796 => "00000000000000000010101111011001",
			2797 => "0000001100000000001010000000000100",
			2798 => "00000000000000000010101111011001",
			2799 => "0000000101000000001000111100000100",
			2800 => "00000000000000000010101111011001",
			2801 => "00000000010010100010101111011001",
			2802 => "00000000000000000010101111011001",
			2803 => "0000000000000000001001101000000100",
			2804 => "00000000000000000010101111011001",
			2805 => "11111111010011110010101111011001",
			2806 => "0000000110000000001110010100001100",
			2807 => "0000000110000000001001011000000100",
			2808 => "00000000000000000010110000100101",
			2809 => "0000001100000000001000111000000100",
			2810 => "00000000011101110010110000100101",
			2811 => "00000000000000000010110000100101",
			2812 => "0000001100000000000011011100001000",
			2813 => "0000000000000000001000011000000100",
			2814 => "11111111010000000010110000100101",
			2815 => "00000000000000000010110000100101",
			2816 => "0000001100000000000100001000010000",
			2817 => "0000001110000000001000001100001100",
			2818 => "0000000000000000000111000000001000",
			2819 => "0000000000000000001011010100000100",
			2820 => "00000000000000000010110000100101",
			2821 => "00000000100011000010110000100101",
			2822 => "00000000000000000010110000100101",
			2823 => "00000000000000000010110000100101",
			2824 => "00000000000000000010110000100101",
			2825 => "0000000001000000001110100000010100",
			2826 => "0000001111000000001011000000000100",
			2827 => "00000000000000000010110001111001",
			2828 => "0000001100000000000100010100001100",
			2829 => "0000000110000000000111101000000100",
			2830 => "00000000111001010010110001111001",
			2831 => "0000000110000000001010011000000100",
			2832 => "00000000000000000010110001111001",
			2833 => "00000000000001000010110001111001",
			2834 => "00000000000000000010110001111001",
			2835 => "0000000101000000000000011100001000",
			2836 => "0000001000000000000111110100000100",
			2837 => "00000000000000000010110001111001",
			2838 => "11111110111001110010110001111001",
			2839 => "0000001001000000001011001100001100",
			2840 => "0000001100000000000100001000001000",
			2841 => "0000000101000000000111110000000100",
			2842 => "00000000010111000010110001111001",
			2843 => "00000000000000000010110001111001",
			2844 => "00000000000000000010110001111001",
			2845 => "11111111110011100010110001111001",
			2846 => "0000001011000000001010111000011000",
			2847 => "0000001100000000001100110000010100",
			2848 => "0000000101000000000100000000000100",
			2849 => "00000000000000000010110010101101",
			2850 => "0000000111000000001110001100001100",
			2851 => "0000000111000000000000110000000100",
			2852 => "00000000000000000010110010101101",
			2853 => "0000001001000000001100100000000100",
			2854 => "00000000000000000010110010101101",
			2855 => "00000000001000110010110010101101",
			2856 => "00000000000000000010110010101101",
			2857 => "00000000000000000010110010101101",
			2858 => "00000000000000000010110010101101",
			2859 => "0000001010000000001000100100011000",
			2860 => "0000001001000000001011001100010100",
			2861 => "0000001111000000001011011100001000",
			2862 => "0000000001000000000110000000000100",
			2863 => "00000000101001100010110100000001",
			2864 => "11111111010100010010110100000001",
			2865 => "0000000000000000001100011100000100",
			2866 => "00000000000000000010110100000001",
			2867 => "0000000101000000001010010100000100",
			2868 => "00000001000000100010110100000001",
			2869 => "00000000000000000010110100000001",
			2870 => "11111111011010000010110100000001",
			2871 => "0000000110000000000001111000010000",
			2872 => "0000000100000000001111100000000100",
			2873 => "11111111111011000010110100000001",
			2874 => "0000001100000000000100010100001000",
			2875 => "0000000011000000000001110100000100",
			2876 => "00000000000000000010110100000001",
			2877 => "00000000110010110010110100000001",
			2878 => "00000000000000000010110100000001",
			2879 => "11111110100110000010110100000001",
			2880 => "0000001000000000000101000100011000",
			2881 => "0000000111000000001110001100010000",
			2882 => "0000001111000000001110110000000100",
			2883 => "00000000000000000010110101100101",
			2884 => "0000001000000000000000001000000100",
			2885 => "00000000000000000010110101100101",
			2886 => "0000001000000000000101000100000100",
			2887 => "00000000101110010010110101100101",
			2888 => "00000000000000000010110101100101",
			2889 => "0000000110000000001001100100000100",
			2890 => "11111111110000010010110101100101",
			2891 => "00000000000000000010110101100101",
			2892 => "0000000110000000001110010100001000",
			2893 => "0000000101000000001101100000000100",
			2894 => "00000000010111010010110101100101",
			2895 => "00000000000000000010110101100101",
			2896 => "0000000000000000000111000000000100",
			2897 => "00000000000000000010110101100101",
			2898 => "0000001001000000000110000000000100",
			2899 => "00000000000000000010110101100101",
			2900 => "0000000101000000000100000000000100",
			2901 => "00000000000000000010110101100101",
			2902 => "0000000111000000001010000000000100",
			2903 => "00000000000000000010110101100101",
			2904 => "11111110110100000010110101100101",
			2905 => "0000000010000000001100010100010100",
			2906 => "0000000110000000000001111000010000",
			2907 => "0000000010000000000111010000000100",
			2908 => "00000000000000000010110110111001",
			2909 => "0000000110000000001011111100001000",
			2910 => "0000000001000000001110100000000100",
			2911 => "00000000010100110010110110111001",
			2912 => "00000000000000000010110110111001",
			2913 => "00000000000000000010110110111001",
			2914 => "11111111011101010010110110111001",
			2915 => "0000000001000000001101011100010100",
			2916 => "0000001100000000000100001000010000",
			2917 => "0000001001000000001100100000000100",
			2918 => "00000000000000000010110110111001",
			2919 => "0000000100000000001101001100001000",
			2920 => "0000000010000000000011000000000100",
			2921 => "00000000101000110010110110111001",
			2922 => "00000000000000000010110110111001",
			2923 => "00000000000000000010110110111001",
			2924 => "00000000000000000010110110111001",
			2925 => "00000000000000000010110110111001",
			2926 => "0000000110000000001110010100010000",
			2927 => "0000001111000000001110110000000100",
			2928 => "00000000000000000010111000100101",
			2929 => "0000000001000000001110100000001000",
			2930 => "0000000100000000000100100000000100",
			2931 => "00000001000111110010111000100101",
			2932 => "00000000000000000010111000100101",
			2933 => "00000000000000000010111000100101",
			2934 => "0000000100000000000000010000001100",
			2935 => "0000000111000000000101101100000100",
			2936 => "00000000000000000010111000100101",
			2937 => "0000001100000000001110001100000100",
			2938 => "00000000110110110010111000100101",
			2939 => "00000000000000000010111000100101",
			2940 => "0000001001000000000110000000010000",
			2941 => "0000001001000000001100100000000100",
			2942 => "00000000000000000010111000100101",
			2943 => "0000001100000000000111111000001000",
			2944 => "0000000011000000000001110100000100",
			2945 => "00000000000000000010111000100101",
			2946 => "00000000101001100010111000100101",
			2947 => "00000000000000000010111000100101",
			2948 => "0000001011000000001001110100000100",
			2949 => "11111110101011010010111000100101",
			2950 => "0000001011000000000001101000000100",
			2951 => "00000000000000000010111000100101",
			2952 => "11111111110100010010111000100101",
			2953 => "0000001000000000000001110000011100",
			2954 => "0000001100000000000100001000011000",
			2955 => "0000001111000000001110110000000100",
			2956 => "00000000000000000010111001111001",
			2957 => "0000000001000000001001011000010000",
			2958 => "0000001000000000000000001000000100",
			2959 => "00000000000000000010111001111001",
			2960 => "0000000101000000001001010100001000",
			2961 => "0000000000000000000111000000000100",
			2962 => "00000000100011010010111001111001",
			2963 => "00000000000000000010111001111001",
			2964 => "00000000000000000010111001111001",
			2965 => "00000000000000000010111001111001",
			2966 => "00000000000000000010111001111001",
			2967 => "0000000110000000001110010100000100",
			2968 => "00000000000000000010111001111001",
			2969 => "0000001100000000000000110000000100",
			2970 => "00000000000000000010111001111001",
			2971 => "0000001001000000000110000000000100",
			2972 => "00000000000000000010111001111001",
			2973 => "11111111000101110010111001111001",
			2974 => "0000001001000000001100110100010000",
			2975 => "0000001111000000001010111100000100",
			2976 => "00000000000000000010111011100101",
			2977 => "0000001011000000001000111100001000",
			2978 => "0000001011000000000000111000000100",
			2979 => "00000000000000000010111011100101",
			2980 => "00000000110010110010111011100101",
			2981 => "00000000000000000010111011100101",
			2982 => "0000001000000000001100000100100000",
			2983 => "0000001111000000001010010100010000",
			2984 => "0000001001000000000010001100000100",
			2985 => "00000000000000000010111011100101",
			2986 => "0000000100000000001100001100001000",
			2987 => "0000000110000000001001011000000100",
			2988 => "00000000000000000010111011100101",
			2989 => "11111111100000110010111011100101",
			2990 => "00000000000000000010111011100101",
			2991 => "0000000111000000001110001100000100",
			2992 => "00000000100111010010111011100101",
			2993 => "0000000110000000001001100100001000",
			2994 => "0000001111000000001100010100000100",
			2995 => "00000000000000000010111011100101",
			2996 => "11111111010111000010111011100101",
			2997 => "00000000000000000010111011100101",
			2998 => "0000001010000000001000100100000100",
			2999 => "00000000000000000010111011100101",
			3000 => "11111110111110110010111011100101",
			3001 => "0000000110000000001101111100011100",
			3002 => "0000000111000000000110000100011000",
			3003 => "0000000110000000001101011100000100",
			3004 => "00000000000000000010111100100001",
			3005 => "0000001010000000000111110100010000",
			3006 => "0000000101000000001000111100000100",
			3007 => "00000000000000000010111100100001",
			3008 => "0000001010000000000011101000001000",
			3009 => "0000000100000000000110110100000100",
			3010 => "00000000000000000010111100100001",
			3011 => "00000000011011100010111100100001",
			3012 => "00000000000000000010111100100001",
			3013 => "00000000000000000010111100100001",
			3014 => "00000000000000000010111100100001",
			3015 => "11111111101100110010111100100001",
			3016 => "0000000110000000000001111000101000",
			3017 => "0000000001000000000110000000001100",
			3018 => "0000001111000000001010111100000100",
			3019 => "00000000000000000010111110101101",
			3020 => "0000001100000000000111111000000100",
			3021 => "00000001010101110010111110101101",
			3022 => "00000000000000000010111110101101",
			3023 => "0000001110000000001000111000001100",
			3024 => "0000000110000000000001000100000100",
			3025 => "00000000000000000010111110101101",
			3026 => "0000000100000000000101010100000100",
			3027 => "11111110101111000010111110101101",
			3028 => "00000000000000000010111110101101",
			3029 => "0000000000000000001100011100000100",
			3030 => "00000000000000000010111110101101",
			3031 => "0000001110000000001001110000000100",
			3032 => "00000000000000000010111110101101",
			3033 => "0000000001000000000111100100000100",
			3034 => "00000001001010010010111110101101",
			3035 => "00000000000000000010111110101101",
			3036 => "0000000000000000000111000000010100",
			3037 => "0000000100000000000110111000001100",
			3038 => "0000001110000000001001010000001000",
			3039 => "0000000011000000000111100000000100",
			3040 => "11111111010100000010111110101101",
			3041 => "00000000101110110010111110101101",
			3042 => "11111110110000000010111110101101",
			3043 => "0000001100000000000000001100000100",
			3044 => "00000001001111100010111110101101",
			3045 => "11111111101001100010111110101101",
			3046 => "0000000001000000001100100000001000",
			3047 => "0000001001000000000000011000000100",
			3048 => "11111111110000000010111110101101",
			3049 => "00000000000000000010111110101101",
			3050 => "11111110011110010010111110101101",
			3051 => "0000001001000000001100110100010000",
			3052 => "0000001111000000001010111100000100",
			3053 => "00000000000000000011000000100001",
			3054 => "0000001011000000001000111100001000",
			3055 => "0000001011000000000000111000000100",
			3056 => "00000000000000000011000000100001",
			3057 => "00000000101111010011000000100001",
			3058 => "00000000000000000011000000100001",
			3059 => "0000001000000000001100000100100100",
			3060 => "0000000100000000000110111000011000",
			3061 => "0000000100000000001010000100001100",
			3062 => "0000001111000000001010010100000100",
			3063 => "00000000000000000011000000100001",
			3064 => "0000000101000000000110110100000100",
			3065 => "00000000100101000011000000100001",
			3066 => "00000000000000000011000000100001",
			3067 => "0000001001000000001001111000000100",
			3068 => "00000000000000000011000000100001",
			3069 => "0000001111000000001010000100000100",
			3070 => "11111111001001010011000000100001",
			3071 => "00000000000000000011000000100001",
			3072 => "0000001100000000001110001100001000",
			3073 => "0000001111000000000001001000000100",
			3074 => "00000000000000000011000000100001",
			3075 => "00000000100110010011000000100001",
			3076 => "00000000000000000011000000100001",
			3077 => "0000001010000000001000100100000100",
			3078 => "00000000000000000011000000100001",
			3079 => "11111111000001010011000000100001",
			3080 => "0000001100000000001010000000100000",
			3081 => "0000001001000000001100110100010000",
			3082 => "0000001111000000001010111100000100",
			3083 => "11111111011010010011000010101101",
			3084 => "0000000100000000001111110000001000",
			3085 => "0000000110000000001101111100000100",
			3086 => "00000001100000110011000010101101",
			3087 => "00000000000000000011000010101101",
			3088 => "00000100000010100011000010101101",
			3089 => "0000001110000000001011000100001000",
			3090 => "0000000001000000000000011000000100",
			3091 => "00000000000000000011000010101101",
			3092 => "11111110101011010011000010101101",
			3093 => "0000000110000000000111101000000100",
			3094 => "00000001010110100011000010101101",
			3095 => "11111111101111100011000010101101",
			3096 => "0000000000000000000111000000011100",
			3097 => "0000001100000000000100001000011000",
			3098 => "0000001100000000001000111000001100",
			3099 => "0000001001000000001001111000001000",
			3100 => "0000001101000000001100110000000100",
			3101 => "00000000000000000011000010101101",
			3102 => "00000000111011110011000010101101",
			3103 => "11111110111111010011000010101101",
			3104 => "0000001000000000000111110100000100",
			3105 => "00000000000000000011000010101101",
			3106 => "0000000001000000001001011000000100",
			3107 => "00000001101001000011000010101101",
			3108 => "00000000000000000011000010101101",
			3109 => "11111110101000110011000010101101",
			3110 => "0000000110000000001011111100000100",
			3111 => "00000000000000000011000010101101",
			3112 => "0000001011000000001010000000000100",
			3113 => "00000000000000000011000010101101",
			3114 => "11111110011011100011000010101101",
			3115 => "0000000001000000000110000000011100",
			3116 => "0000001111000000001110110000001000",
			3117 => "0000000110000000000101011100000100",
			3118 => "00000000000000000011000100111001",
			3119 => "11111111100010100011000100111001",
			3120 => "0000001100000000000100010100010000",
			3121 => "0000000001000000000000011000001000",
			3122 => "0000001101000000000100000000000100",
			3123 => "00000000000000000011000100111001",
			3124 => "00000001100111110011000100111001",
			3125 => "0000001101000000000011011100000100",
			3126 => "11111111111010110011000100111001",
			3127 => "00000000110001110011000100111001",
			3128 => "00000000000000000011000100111001",
			3129 => "0000000000000000000111000000011100",
			3130 => "0000001010000000001000100100010100",
			3131 => "0000001100000000001000111000010000",
			3132 => "0000000000000000001001101000001000",
			3133 => "0000001111000000000110100100000100",
			3134 => "00000000000000000011000100111001",
			3135 => "00000000110101110011000100111001",
			3136 => "0000001101000000001100101100000100",
			3137 => "00000000000000000011000100111001",
			3138 => "11111111011010000011000100111001",
			3139 => "11111110110101010011000100111001",
			3140 => "0000001100000000000000001100000100",
			3141 => "00000001001111100011000100111001",
			3142 => "11111111110011110011000100111001",
			3143 => "0000000101000000001001110000000100",
			3144 => "00000000000000000011000100111001",
			3145 => "0000001001000000000010001100000100",
			3146 => "00000000000000000011000100111001",
			3147 => "0000001010000000000011101000000100",
			3148 => "00000000000000000011000100111001",
			3149 => "11111110100000100011000100111001",
			3150 => "0000001010000000001000100100100000",
			3151 => "0000001001000000001011001100011100",
			3152 => "0000001111000000001011011100001000",
			3153 => "0000000001000000000110000000000100",
			3154 => "00000000100101100011000110110101",
			3155 => "11111111011001010011000110110101",
			3156 => "0000000000000000001100011100000100",
			3157 => "00000000000000000011000110110101",
			3158 => "0000000101000000001010010100001100",
			3159 => "0000001010000000000011101000000100",
			3160 => "00000001000000100011000110110101",
			3161 => "0000001000000000000101000100000100",
			3162 => "00000000000000000011000110110101",
			3163 => "00000000001110010011000110110101",
			3164 => "00000000000000000011000110110101",
			3165 => "11111111011110010011000110110101",
			3166 => "0000001001000000001100110100011000",
			3167 => "0000000110000000000001111000010000",
			3168 => "0000000111000000000100010100001100",
			3169 => "0000001111000000001101010100000100",
			3170 => "00000000000000000011000110110101",
			3171 => "0000000100000000001101110100000100",
			3172 => "00000000000000000011000110110101",
			3173 => "00000000101010010011000110110101",
			3174 => "00000000000000000011000110110101",
			3175 => "0000001111000000001111011100000100",
			3176 => "11111111111111010011000110110101",
			3177 => "00000000000000000011000110110101",
			3178 => "0000000101000000000100000000000100",
			3179 => "00000000000000000011000110110101",
			3180 => "11111110100110100011000110110101",
			3181 => "0000000110000000000111101000011100",
			3182 => "0000000001000000001110100000011000",
			3183 => "0000000110000000001110010100010000",
			3184 => "0000001100000000000100010100001100",
			3185 => "0000001111000000000111001000000100",
			3186 => "00000000011001110011001001000001",
			3187 => "0000001001000000001001111000000100",
			3188 => "00000001111001110011001001000001",
			3189 => "00000000000000000011001001000001",
			3190 => "00000011101101010011001001000001",
			3191 => "0000000010000000001110010000000100",
			3192 => "11111110001011010011001001000001",
			3193 => "00000001101111100011001001000001",
			3194 => "11111110011101100011001001000001",
			3195 => "0000000111000000001110111100001100",
			3196 => "0000000010000000000011001000000100",
			3197 => "11111110011011010011001001000001",
			3198 => "0000001111000000000110110100000100",
			3199 => "00000010011011000011001001000001",
			3200 => "00000001001001110011001001000001",
			3201 => "0000001010000000000011101000010000",
			3202 => "0000001011000000000110100100001100",
			3203 => "0000001011000000000100001000000100",
			3204 => "11111110110001110011001001000001",
			3205 => "0000000010000000001100000000000100",
			3206 => "00001001101101000011001001000001",
			3207 => "11111111100110000011001001000001",
			3208 => "11111110011010010011001001000001",
			3209 => "0000001100000000000000110000001100",
			3210 => "0000000011000000000011010000001000",
			3211 => "0000000011000000000001110100000100",
			3212 => "11111110101110000011001001000001",
			3213 => "00000001011101010011001001000001",
			3214 => "11111110011101010011001001000001",
			3215 => "11111110011010010011001001000001",
			3216 => "0000000110000000000001111000100100",
			3217 => "0000000001000000000110000000010000",
			3218 => "0000001111000000001010111100000100",
			3219 => "11111111001001000011001011010101",
			3220 => "0000000111000000000000101000001000",
			3221 => "0000000110000000001110010100000100",
			3222 => "00000001100101010011001011010101",
			3223 => "00000000101011010011001011010101",
			3224 => "00000000000000000011001011010101",
			3225 => "0000001111000000000100010000001000",
			3226 => "0000001001000000000010001100000100",
			3227 => "00000000000000000011001011010101",
			3228 => "11111110100100010011001011010101",
			3229 => "0000000011000000000101110100001000",
			3230 => "0000001111000000001010010100000100",
			3231 => "00000000000000000011001011010101",
			3232 => "00000001111011000011001011010101",
			3233 => "11111111011111100011001011010101",
			3234 => "0000000100000000000110101100001100",
			3235 => "0000000000000000001011010100000100",
			3236 => "11111110101101110011001011010101",
			3237 => "0000001110000000001110101000000100",
			3238 => "00000000000000000011001011010101",
			3239 => "00000001001000000011001011010101",
			3240 => "0000000111000000001110111100011000",
			3241 => "0000001001000000001110100000010100",
			3242 => "0000001101000000001000111100001100",
			3243 => "0000000111000000001110111100001000",
			3244 => "0000001101000000000100000000000100",
			3245 => "11111111110011100011001011010101",
			3246 => "00000000000000000011001011010101",
			3247 => "00000000000000000011001011010101",
			3248 => "0000000001000000001110011100000100",
			3249 => "00000000000000000011001011010101",
			3250 => "00000000100000100011001011010101",
			3251 => "11111111001001110011001011010101",
			3252 => "11111110011111100011001011010101",
			3253 => "0000000001000000000000011000010000",
			3254 => "0000001111000000001110110000000100",
			3255 => "00000000000000000011001101011001",
			3256 => "0000000101000000001100101000001000",
			3257 => "0000001101000000000100000000000100",
			3258 => "00000000000000000011001101011001",
			3259 => "00000001000011010011001101011001",
			3260 => "00000000000000000011001101011001",
			3261 => "0000000000000000001000110000101000",
			3262 => "0000000100000000000110111000011100",
			3263 => "0000000100000000001010000100010000",
			3264 => "0000001111000000001011000000000100",
			3265 => "00000000000000000011001101011001",
			3266 => "0000000111000000000110000100001000",
			3267 => "0000001000000000000000001000000100",
			3268 => "00000000000000000011001101011001",
			3269 => "00000000110101010011001101011001",
			3270 => "00000000000000000011001101011001",
			3271 => "0000000111000000000111001000001000",
			3272 => "0000000001000000001110100000000100",
			3273 => "00000000000000000011001101011001",
			3274 => "11111110111010000011001101011001",
			3275 => "00000000000000000011001101011001",
			3276 => "0000001100000000001110001100001000",
			3277 => "0000000000000000001000101100000100",
			3278 => "00000000110111100011001101011001",
			3279 => "00000000000000000011001101011001",
			3280 => "00000000000000000011001101011001",
			3281 => "0000000110000000001011111100000100",
			3282 => "00000000000000000011001101011001",
			3283 => "0000000101000000000100000000000100",
			3284 => "00000000000000000011001101011001",
			3285 => "11111110101101100011001101011001",
			3286 => "0000000001000000000000011000010100",
			3287 => "0000000001000000001110011100000100",
			3288 => "00000000000000000011001111001101",
			3289 => "0000001100000000000111111000001100",
			3290 => "0000001111000000001010111100000100",
			3291 => "00000000000000000011001111001101",
			3292 => "0000001101000000000100000000000100",
			3293 => "00000000000000000011001111001101",
			3294 => "00000001011100010011001111001101",
			3295 => "00000000000000000011001111001101",
			3296 => "0000001000000000000001110000100000",
			3297 => "0000001100000000000100001000011100",
			3298 => "0000001110000000000100000000001000",
			3299 => "0000000100000000001000110100000100",
			3300 => "11111111001111000011001111001101",
			3301 => "00000000000000000011001111001101",
			3302 => "0000000001000000001101011100010000",
			3303 => "0000000111000000000111001000001000",
			3304 => "0000000110000000000001111000000100",
			3305 => "00000000111101010011001111001101",
			3306 => "11111111011110110011001111001101",
			3307 => "0000000001000000001101011100000100",
			3308 => "00000000000000000011001111001101",
			3309 => "00000001010000100011001111001101",
			3310 => "00000000000000000011001111001101",
			3311 => "11111111010000010011001111001101",
			3312 => "0000000110000000001110010100000100",
			3313 => "00000000000000000011001111001101",
			3314 => "11111110100001010011001111001101",
			3315 => "0000000001000000000000011000010000",
			3316 => "0000001111000000001011000000000100",
			3317 => "00000000000000000011010001010001",
			3318 => "0000000101000000001100101000001000",
			3319 => "0000001101000000000100000000000100",
			3320 => "00000000000000000011010001010001",
			3321 => "00000001001001000011010001010001",
			3322 => "00000000000000000011010001010001",
			3323 => "0000000000000000001000110000101000",
			3324 => "0000001001000000001011001100011100",
			3325 => "0000001001000000001100011000010100",
			3326 => "0000000110000000000001111000010000",
			3327 => "0000001110000000001011000100001000",
			3328 => "0000001101000000000110000100000100",
			3329 => "11111111110100100011010001010001",
			3330 => "00000000000000000011010001010001",
			3331 => "0000000101000000000110100100000100",
			3332 => "00000000101110010011010001010001",
			3333 => "00000000000000000011010001010001",
			3334 => "11111111001101010011010001010001",
			3335 => "0000001101000000001110101100000100",
			3336 => "00000000111000000011010001010001",
			3337 => "00000000000000000011010001010001",
			3338 => "0000001010000000001001000100000100",
			3339 => "11111111001100000011010001010001",
			3340 => "0000001001000000001001111100000100",
			3341 => "00000000001100110011010001010001",
			3342 => "00000000000000000011010001010001",
			3343 => "0000000110000000001011111100000100",
			3344 => "00000000000000000011010001010001",
			3345 => "0000000101000000000100000000000100",
			3346 => "00000000000000000011010001010001",
			3347 => "11111110101011110011010001010001",
			3348 => "0000000110000000000111101000100000",
			3349 => "0000001001000000001001111000011100",
			3350 => "0000001111000000001101010100001000",
			3351 => "0000000111000000000000110000000100",
			3352 => "00000000000010010011010011011101",
			3353 => "11111110011010100011010011011101",
			3354 => "0000000010000000000101110100000100",
			3355 => "00000100001001000011010011011101",
			3356 => "0000001100000000000111111000001100",
			3357 => "0000000110000000001110010100000100",
			3358 => "00000010000010000011010011011101",
			3359 => "0000000010000000001110010000000100",
			3360 => "11111110101001110011010011011101",
			3361 => "00000010000010000011010011011101",
			3362 => "11111110100100110011010011011101",
			3363 => "11111110011011000011010011011101",
			3364 => "0000000111000000001110111100001100",
			3365 => "0000000010000000000011001000000100",
			3366 => "11111110011010010011010011011101",
			3367 => "0000001111000000000110110100000100",
			3368 => "00000010110011100011010011011101",
			3369 => "00000001010110010011010011011101",
			3370 => "0000001100000000000000111000001000",
			3371 => "0000001000000000001110111100000100",
			3372 => "11111111100011010011010011011101",
			3373 => "00000000100010000011010011011101",
			3374 => "0000000100000000001000110100010000",
			3375 => "0000000100000000001000000100000100",
			3376 => "11111110100001100011010011011101",
			3377 => "0000001000000000000001110000000100",
			3378 => "11111110101100100011010011011101",
			3379 => "0000001000000000001100000100000100",
			3380 => "00000101100010110011010011011101",
			3381 => "11111110111101000011010011011101",
			3382 => "11111110011001100011010011011101",
			3383 => "0000000001000000000000011000011000",
			3384 => "0000001100000000000100010100010100",
			3385 => "0000000011000000001010101100001000",
			3386 => "0000000111000000000000110000000100",
			3387 => "00000000000000000011010101011001",
			3388 => "11111111011101110011010101011001",
			3389 => "0000000100000000001111110000001000",
			3390 => "0000000010000000001110101000000100",
			3391 => "00000000001011110011010101011001",
			3392 => "00000001011010110011010101011001",
			3393 => "00000011011010100011010101011001",
			3394 => "11111110111111100011010101011001",
			3395 => "0000001000000000000001110000100100",
			3396 => "0000001100000000000100001000100000",
			3397 => "0000001110000000001101010100001100",
			3398 => "0000001001000000001001111000001000",
			3399 => "0000000011000000000000101000000100",
			3400 => "11111111000110100011010101011001",
			3401 => "00000001000010000011010101011001",
			3402 => "11111110110100110011010101011001",
			3403 => "0000000001000000001101011100010000",
			3404 => "0000000000000000000110001000001000",
			3405 => "0000001011000000000001111100000100",
			3406 => "00000001100001000011010101011001",
			3407 => "11111110110110110011010101011001",
			3408 => "0000000010000000001110010000000100",
			3409 => "00000000000000000011010101011001",
			3410 => "00000001110101100011010101011001",
			3411 => "00000000000000000011010101011001",
			3412 => "11111110101010000011010101011001",
			3413 => "11111110011101110011010101011001",
			3414 => "0000000110000000001110010100100000",
			3415 => "0000000101000000000100011000011100",
			3416 => "0000000010000000000001001000001100",
			3417 => "0000000011000000000100000000000100",
			3418 => "11111110100111000011010111111101",
			3419 => "0000000001000000001110100000000100",
			3420 => "00000001011100110011010111111101",
			3421 => "00000000000000000011010111111101",
			3422 => "0000000001000000001110100000001100",
			3423 => "0000000001000000000110000000000100",
			3424 => "00000001101010100011010111111101",
			3425 => "0000000110000000001011111100000100",
			3426 => "00000001101000000011010111111101",
			3427 => "00000000000000000011010111111101",
			3428 => "11111111101011100011010111111101",
			3429 => "11111110100100100011010111111101",
			3430 => "0000001001000000001110100000010000",
			3431 => "0000000010000000001000101000001100",
			3432 => "0000000100000000001111110100001000",
			3433 => "0000000010000000001110010000000100",
			3434 => "11111110101001110011010111111101",
			3435 => "00000001100010010011010111111101",
			3436 => "11111110100000100011010111111101",
			3437 => "00001000111011100011010111111101",
			3438 => "0000000100000000000110101100010000",
			3439 => "0000001000000000000110011000000100",
			3440 => "11111110011111100011010111111101",
			3441 => "0000001110000000001110101000000100",
			3442 => "11111111001111000011010111111101",
			3443 => "0000001001000000001001111100000100",
			3444 => "00000010100001000011010111111101",
			3445 => "11111111101110110011010111111101",
			3446 => "0000001000000000000001110000010000",
			3447 => "0000001001000000000100111100001100",
			3448 => "0000000010000000001000001100001000",
			3449 => "0000000100000000000101000000000100",
			3450 => "11111110100010110011010111111101",
			3451 => "00000000000000000011010111111101",
			3452 => "00000010000101110011010111111101",
			3453 => "11111110011101100011010111111101",
			3454 => "11111110011001110011010111111101",
			3455 => "0000000110000000000001111000101100",
			3456 => "0000000010000000000101001000100000",
			3457 => "0000001010000000000011101000011000",
			3458 => "0000001111000000001110110000000100",
			3459 => "11111111010011100011011010010001",
			3460 => "0000000001000000000111100100010000",
			3461 => "0000001010000000001010100000001000",
			3462 => "0000001000000000000000001000000100",
			3463 => "00000000000000000011011010010001",
			3464 => "00000001101101100011011010010001",
			3465 => "0000000111000000000100010100000100",
			3466 => "00000000111101100011011010010001",
			3467 => "11111111011010010011011010010001",
			3468 => "11111111110101100011011010010001",
			3469 => "0000000110000000001011111100000100",
			3470 => "00000000001011010011011010010001",
			3471 => "11111110100101000011011010010001",
			3472 => "0000000111000000000000101000001000",
			3473 => "0000000001000000001110100000000100",
			3474 => "00000001100100000011011010010001",
			3475 => "00000000000000000011011010010001",
			3476 => "11111111001100100011011010010001",
			3477 => "0000000010000000001110110100000100",
			3478 => "11111110011011110011011010010001",
			3479 => "0000001100000000000100001000011000",
			3480 => "0000000000000000000111000000010000",
			3481 => "0000001011000000001001110100001000",
			3482 => "0000001111000000000010000100000100",
			3483 => "00000000100011000011011010010001",
			3484 => "11111111011010100011011010010001",
			3485 => "0000001011000000000001101000000100",
			3486 => "00000001010010110011011010010001",
			3487 => "00000000000000000011011010010001",
			3488 => "0000001011000000001011000100000100",
			3489 => "00000000100011000011011010010001",
			3490 => "11111110101011100011011010010001",
			3491 => "11111110100010110011011010010001",
			3492 => "0000000110000000000111101000100100",
			3493 => "0000000001000000001110100000011000",
			3494 => "0000000010000000000101110100000100",
			3495 => "00000110110111010011011100110101",
			3496 => "0000000001000000001110011100000100",
			3497 => "11111110011101010011011100110101",
			3498 => "0000000010000000000111100000001000",
			3499 => "0000000110000000001110010100000100",
			3500 => "00000010111001100011011100110101",
			3501 => "11111101110011110011011100110101",
			3502 => "0000000011000000000000001100000100",
			3503 => "00000010110000000011011100110101",
			3504 => "00000011110010010011011100110101",
			3505 => "0000000001000000001110100000001000",
			3506 => "0000000001000000001110100000000100",
			3507 => "11111110110010100011011100110101",
			3508 => "00000000101110000011011100110101",
			3509 => "11111110011001110011011100110101",
			3510 => "0000000111000000001110111100001100",
			3511 => "0000000010000000000011001000000100",
			3512 => "11111110011000010011011100110101",
			3513 => "0000001010000000000001010100000100",
			3514 => "00000100010101110011011100110101",
			3515 => "00000010110100010011011100110101",
			3516 => "0000000100000000000101110000000100",
			3517 => "00000100001000000011011100110101",
			3518 => "0000000100000000001000110100010000",
			3519 => "0000000111000000001110110000001100",
			3520 => "0000001101000000000101100100000100",
			3521 => "11111110011000010011011100110101",
			3522 => "0000001000000000000110011100000100",
			3523 => "00000011001010110011011100110101",
			3524 => "00010000100110000011011100110101",
			3525 => "11111110011000000011011100110101",
			3526 => "0000000101000000001001110000001100",
			3527 => "0000001101000000001000111000000100",
			3528 => "11111110011111110011011100110101",
			3529 => "0000000101000000001000111100000100",
			3530 => "00000000101110010011011100110101",
			3531 => "11111110110101010011011100110101",
			3532 => "11111110010111100011011100110101",
			3533 => "0000000110000000000111101000011100",
			3534 => "0000001001000000000110101000011000",
			3535 => "0000000010000000000010110100001100",
			3536 => "0000000110000000001011111100001000",
			3537 => "0000000011000000000100000000000100",
			3538 => "00000000001111010011011111001001",
			3539 => "00000001110010000011011111001001",
			3540 => "11111110011011010011011111001001",
			3541 => "0000001100000000000111111000001000",
			3542 => "0000000110000000001110010100000100",
			3543 => "00000001101011110011011111001001",
			3544 => "00000000110111000011011111001001",
			3545 => "00000000010010100011011111001001",
			3546 => "11111110100101110011011111001001",
			3547 => "0000000100000000000101110000000100",
			3548 => "00000100001100000011011111001001",
			3549 => "0000000000000000000111000000010100",
			3550 => "0000001100000000000100001000010000",
			3551 => "0000001111000000000011001000000100",
			3552 => "11111110101101100011011111001001",
			3553 => "0000000001000000001001011000001000",
			3554 => "0000000110000000001101111100000100",
			3555 => "00000000000000000011011111001001",
			3556 => "00000011000101110011011111001001",
			3557 => "11111110111001010011011111001001",
			3558 => "11111110011011010011011111001001",
			3559 => "0000000111000000001110111100001000",
			3560 => "0000000010000000000011001000000100",
			3561 => "11111110100001110011011111001001",
			3562 => "00000001010000110011011111001001",
			3563 => "0000001100000000000000110000001100",
			3564 => "0000001110000000000001110100001000",
			3565 => "0000001101000000000100000000000100",
			3566 => "11111111011100100011011111001001",
			3567 => "00000000101001010011011111001001",
			3568 => "11111110111100010011011111001001",
			3569 => "11111110011001100011011111001001",
			3570 => "0000000110000000000111101000100000",
			3571 => "0000000001000000001110100000011100",
			3572 => "0000001111000000001101010100001000",
			3573 => "0000000111000000000000110000000100",
			3574 => "00000000000000110011100001110101",
			3575 => "11111110011110100011100001110101",
			3576 => "0000000110000000001110010100001000",
			3577 => "0000000100000000000010000000000100",
			3578 => "00000011010001000011100001110101",
			3579 => "00000001111100110011100001110101",
			3580 => "0000000111000000000100010100001000",
			3581 => "0000000100000000001111100000000100",
			3582 => "11111111111001000011100001110101",
			3583 => "00000001111100000011100001110101",
			3584 => "11111101111101110011100001110101",
			3585 => "11111110011011010011100001110101",
			3586 => "0000000111000000001110111100001100",
			3587 => "0000001111000000001110110000000100",
			3588 => "11111110011011010011100001110101",
			3589 => "0000000001000000000000011000000100",
			3590 => "00000010100000000011100001110101",
			3591 => "11111110100100010011100001110101",
			3592 => "0000001100000000000000111000001000",
			3593 => "0000001000000000001110111100000100",
			3594 => "11111111101000010011100001110101",
			3595 => "00000000011100010011100001110101",
			3596 => "0000000100000000001000110100011000",
			3597 => "0000000100000000001000000100001100",
			3598 => "0000001100000000000100001000001000",
			3599 => "0000001100000000000000001100000100",
			3600 => "11111110100110000011100001110101",
			3601 => "00000001110110110011100001110101",
			3602 => "11111110011001010011100001110101",
			3603 => "0000001100000000000000001100001000",
			3604 => "0000001100000000000000101000000100",
			3605 => "11111111000110010011100001110101",
			3606 => "00000100101101110011100001110101",
			3607 => "11111110101100110011100001110101",
			3608 => "0000001100000000001010000000001000",
			3609 => "0000001100000000001010000000000100",
			3610 => "11111110100001100011100001110101",
			3611 => "00000010000100000011100001110101",
			3612 => "11111110011000110011100001110101",
			3613 => "0000001100000000001010000000101000",
			3614 => "0000001111000000001010111100000100",
			3615 => "11111110010111110011100101100011",
			3616 => "0000000001000000000110000000010100",
			3617 => "0000000010000000001110000100001100",
			3618 => "0000001010000000000110011000000100",
			3619 => "00000011000011100011100101100011",
			3620 => "0000000000000000001100001000000100",
			3621 => "11111110101000100011100101100011",
			3622 => "00000000001111000011100101100011",
			3623 => "0000000000000000000100000100000100",
			3624 => "00000011001010110011100101100011",
			3625 => "00000100100011000011100101100011",
			3626 => "0000001010000000001000100100001000",
			3627 => "0000000101000000001101100000000100",
			3628 => "00000011100110110011100101100011",
			3629 => "00000000001110000011100101100011",
			3630 => "0000000100000000000011011000000100",
			3631 => "11111110010101100011100101100011",
			3632 => "00000000101101100011100101100011",
			3633 => "0000000111000000000100010100011100",
			3634 => "0000001010000000000111110100001000",
			3635 => "0000000010000000001101000100000100",
			3636 => "00000000101001100011100101100011",
			3637 => "00000011001001110011100101100011",
			3638 => "0000000010000000001010001000001100",
			3639 => "0000001011000000001010000000001000",
			3640 => "0000000101000000000100000000000100",
			3641 => "11111110100110100011100101100011",
			3642 => "00000000011101100011100101100011",
			3643 => "11111110011000010011100101100011",
			3644 => "0000000001000000000000011000000100",
			3645 => "00000011000000000011100101100011",
			3646 => "11111110100100010011100101100011",
			3647 => "0000000010000000000001001000010100",
			3648 => "0000001001000000000010001100001000",
			3649 => "0000000100000000000000010100000100",
			3650 => "00000100101011010011100101100011",
			3651 => "11111111000100000011100101100011",
			3652 => "0000001111000000001010011100000100",
			3653 => "11111110010110000011100101100011",
			3654 => "0000000101000000001000011000000100",
			3655 => "00000100110100000011100101100011",
			3656 => "11111110100011010011100101100011",
			3657 => "0000001000000000000101000100010100",
			3658 => "0000000111000000001110110000010000",
			3659 => "0000000010000000001110010000001000",
			3660 => "0000001010000000001010100000000100",
			3661 => "00000001111001100011100101100011",
			3662 => "11111110110100010011100101100011",
			3663 => "0000001101000000001011110100000100",
			3664 => "00001101000010110011100101100011",
			3665 => "00000000100100010011100101100011",
			3666 => "11111110010111110011100101100011",
			3667 => "0000001101000000001000111100001000",
			3668 => "0000000101000000001000111000000100",
			3669 => "11111110101000010011100101100011",
			3670 => "00000000000111000011100101100011",
			3671 => "11111110010111010011100101100011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1192, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(2454, initial_addr_3'length));
	end generate gen_rom_15;

	process (Clk)
	begin
		if rising_edge(Clk) then
			if (Re = '1') then
				-- Read from Addr
				Dout <= bank(to_integer(unsigned(Addr)));
			else
				Dout <= (others => '0');
			end if;
		end if;
	end process;
end Behavioral;
